
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal DATA2_I_30_port, DATA2_I_28_port, DATA2_I_27_port, DATA2_I_26_port, 
      DATA2_I_25_port, DATA2_I_24_port, DATA2_I_23_port, DATA2_I_22_port, 
      DATA2_I_21_port, DATA2_I_20_port, DATA2_I_19_port, DATA2_I_18_port, 
      DATA2_I_17_port, DATA2_I_16_port, DATA2_I_15_port, DATA2_I_14_port, 
      DATA2_I_13_port, DATA2_I_12_port, DATA2_I_11_port, DATA2_I_10_port, 
      DATA2_I_9_port, DATA2_I_8_port, DATA2_I_7_port, DATA2_I_6_port, 
      DATA2_I_5_port, DATA2_I_4_port, DATA2_I_3_port, DATA2_I_2_port, 
      DATA2_I_1_port, DATA2_I_0_port, data1_mul_15_port, data1_mul_0_port, 
      data2_mul_2_port, data2_mul_1_port, N2517, N2518, N2519, N2520, N2521, 
      N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n554, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_34_port, 
      boothmul_pipelined_i_muxes_in_4_33_port, 
      boothmul_pipelined_i_muxes_in_4_32_port, 
      boothmul_pipelined_i_muxes_in_4_31_port, 
      boothmul_pipelined_i_muxes_in_4_30_port, 
      boothmul_pipelined_i_muxes_in_4_29_port, 
      boothmul_pipelined_i_muxes_in_4_28_port, 
      boothmul_pipelined_i_muxes_in_4_27_port, 
      boothmul_pipelined_i_sum_B_in_7_14_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_6_12_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_5_10_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_4_8_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_3_6_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_4_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n1353, 
      n1429, n2808, n3020, n3026, n3027, n3028, n3029, n3030, n3036, n3794, 
      n3800, n3820, n3821, n3822, n3831, n3834, n3835, n3836, n3837, n3838, 
      n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, 
      n3854, n3856, n3858, n3859, n3860, n3861, n3862, n3863, n3865, n3866, 
      n3867, n3875, n3885, n3888, n3892, n3893, n3894, n3895, n3896, n3897, 
      n3900, n3902, n3904, n3905, n3910, n3911, n3918, n3919, n3920, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3940, n3941, n3943, n3944, 
      n3945, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3956, 
      n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
      n3967, n3968, n3970, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
      n3979, n3980, n3981, n3982, n3983, n3984, n3986, n3989, n3990, n3991, 
      n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, 
      n4003, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, 
      n4016, n4017, n4018, n4020, n4025, n4026, n4027, n4033, n4034, n4035, 
      n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, 
      n4046, n4048, n4055, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
      n4067, n4068, n4069, n4070, n4073, n4074, n4075, n4078, n4111, n4175, 
      n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, 
      n4186, n4187, n4188, n4189, n4190, n4192, n4199, n4200, n4205, n4212, 
      n4216, n4220, n4257, n4263, n4266, n4270, n4274, n4280, n4293, n4295, 
      n4298, n4302, n4303, n4308, n4310, n4316, n4319, n4325, n4395, n4421, 
      n4476, n4506, n6095, n6106, n6174, n6177, n6179, n6184, n6187, n6191, 
      n6192, n6196, n6197, n6198, n6204, n6205, n6206, n6207, n6208, n6212, 
      n6213, n6214, n6215, n6237, n6238, n6240, n6241, n6260, n6261, n6267, 
      n6268, n6294, n6314, n6338, n6340, n6351, n6367, n6381, n6422, n6502, 
      n6505, n6506, n6510, n6516, n6517, n6523, n6524, n6525, n6529, n6530, 
      n6533, n6541, n6561, n6617, n6618, n6671, n6675, n6676, n6677, n6733, 
      n6739, n6740, n6742, n6744, n6749, n6762, n6763, n6793, n6837, n6850, 
      n6852, n6853, n6858, n6860, n6862, n6865, n6869, n6870, n6871, n6874, 
      n6876, n6880, n6881, n6888, n6889, n6896, n6899, n6905, n6908, n6932, 
      n6935, n6938, n6949, n6957, n6980, n7007, n7047, n7086, n7097, n7114, 
      n7134, n7147, n7150, n7153, n7166, n7284, n7285, n7286, n7287, n7325, 
      n7326, n7332, n7333, n7339, n7340, n7449, n7481, n7483, n7485, n7654, 
      n7659, n7759, n7769, n7822, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, 
      n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8553, n8554, n8555, 
      n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, 
      n8566, n8567, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, 
      n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8586, n8587, n8588, 
      n8589, n8591, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, 
      n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, 
      n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, 
      n8621, n8622, n8623, n8626, n8627, n8628, n8629, n8630, n8631, n8632, 
      n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, 
      n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, 
      n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, 
      n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, 
      n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, 
      n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, 
      n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, 
      n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, 
      n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, 
      n8723, n8724, n8725, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8744, 
      n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, 
      n8755, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, 
      n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, 
      n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, 
      n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, 
      n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, 
      n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, 
      n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, 
      n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, 
      n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, 
      n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8856, 
      n8857, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, 
      n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, 
      n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, 
      n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, 
      n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, 
      n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, 
      n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, 
      n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, 
      n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, 
      n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, 
      n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, 
      n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, 
      n8980, n8981, n8983, n8984, n8985, n8986, n8988, n8989, n8990, n8991, 
      n8992, n8993, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, 
      n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, 
      n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, 
      n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, 
      n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9044, 
      n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, 
      n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, 
      n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, 
      n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, 
      n9085, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, 
      n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, 
      n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, 
      n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, 
      n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, 
      n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, 
      n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, 
      n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, 
      n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, 
      n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, 
      n9192, n9193, n9194, n9195, n9196, n9198, n9199, n9200, n9201, n9202, 
      n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, 
      n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, 
      n9223, n9225, n11300, n11301, n11302, n11303, n11304, n11305, n11306, 
      n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, 
      n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, 
      n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
      n11334, n11335, n11337, n11338, n11339, n11340, n1799, n1800, n1801, 
      n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, 
      n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, 
      n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n11377, n11378, n11379, n11380, n11381, n11382, n11383, 
      n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, 
      n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, 
      n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, 
      n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, 
      n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, 
      n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, 
      n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, 
      n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, 
      n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, 
      n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, 
      n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, 
      n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, 
      n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, 
      n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, 
      n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, 
      n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, 
      n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, 
      n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, 
      n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, 
      n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, 
      n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, 
      n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, 
      n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, 
      n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, 
      n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, 
      n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, 
      n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, 
      n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, 
      n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, 
      n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, 
      n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, 
      n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, 
      n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, 
      n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, 
      n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, 
      n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, 
      n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, 
      n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, 
      n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, 
      n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, 
      n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, 
      n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, 
      n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, 
      n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, 
      n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, 
      n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, 
      n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, 
      n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, 
      n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, 
      n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, 
      n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, 
      n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, 
      n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, 
      n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, 
      n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, 
      n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, 
      n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, 
      n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, 
      n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, 
      n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, 
      n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, 
      n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, 
      n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, 
      n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, 
      n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, 
      n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, 
      n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, 
      n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, 
      n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, 
      n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, 
      n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, 
      n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, 
      n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, 
      n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, 
      n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, 
      n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, 
      n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, 
      n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, 
      n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, 
      n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, 
      n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, 
      n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, 
      n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, 
      n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, 
      n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, 
      n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, 
      n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, 
      n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, 
      n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, 
      n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, 
      n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, 
      n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, 
      n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, 
      n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, 
      n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, 
      n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, 
      n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, 
      n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, 
      n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, 
      n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, 
      n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, 
      n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, 
      n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, 
      n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, 
      n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, 
      n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, 
      n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, 
      n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, 
      n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, 
      n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, 
      n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, 
      n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, 
      n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, 
      n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, 
      n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, 
      n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, 
      n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, 
      n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, 
      n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, 
      n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, 
      n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, 
      n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, 
      n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, 
      n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, 
      n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, 
      n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, 
      n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, 
      n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, 
      n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, 
      n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, 
      n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, 
      n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, 
      n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, 
      n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, 
      n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, 
      n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, 
      n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, 
      n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, 
      n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, 
      n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, 
      n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, 
      n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, 
      n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, 
      n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, 
      n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, 
      n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, 
      n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, 
      n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, 
      n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, 
      n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, 
      n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, 
      n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, 
      n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, 
      n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, 
      n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, 
      n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, 
      n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, 
      n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, 
      n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, 
      n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, 
      n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, 
      n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, 
      n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, 
      n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, 
      n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, 
      n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, 
      n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, 
      n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, 
      n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, 
      n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, 
      n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, 
      n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, 
      n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, 
      n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, 
      n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, 
      n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, 
      n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, 
      n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, 
      n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, 
      n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, 
      n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, 
      n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, 
      n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, 
      n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, 
      n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, 
      n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, 
      n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, 
      n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, 
      n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, 
      n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, 
      n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, 
      n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, 
      n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, 
      n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, 
      n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, 
      n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, 
      n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, 
      n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, 
      n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, 
      n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, 
      n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, 
      n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, 
      n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, 
      n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, 
      n13220, n13221, n13222, n13223, n13224, n13225, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634 : std_logic;

begin
   
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n554, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n554, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n13225, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n13225, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n554, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n554, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n554, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n554, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n554, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n554, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n13225, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n554, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n554, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n554, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n554, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n554, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n554, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n13225, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n554, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n13225, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n13225, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n13225, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n13225, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n554, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n554, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n554, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n554, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n554, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n13225, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n7822, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_27_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_28_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_29_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_30_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_31_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_32_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_33_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_34_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => n9225, GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => n9223, GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => n9222, GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => n9221, GN => n7822, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n7822, Q => 
                           n4325);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n7822, Q => 
                           n4319);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n7822, Q => 
                           n4316);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n7822, Q => 
                           n4310);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n7822, Q => 
                           n4308);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n7822, Q => 
                           n4303);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n7822, Q => 
                           n4302);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n7822, Q => 
                           n4298);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n7822, Q => 
                           n7769);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n7822, Q => 
                           n4295);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n7822, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n7822, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n554, Q => n4293);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1825, B => n1826, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1824, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1823, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1822, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1820, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1819, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1818, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1817, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1816, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1815, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1814, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1813, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1812, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1811, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1810, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3036,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => n4048);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => n4046);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => n4045);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => n4044);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => n4043);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => n4042);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => n4041);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => n4040);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => n4039);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => n4038);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => n4037);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => n4036);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => n4035);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => n4034);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1004, S => n4033);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => n8792, 
                           CI => n3026, CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => n4027);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => n8791, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => n8790, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => n8789, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => n8788, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => n8787, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => n8786, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => n8785, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => n8784, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => n8783, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => n8782, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => n8781, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => n8780, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => n8779, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => n8779, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => n4026, S => n4025);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n8535, B => n8778, CI => n8771, CO => n_1005, S => 
                           boothmul_pipelined_i_sum_B_in_3_22_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3030,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => n4020);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => n4018);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => n4017);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => n4016);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => n4015);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => n4014);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => n4013);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => n4012);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => n4011);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => n4010);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n8813, B => n8772, CI => n8763, CO => n4009, S => 
                           n4008);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n8812, B => n8770, CI => n4009, CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n8811, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n8810, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n8534, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1006, S => n4007);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => n4018, 
                           CI => n3029, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => n4003);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => n4017, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => n4016, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => n4001);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => n4015, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => n4000);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => n4014, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => n3999);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => n4013, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => n3998);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => n4012, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => n3997);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           n8928, B => n8764, CI => n8751, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => n3996);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           n8927, B => n8762, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => n3995);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           n8926, B => n4008, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => n3994);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n8925, B => boothmul_pipelined_i_sum_B_in_4_19_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => n3993);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n8924, B => boothmul_pipelined_i_sum_B_in_4_20_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => n3992);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n8923, B => boothmul_pipelined_i_sum_B_in_4_21_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => n3991, S => n3990);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n8922, B => n4007, CI => n3991, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n8921, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n8549, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1007, S => n3989);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => n8755, 
                           CI => n3028, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => n3986);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => n8754, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => n8753, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => n3984);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => n8752, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => n3983);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => n8750, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => n3982);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => n3996, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => n3981);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => n3995, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => n3980);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => n3994, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => n3979);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => n3993, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => n3978);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => n3992, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => n3977);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => n3990, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => n3976);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => n3975);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n8920, B => n8749, CI => n8733, CO => n3974, S => 
                           n3973);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n8919, B => n8748, CI => n3974, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n8918, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n8548, B => n8748, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1008, S => n3972);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => n8742, 
                           CI => n3027, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => n3970);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => n8741, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => n8740, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => n3968);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => n8739, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => n3967);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => n8738, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => n3966);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => n8737, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => n3965);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => n8736, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => n3964);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => n8735, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => n3963);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => n8734, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => n3962);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => n8732, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => n3961);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => n3973, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => n3960);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => n3959);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n8917, B => n8731, CI => n8716, CO => n3958, S => 
                           n3957);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n8916, B => n8730, CI => n3958, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n8915, B => n8730, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n8547, B => n8730, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1009, S => n3956);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => n8725, 
                           CI => n3020, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => n3954);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => n8724, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => n3953);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => n8723, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => n3952);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => n8722, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => n3951);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => n8721, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => n3950);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => n8720, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => n3949);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => n8719, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => n3948);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => n8718, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => n3947);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => n8717, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => n3945);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => n8715, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => n3944);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => n3957, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => n3943);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => n3941);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n8914, B => n8714, CI => n8689, CO => n3940, S => 
                           n3938);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n8913, B => n8713, CI => n3940, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => n3937);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           n8912, B => n8713, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => n3936);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           n8911, B => n8713, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => n3935);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           n8911, B => n8713, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1010, S => n3934);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n7822, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n554, Q => 
                           DATA2_I_30_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port);
   clk_r_REG4782_S3 : DFFS_X1 port map( D => n1859, CK => clk, SN => rst_BAR, Q
                           => n13149, QN => n9225);
   clk_r_REG4928_S3 : DFFS_X1 port map( D => n1860, CK => clk, SN => rst_BAR, Q
                           => n_1011, QN => n9223);
   clk_r_REG5584_S3 : DFFR_X1 port map( D => DATA1(1), CK => clk, RN => n11392,
                           Q => n9222, QN => n11332);
   clk_r_REG5920_S5 : DFFR_X1 port map( D => DATA1(0), CK => clk, RN => n11377,
                           Q => n9221, QN => n13173);
   clk_r_REG6781_S1 : DFFR_X1 port map( D => cin, CK => clk, RN => n11390, Q =>
                           n9220, QN => n_1012);
   clk_r_REG4486_S4 : DFFR_X1 port map( D => n7654, CK => clk, RN => n11397, Q 
                           => n_1013, QN => n9219);
   clk_r_REG4365_S4 : DFFS_X1 port map( D => n4506, CK => clk, SN => n11389, Q 
                           => n_1014, QN => n9218);
   clk_r_REG4348_S4 : DFFR_X1 port map( D => n7659, CK => clk, RN => n11392, Q 
                           => n13169, QN => n9217);
   clk_r_REG4440_S4 : DFFS_X1 port map( D => n7759, CK => clk, SN => n11378, Q 
                           => n13145, QN => n9216);
   clk_r_REG4443_S4 : DFFR_X1 port map( D => n4476, CK => clk, RN => n11382, Q 
                           => n13140, QN => n9215);
   clk_r_REG6651_S3 : DFFS_X1 port map( D => n1832, CK => clk, SN => n11388, Q 
                           => n9214, QN => n_1015);
   clk_r_REG6648_S3 : DFFR_X1 port map( D => FUNC(2), CK => clk, RN => n11399, 
                           Q => n_1016, QN => n9213);
   clk_r_REG6652_S3 : DFFS_X1 port map( D => FUNC(3), CK => clk, SN => n11400, 
                           Q => n_1017, QN => n9212);
   clk_r_REG3851_S4 : DFFS_X1 port map( D => n13224, CK => clk, SN => n11388, Q
                           => n9211, QN => n_1018);
   clk_r_REG3850_S4 : DFFR_X1 port map( D => n6095, CK => clk, RN => n11389, Q 
                           => n9210, QN => n_1019);
   clk_r_REG6647_S3 : DFFS_X1 port map( D => n1835, CK => clk, SN => n11384, Q 
                           => n_1020, QN => n9209);
   clk_r_REG5658_S4 : DFFS_X1 port map( D => n1846, CK => clk, SN => n11400, Q 
                           => n9208, QN => n_1021);
   clk_r_REG3557_S5 : DFFR_X1 port map( D => n6106, CK => clk, RN => n11382, Q 
                           => n_1022, QN => n9207);
   clk_r_REG4783_S3 : DFFS_X1 port map( D => n1859, CK => clk, SN => rst_BAR, Q
                           => n9206, QN => n_1023);
   clk_r_REG4929_S3 : DFFS_X1 port map( D => n1860, CK => clk, SN => n11378, Q 
                           => n9205, QN => n13177);
   clk_r_REG5258_S4 : DFFS_X1 port map( D => n1839, CK => clk, SN => n11396, Q 
                           => n9204, QN => n_1024);
   clk_r_REG4400_S4 : DFFS_X1 port map( D => n1841, CK => clk, SN => n11378, Q 
                           => n9203, QN => n_1025);
   clk_r_REG4416_S4 : DFFR_X1 port map( D => n1849, CK => clk, RN => n11392, Q 
                           => n9202, QN => n_1026);
   clk_r_REG4122_S4 : DFFR_X1 port map( D => n1854, CK => clk, RN => n11401, Q 
                           => n9201, QN => n_1027);
   clk_r_REG3764_S4 : DFFR_X1 port map( D => n1844, CK => clk, RN => n11401, Q 
                           => n9200, QN => n_1028);
   clk_r_REG3779_S4 : DFFS_X1 port map( D => n1842, CK => clk, SN => n11403, Q 
                           => n9199, QN => n_1029);
   clk_r_REG3927_S4 : DFFS_X1 port map( D => n1850, CK => clk, SN => n11400, Q 
                           => n9198, QN => n_1030);
   clk_r_REG3924_S4 : DFFS_X1 port map( D => n1851, CK => clk, SN => n11378, Q 
                           => n_1031, QN => n13201);
   clk_r_REG3974_S4 : DFFR_X1 port map( D => n1856, CK => clk, RN => n11401, Q 
                           => n9196, QN => n_1032);
   clk_r_REG3972_S4 : DFFS_X1 port map( D => n1857, CK => clk, SN => n11377, Q 
                           => n9195, QN => n13152);
   clk_r_REG3922_S4 : DFFR_X1 port map( D => n1855, CK => clk, RN => n11388, Q 
                           => n9194, QN => n_1033);
   clk_r_REG4607_S5 : DFFR_X1 port map( D => n1828, CK => clk, RN => n11379, Q 
                           => n9193, QN => n13209);
   clk_r_REG3633_S5 : DFFR_X1 port map( D => n1799, CK => clk, RN => n11379, Q 
                           => n9192, QN => n13211);
   clk_r_REG3933_S4 : DFFS_X1 port map( D => n1858, CK => clk, SN => n11396, Q 
                           => n9191, QN => n_1034);
   clk_r_REG4615_S4 : DFFS_X1 port map( D => n1836, CK => clk, SN => n11377, Q 
                           => n9190, QN => n_1035);
   clk_r_REG4133_S5 : DFFS_X1 port map( D => n11327, CK => clk, SN => n11378, Q
                           => n9189, QN => n_1036);
   clk_r_REG4144_S5 : DFFS_X1 port map( D => n11305, CK => clk, SN => n11381, Q
                           => n9188, QN => n_1037);
   clk_r_REG4392_S4 : DFFS_X1 port map( D => n13221, CK => clk, SN => n11379, Q
                           => n9187, QN => n_1038);
   clk_r_REG4397_S4 : DFFS_X1 port map( D => n13221, CK => clk, SN => n11396, Q
                           => n9186, QN => n_1039);
   clk_r_REG4458_S4 : DFFR_X1 port map( D => n1872, CK => clk, RN => n11398, Q 
                           => n9185, QN => n_1040);
   clk_r_REG4424_S4 : DFFS_X1 port map( D => n13220, CK => clk, SN => n11390, Q
                           => n9184, QN => n_1041);
   clk_r_REG4362_S4 : DFFS_X1 port map( D => n1876, CK => clk, SN => n11377, Q 
                           => n9183, QN => n13143);
   clk_r_REG4454_S4 : DFFS_X1 port map( D => n11312, CK => clk, SN => n11401, Q
                           => n9182, QN => n13141);
   clk_r_REG4374_S4 : DFFS_X1 port map( D => n11318, CK => clk, SN => n11399, Q
                           => n9181, QN => n13144);
   clk_r_REG4382_S4 : DFFS_X1 port map( D => n11315, CK => clk, SN => n11377, Q
                           => n9180, QN => n_1042);
   clk_r_REG3585_S4 : DFFS_X1 port map( D => DATA2(31), CK => clk, SN => n11400
                           , Q => n9179, QN => n_1043);
   clk_r_REG4408_S4 : DFFS_X1 port map( D => n1848, CK => clk, SN => n11378, Q 
                           => n9178, QN => n_1044);
   clk_r_REG4407_S4 : DFFS_X1 port map( D => n1847, CK => clk, SN => n11402, Q 
                           => n9177, QN => n_1045);
   clk_r_REG4425_S4 : DFFS_X1 port map( D => n1843, CK => clk, SN => n11378, Q 
                           => n9176, QN => n_1046);
   clk_r_REG4488_S4 : DFFS_X1 port map( D => n7654, CK => clk, SN => n11379, Q 
                           => n9175, QN => n_1047);
   clk_r_REG4140_S4 : DFFR_X1 port map( D => n1829, CK => clk, RN => n11398, Q 
                           => n9174, QN => n_1048);
   clk_r_REG4353_S4 : DFFR_X1 port map( D => n11321, CK => clk, RN => n11397, Q
                           => n9173, QN => n_1049);
   clk_r_REG4493_S5 : DFFS_X1 port map( D => n1821, CK => clk, SN => n11396, Q 
                           => n9172, QN => n_1050);
   clk_r_REG6451_S5 : DFFS_X1 port map( D => n1801, CK => clk, SN => n11403, Q 
                           => n9171, QN => n_1051);
   clk_r_REG4670_S5 : DFFS_X1 port map( D => n1807, CK => clk, SN => n11401, Q 
                           => n9170, QN => n_1052);
   clk_r_REG4476_S4 : DFFS_X1 port map( D => n11316, CK => clk, SN => n11402, Q
                           => n9169, QN => n_1053);
   clk_r_REG4336_S4 : DFFR_X1 port map( D => n1877, CK => clk, RN => n11388, Q 
                           => n9168, QN => n_1054);
   clk_r_REG4347_S4 : DFFS_X1 port map( D => n11319, CK => clk, SN => n11394, Q
                           => n9167, QN => n13172);
   clk_r_REG4463_S4 : DFFS_X1 port map( D => n11322, CK => clk, SN => n11377, Q
                           => n9166, QN => n13157);
   clk_r_REG4446_S4 : DFFS_X1 port map( D => n1866, CK => clk, SN => n11403, Q 
                           => n9165, QN => n13153);
   clk_r_REG4345_S4 : DFFR_X1 port map( D => n1873, CK => clk, RN => n11394, Q 
                           => n9164, QN => n_1055);
   clk_r_REG4470_S4 : DFFS_X1 port map( D => n11324, CK => clk, SN => n11378, Q
                           => n9163, QN => n_1056);
   clk_r_REG4339_S4 : DFFR_X1 port map( D => n1871, CK => clk, RN => n11387, Q 
                           => n9162, QN => n13180);
   clk_r_REG3911_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_102_port, CK => clk,
                           RN => n11398, Q => n9161, QN => n_1057);
   clk_r_REG3912_S6 : DFFR_X1 port map( D => n9161, CK => clk, RN => n11388, Q 
                           => n9160, QN => n_1058);
   clk_r_REG3913_S7 : DFFR_X1 port map( D => n9160, CK => clk, RN => n11380, Q 
                           => n9159, QN => n_1059);
   clk_r_REG3902_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_103_port, CK => clk,
                           RN => n11391, Q => n9158, QN => n_1060);
   clk_r_REG3905_S6 : DFFR_X1 port map( D => n9158, CK => clk, RN => n11385, Q 
                           => n9157, QN => n_1061);
   clk_r_REG3906_S7 : DFFR_X1 port map( D => n9157, CK => clk, RN => n11390, Q 
                           => n9156, QN => n_1062);
   clk_r_REG3963_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_104_port, CK => clk,
                           RN => n11384, Q => n9155, QN => n_1063);
   clk_r_REG3965_S6 : DFFR_X1 port map( D => n9155, CK => clk, RN => n11397, Q 
                           => n9154, QN => n_1064);
   clk_r_REG3966_S7 : DFFR_X1 port map( D => n9154, CK => clk, RN => n11391, Q 
                           => n9153, QN => n_1065);
   clk_r_REG4109_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_105_port, CK => clk,
                           RN => n11398, Q => n9152, QN => n_1066);
   clk_r_REG4110_S6 : DFFR_X1 port map( D => n9152, CK => clk, RN => n11388, Q 
                           => n9151, QN => n_1067);
   clk_r_REG4111_S7 : DFFR_X1 port map( D => n9151, CK => clk, RN => n11380, Q 
                           => n9150, QN => n_1068);
   clk_r_REG4106_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_106_port, CK => clk,
                           RN => n11379, Q => n9149, QN => n_1069);
   clk_r_REG4107_S6 : DFFR_X1 port map( D => n9149, CK => clk, RN => n11381, Q 
                           => n9148, QN => n_1070);
   clk_r_REG4108_S7 : DFFR_X1 port map( D => n9148, CK => clk, RN => n11393, Q 
                           => n9147, QN => n_1071);
   clk_r_REG4102_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_107_port, CK => clk,
                           RN => n11394, Q => n9146, QN => n_1072);
   clk_r_REG4103_S6 : DFFR_X1 port map( D => n9146, CK => clk, RN => n11402, Q 
                           => n9145, QN => n_1073);
   clk_r_REG4104_S7 : DFFR_X1 port map( D => n9145, CK => clk, RN => n11380, Q 
                           => n9144, QN => n_1074);
   clk_r_REG4099_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_108_port, CK => clk,
                           RN => n11390, Q => n9143, QN => n_1075);
   clk_r_REG4100_S6 : DFFR_X1 port map( D => n9143, CK => clk, RN => n11388, Q 
                           => n9142, QN => n_1076);
   clk_r_REG4101_S7 : DFFR_X1 port map( D => n9142, CK => clk, RN => n11392, Q 
                           => n9141, QN => n_1077);
   clk_r_REG4156_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_109_port, CK => clk,
                           RN => n11383, Q => n9140, QN => n_1078);
   clk_r_REG4157_S6 : DFFR_X1 port map( D => n9140, CK => clk, RN => n11384, Q 
                           => n9139, QN => n_1079);
   clk_r_REG4158_S7 : DFFR_X1 port map( D => n9139, CK => clk, RN => n11403, Q 
                           => n9138, QN => n_1080);
   clk_r_REG4153_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_110_port, CK => clk,
                           RN => n11401, Q => n9137, QN => n_1081);
   clk_r_REG4154_S6 : DFFR_X1 port map( D => n9137, CK => clk, RN => n11399, Q 
                           => n9136, QN => n_1082);
   clk_r_REG4155_S7 : DFFR_X1 port map( D => n9136, CK => clk, RN => n11383, Q 
                           => n9135, QN => n_1083);
   clk_r_REG4500_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_111_port, CK => clk,
                           RN => n11393, Q => n9134, QN => n_1084);
   clk_r_REG4501_S6 : DFFR_X1 port map( D => n9134, CK => clk, RN => n11401, Q 
                           => n9133, QN => n_1085);
   clk_r_REG4502_S7 : DFFR_X1 port map( D => n9133, CK => clk, RN => n11382, Q 
                           => n9132, QN => n_1086);
   clk_r_REG4497_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_112_port, CK => clk,
                           RN => n11380, Q => n9131, QN => n_1087);
   clk_r_REG4498_S6 : DFFR_X1 port map( D => n9131, CK => clk, RN => n11385, Q 
                           => n9130, QN => n_1088);
   clk_r_REG4499_S7 : DFFR_X1 port map( D => n9130, CK => clk, RN => n11391, Q 
                           => n9129, QN => n_1089);
   clk_r_REG4494_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_113_port, CK => clk,
                           RN => n11387, Q => n9128, QN => n_1090);
   clk_r_REG4495_S6 : DFFR_X1 port map( D => n9128, CK => clk, RN => n11392, Q 
                           => n9127, QN => n_1091);
   clk_r_REG4496_S7 : DFFR_X1 port map( D => n9127, CK => clk, RN => n11389, Q 
                           => n9126, QN => n_1092);
   clk_r_REG4784_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_114_port, CK => clk,
                           RN => n11403, Q => n9125, QN => n_1093);
   clk_r_REG4785_S6 : DFFR_X1 port map( D => n9125, CK => clk, RN => n11394, Q 
                           => n9124, QN => n_1094);
   clk_r_REG4786_S7 : DFFR_X1 port map( D => n9124, CK => clk, RN => rst_BAR, Q
                           => n9123, QN => n_1095);
   clk_r_REG4930_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_115_port, CK => clk,
                           RN => n11384, Q => n9122, QN => n_1096);
   clk_r_REG4931_S6 : DFFR_X1 port map( D => n9122, CK => clk, RN => n11386, Q 
                           => n9121, QN => n_1097);
   clk_r_REG4932_S7 : DFFR_X1 port map( D => n9121, CK => clk, RN => n11393, Q 
                           => n9120, QN => n_1098);
   clk_r_REG5586_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_0_116_port, CK => clk,
                           RN => n11383, Q => n9119, QN => n_1099);
   clk_r_REG5587_S6 : DFFR_X1 port map( D => n9119, CK => clk, RN => n11401, Q 
                           => n9118, QN => n_1100);
   clk_r_REG5588_S7 : DFFR_X1 port map( D => n9118, CK => clk, RN => n11383, Q 
                           => n9117, QN => n_1101);
   clk_r_REG3984_S5 : DFFS_X1 port map( D => n11330, CK => clk, SN => n11380, Q
                           => n9116, QN => n_1102);
   clk_r_REG6000_S5 : DFFS_X1 port map( D => n1803, CK => clk, SN => n11400, Q 
                           => n9115, QN => n_1103);
   clk_r_REG5997_S5 : DFFS_X1 port map( D => n1804, CK => clk, SN => n11403, Q 
                           => n9114, QN => n_1104);
   clk_r_REG4473_S4 : DFFR_X1 port map( D => n11311, CK => clk, RN => n11386, Q
                           => n9113, QN => n_1105);
   clk_r_REG4330_S4 : DFFS_X1 port map( D => n11317, CK => clk, SN => n11378, Q
                           => n9112, QN => n_1106);
   clk_r_REG4467_S4 : DFFS_X1 port map( D => n11313, CK => clk, SN => n11399, Q
                           => n9111, QN => n_1107);
   clk_r_REG6649_S3 : DFFS_X1 port map( D => n7166, CK => clk, SN => n11390, Q 
                           => n9110, QN => n_1108);
   clk_r_REG4483_S4 : DFFS_X1 port map( D => n1834, CK => clk, SN => n11381, Q 
                           => n9109, QN => n13207);
   clk_r_REG4146_S5 : DFFS_X1 port map( D => n7147, CK => clk, SN => n11399, Q 
                           => n9108, QN => n_1109);
   clk_r_REG4341_S4 : DFFS_X1 port map( D => n11320, CK => clk, SN => n11403, Q
                           => n9107, QN => n13193);
   clk_r_REG4361_S4 : DFFS_X1 port map( D => n11323, CK => clk, SN => n11395, Q
                           => n9106, QN => n13167);
   clk_r_REG4439_S4 : DFFS_X1 port map( D => n1868, CK => clk, SN => n11397, Q 
                           => n9105, QN => n13179);
   clk_r_REG4375_S4 : DFFS_X1 port map( D => n11318, CK => clk, SN => n11389, Q
                           => n9104, QN => n_1110);
   clk_r_REG4368_S4 : DFFS_X1 port map( D => n11314, CK => clk, SN => n11401, Q
                           => n9103, QN => n_1111);
   clk_r_REG4350_S4 : DFFS_X1 port map( D => n7659, CK => clk, SN => n11379, Q 
                           => n9102, QN => n13196);
   clk_r_REG4371_S4 : DFFS_X1 port map( D => n1874, CK => clk, SN => n11400, Q 
                           => n9101, QN => n_1112);
   clk_r_REG4481_S4 : DFFS_X1 port map( D => n1833, CK => clk, SN => n11379, Q 
                           => n9100, QN => n13161);
   clk_r_REG4485_S4 : DFFS_X1 port map( D => n1878, CK => clk, SN => n11398, Q 
                           => n9099, QN => n_1113);
   clk_r_REG4356_S4 : DFFS_X1 port map( D => n1870, CK => clk, SN => n11377, Q 
                           => n9098, QN => n_1114);
   clk_r_REG3914_S5 : DFFR_X1 port map( D => n1809, CK => clk, RN => n11397, Q 
                           => n9097, QN => n_1115);
   clk_r_REG3915_S6 : DFFR_X1 port map( D => n9097, CK => clk, RN => n11398, Q 
                           => n9096, QN => n_1116);
   clk_r_REG3916_S7 : DFFR_X1 port map( D => n9096, CK => clk, RN => n11383, Q 
                           => n9095, QN => n_1117);
   clk_r_REG4450_S4 : DFFS_X1 port map( D => n1869, CK => clk, SN => n11387, Q 
                           => n9094, QN => n_1118);
   clk_r_REG4322_S5 : DFFR_X1 port map( D => n11331, CK => clk, RN => n11391, Q
                           => n9093, QN => n_1119);
   clk_r_REG4141_S5 : DFFS_X1 port map( D => n1827, CK => clk, SN => n11381, Q 
                           => n_1120, QN => n11306);
   clk_r_REG4066_S6 : DFFS_X1 port map( D => n11328, CK => clk, SN => n11377, Q
                           => n_1121, QN => n11307);
   clk_r_REG3861_S7 : DFFS_X1 port map( D => n11326, CK => clk, SN => n11386, Q
                           => n_1122, QN => n11308);
   clk_r_REG3956_S8 : DFFS_X1 port map( D => n11329, CK => clk, SN => n11379, Q
                           => n_1123, QN => n11309);
   clk_r_REG5921_S7 : DFFR_X1 port map( D => data1_mul_0_port, CK => clk, RN =>
                           n11387, Q => n_1124, QN => n11310);
   clk_r_REG5922_S8 : DFFS_X1 port map( D => n11310, CK => clk, SN => n11402, Q
                           => n11300, QN => n_1125);
   clk_r_REG5923_S9 : DFFS_X1 port map( D => n11300, CK => clk, SN => n11378, Q
                           => n11301, QN => n_1126);
   clk_r_REG5589_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_64_port, CK => clk, 
                           RN => n11402, Q => n9085, QN => n_1127);
   clk_r_REG5590_S6 : DFFR_X1 port map( D => n9085, CK => clk, RN => n11383, Q 
                           => n9084, QN => n_1128);
   clk_r_REG5591_S7 : DFFR_X1 port map( D => n9084, CK => clk, RN => n11388, Q 
                           => n9083, QN => n_1129);
   clk_r_REG4933_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_63_port, CK => clk, 
                           RN => n11387, Q => n9082, QN => n_1130);
   clk_r_REG4934_S6 : DFFR_X1 port map( D => n9082, CK => clk, RN => n11379, Q 
                           => n9081, QN => n_1131);
   clk_r_REG4935_S7 : DFFR_X1 port map( D => n9081, CK => clk, RN => n11399, Q 
                           => n9080, QN => n_1132);
   clk_r_REG4787_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_62_port, CK => clk, 
                           RN => n11380, Q => n9079, QN => n_1133);
   clk_r_REG4788_S6 : DFFR_X1 port map( D => n9079, CK => clk, RN => n11394, Q 
                           => n9078, QN => n_1134);
   clk_r_REG4789_S7 : DFFR_X1 port map( D => n9078, CK => clk, RN => n11384, Q 
                           => n9077, QN => n_1135);
   clk_r_REG4503_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_61_port, CK => clk, 
                           RN => n11390, Q => n9076, QN => n_1136);
   clk_r_REG4504_S6 : DFFR_X1 port map( D => n9076, CK => clk, RN => n11394, Q 
                           => n9075, QN => n_1137);
   clk_r_REG4505_S7 : DFFR_X1 port map( D => n9075, CK => clk, RN => n11382, Q 
                           => n9074, QN => n_1138);
   clk_r_REG4575_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_60_port, CK => clk, 
                           RN => n11382, Q => n9073, QN => n_1139);
   clk_r_REG4576_S10 : DFFR_X1 port map( D => n9073, CK => clk, RN => n11385, Q
                           => n9072, QN => n_1140);
   clk_r_REG4577_S11 : DFFR_X1 port map( D => n9072, CK => clk, RN => n11386, Q
                           => n9071, QN => n_1141);
   clk_r_REG5911_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_59_port, CK => clk, 
                           RN => n11387, Q => n9070, QN => n_1142);
   clk_r_REG5912_S10 : DFFR_X1 port map( D => n9070, CK => clk, RN => n11387, Q
                           => n9069, QN => n_1143);
   clk_r_REG5913_S11 : DFFR_X1 port map( D => n9069, CK => clk, RN => n11400, Q
                           => n9068, QN => n_1144);
   clk_r_REG4159_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_34_port, CK => clk, 
                           RN => n11389, Q => n9067, QN => n_1145);
   clk_r_REG4160_S6 : DFFR_X1 port map( D => n9067, CK => clk, RN => n11402, Q 
                           => n9066, QN => n_1146);
   clk_r_REG4161_S7 : DFFR_X1 port map( D => n9066, CK => clk, RN => n11395, Q 
                           => n9065, QN => n_1147);
   clk_r_REG4250_S7 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_33_port, CK => clk, 
                           RN => n11403, Q => n9064, QN => n_1148);
   clk_r_REG4251_S8 : DFFR_X1 port map( D => n9064, CK => clk, RN => n11389, Q 
                           => n9063, QN => n_1149);
   clk_r_REG4252_S9 : DFFR_X1 port map( D => n9063, CK => clk, RN => n11397, Q 
                           => n9062, QN => n_1150);
   clk_r_REG4112_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_32_port, CK => clk, 
                           RN => n11379, Q => n9061, QN => n_1151);
   clk_r_REG4113_S6 : DFFR_X1 port map( D => n9061, CK => clk, RN => n11381, Q 
                           => n9060, QN => n_1152);
   clk_r_REG4114_S7 : DFFR_X1 port map( D => n9060, CK => clk, RN => n11389, Q 
                           => n9059, QN => n_1153);
   clk_r_REG4699_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_31_port, CK => clk, 
                           RN => n11386, Q => n9058, QN => n_1154);
   clk_r_REG4700_S12 : DFFR_X1 port map( D => n9058, CK => clk, RN => n11403, Q
                           => n9057, QN => n_1155);
   clk_r_REG4701_S13 : DFFR_X1 port map( D => n9057, CK => clk, RN => n11399, Q
                           => n9056, QN => n_1156);
   clk_r_REG4693_S17 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_30_port, CK => clk, 
                           RN => n11381, Q => n9055, QN => n_1157);
   clk_r_REG4694_S18 : DFFR_X1 port map( D => n9055, CK => clk, RN => n11395, Q
                           => n9054, QN => n_1158);
   clk_r_REG4695_S19 : DFFR_X1 port map( D => n9054, CK => clk, RN => n11394, Q
                           => n9053, QN => n_1159);
   clk_r_REG4687_S17 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_29_port, CK => clk, 
                           RN => n11387, Q => n9052, QN => n_1160);
   clk_r_REG4688_S18 : DFFR_X1 port map( D => n9052, CK => clk, RN => n11392, Q
                           => n9051, QN => n_1161);
   clk_r_REG4689_S19 : DFFR_X1 port map( D => n9051, CK => clk, RN => n11392, Q
                           => n9050, QN => n_1162);
   clk_r_REG3967_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_28_port, CK => clk, 
                           RN => n11382, Q => n9049, QN => n_1163);
   clk_r_REG3968_S6 : DFFR_X1 port map( D => n9049, CK => clk, RN => n11385, Q 
                           => n9048, QN => n_1164);
   clk_r_REG3969_S7 : DFFR_X1 port map( D => n9048, CK => clk, RN => n11398, Q 
                           => n9047, QN => n_1165);
   clk_r_REG3917_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_muxes_in_4_27_port, CK => clk, 
                           RN => n11384, Q => n9046, QN => n_1166);
   clk_r_REG3918_S6 : DFFR_X1 port map( D => n9046, CK => clk, RN => n11396, Q 
                           => n9045, QN => n_1167);
   clk_r_REG3919_S7 : DFFR_X1 port map( D => n9045, CK => clk, RN => n11386, Q 
                           => n9044, QN => n_1168);
   clk_r_REG4675_S17 : DFFR_X1 port map( D => data1_mul_15_port, CK => clk, RN 
                           => n11383, Q => n_1169, QN => n11302);
   clk_r_REG4676_S18 : DFFS_X1 port map( D => n11302, CK => clk, SN => n11397, 
                           Q => n11303, QN => n_1170);
   clk_r_REG4677_S19 : DFFS_X1 port map( D => n11303, CK => clk, SN => n11399, 
                           Q => n_1171, QN => n9041);
   clk_r_REG4475_S4 : DFFS_X1 port map( D => n11316, CK => clk, SN => n11378, Q
                           => n9040, QN => n_1172);
   clk_r_REG3625_S5 : DFFS_X1 port map( D => n1804, CK => clk, SN => n11395, Q 
                           => n9039, QN => n_1173);
   clk_r_REG6001_S5 : DFFR_X1 port map( D => n1803, CK => clk, RN => n11381, Q 
                           => n9038, QN => n_1174);
   clk_r_REG4472_S4 : DFFR_X1 port map( D => n11311, CK => clk, RN => n11385, Q
                           => n9037, QN => n_1175);
   clk_r_REG4464_S4 : DFFR_X1 port map( D => n11322, CK => clk, RN => n11392, Q
                           => n9036, QN => n_1176);
   clk_r_REG4466_S4 : DFFS_X1 port map( D => n11313, CK => clk, SN => n11398, Q
                           => n9035, QN => n_1177);
   clk_r_REG4487_S4 : DFFR_X1 port map( D => n7654, CK => clk, RN => n11399, Q 
                           => n9034, QN => n_1178);
   clk_r_REG4484_S4 : DFFS_X1 port map( D => n1834, CK => clk, SN => n11377, Q 
                           => n9033, QN => n_1179);
   clk_r_REG4342_S4 : DFFS_X1 port map( D => n11320, CK => clk, SN => n11401, Q
                           => n9032, QN => n_1180);
   clk_r_REG4360_S4 : DFFS_X1 port map( D => n11323, CK => clk, SN => n11385, Q
                           => n9031, QN => n13199);
   clk_r_REG4366_S4 : DFFS_X1 port map( D => n4506, CK => clk, SN => n11395, Q 
                           => n9030, QN => n13147);
   clk_r_REG4369_S4 : DFFS_X1 port map( D => n11314, CK => clk, SN => n11381, Q
                           => n9029, QN => n13171);
   clk_r_REG4451_S4 : DFFR_X1 port map( D => n1869, CK => clk, RN => n11384, Q 
                           => n9028, QN => n_1181);
   clk_r_REG4372_S4 : DFFS_X1 port map( D => n1874, CK => clk, SN => n11403, Q 
                           => n9027, QN => n13212);
   clk_r_REG4349_S4 : DFFR_X1 port map( D => n7659, CK => clk, RN => n11390, Q 
                           => n9026, QN => n13168);
   clk_r_REG4338_S4 : DFFR_X1 port map( D => n1871, CK => clk, RN => n11381, Q 
                           => n9025, QN => n_1182);
   clk_r_REG4358_S4 : DFFS_X1 port map( D => n1876, CK => clk, SN => n11402, Q 
                           => n9024, QN => n13189);
   clk_r_REG4455_S4 : DFFS_X1 port map( D => n11312, CK => clk, SN => n11380, Q
                           => n9023, QN => n13162);
   clk_r_REG4447_S4 : DFFS_X1 port map( D => n1866, CK => clk, SN => n11393, Q 
                           => n9022, QN => n13170);
   clk_r_REG4441_S4 : DFFS_X1 port map( D => n7759, CK => clk, SN => n11381, Q 
                           => n9021, QN => n_1183);
   clk_r_REG4442_S4 : DFFS_X1 port map( D => n7759, CK => clk, SN => n11396, Q 
                           => n9020, QN => n13146);
   clk_r_REG4444_S4 : DFFR_X1 port map( D => n4476, CK => clk, RN => n11399, Q 
                           => n9019, QN => n13195);
   clk_r_REG4456_S4 : DFFS_X1 port map( D => n11312, CK => clk, SN => n11378, Q
                           => n9018, QN => n_1184);
   clk_r_REG4437_S4 : DFFS_X1 port map( D => n1867, CK => clk, SN => n11401, Q 
                           => n9017, QN => n13190);
   clk_r_REG4459_S4 : DFFR_X1 port map( D => n1872, CK => clk, RN => n11402, Q 
                           => n9016, QN => n13208);
   clk_r_REG4423_S4 : DFFS_X1 port map( D => n13223, CK => clk, SN => n11378, Q
                           => n9015, QN => n_1185);
   clk_r_REG4404_S4 : DFFR_X1 port map( D => n13222, CK => clk, RN => n11386, Q
                           => n9014, QN => n_1186);
   clk_r_REG4418_S4 : DFFS_X1 port map( D => n1865, CK => clk, SN => n11399, Q 
                           => n9013, QN => n_1187);
   clk_r_REG4452_S4 : DFFS_X1 port map( D => n1869, CK => clk, SN => n11392, Q 
                           => n9012, QN => n_1188);
   clk_r_REG4364_S4 : DFFS_X1 port map( D => n1875, CK => clk, SN => n11378, Q 
                           => n9011, QN => n13185);
   clk_r_REG4344_S4 : DFFR_X1 port map( D => n1873, CK => clk, RN => n11385, Q 
                           => n9010, QN => n_1189);
   clk_r_REG4480_S4 : DFFS_X1 port map( D => n1833, CK => clk, SN => n11400, Q 
                           => n9009, QN => n13204);
   clk_r_REG4460_S4 : DFFR_X1 port map( D => n1870, CK => clk, RN => n11390, Q 
                           => n9008, QN => n_1190);
   clk_r_REG6653_S3 : DFFS_X1 port map( D => FUNC(3), CK => clk, SN => n11381, 
                           Q => n9007, QN => n_1191);
   clk_r_REG5585_S4 : DFFS_X1 port map( D => n9222, CK => clk, SN => n11387, Q 
                           => n9006, QN => n_1192);
   clk_r_REG4857_S4 : DFFS_X1 port map( D => DATA1(13), CK => clk, SN => n11378
                           , Q => n9005, QN => n_1193);
   clk_r_REG4671_S16 : DFFS_X1 port map( D => DATA1(16), CK => clk, SN => 
                           n11403, Q => n9004, QN => n_1194);
   clk_r_REG4662_S16 : DFFS_X1 port map( D => DATA1(18), CK => clk, SN => 
                           n11398, Q => n9003, QN => n_1195);
   clk_r_REG4631_S16 : DFFS_X1 port map( D => DATA1(27), CK => clk, SN => 
                           n11386, Q => n9002, QN => n_1196);
   clk_r_REG4612_S16 : DFFR_X1 port map( D => n1837, CK => clk, RN => n11380, Q
                           => n9001, QN => n_1197);
   clk_r_REG6654_S3 : DFFR_X1 port map( D => FUNC(3), CK => clk, RN => n11391, 
                           Q => n9000, QN => n_1198);
   clk_r_REG6650_S3 : DFFS_X1 port map( D => FUNC(2), CK => clk, SN => n11377, 
                           Q => n8999, QN => n_1199);
   clk_r_REG6822_S8 : DFFS_X1 port map( D => FUNC(1), CK => clk, SN => n11393, 
                           Q => n8998, QN => n_1200);
   clk_r_REG3834_S5 : DFFR_X1 port map( D => n4325, CK => clk, RN => n11389, Q 
                           => n8997, QN => n_1201);
   clk_r_REG3835_S6 : DFFR_X1 port map( D => n8997, CK => clk, RN => n11396, Q 
                           => n8996, QN => n_1202);
   clk_r_REG3836_S7 : DFFR_X1 port map( D => n8996, CK => clk, RN => n11397, Q 
                           => n8995, QN => n_1203);
   clk_r_REG3837_S8 : DFFR_X1 port map( D => n8995, CK => clk, RN => n11389, Q 
                           => n13182, QN => n11325);
   clk_r_REG3884_S5 : DFFR_X1 port map( D => n4319, CK => clk, RN => n11399, Q 
                           => n8993, QN => n_1204);
   clk_r_REG3885_S6 : DFFR_X1 port map( D => n8993, CK => clk, RN => n11392, Q 
                           => n8992, QN => n_1205);
   clk_r_REG3886_S7 : DFFR_X1 port map( D => n8992, CK => clk, RN => n11385, Q 
                           => n8991, QN => n_1206);
   clk_r_REG3887_S8 : DFFR_X1 port map( D => n8991, CK => clk, RN => n11383, Q 
                           => n8990, QN => n_1207);
   clk_r_REG3953_S5 : DFFR_X1 port map( D => n4316, CK => clk, RN => rst_BAR, Q
                           => n8989, QN => n_1208);
   clk_r_REG3954_S6 : DFFR_X1 port map( D => n8989, CK => clk, RN => n11383, Q 
                           => n8988, QN => n_1209);
   clk_r_REG3955_S7 : DFFR_X1 port map( D => n8988, CK => clk, RN => n11379, Q 
                           => n13175, QN => n11329);
   clk_r_REG3788_S5 : DFFR_X1 port map( D => n4310, CK => clk, RN => n11400, Q 
                           => n8986, QN => n_1210);
   clk_r_REG3789_S6 : DFFR_X1 port map( D => n8986, CK => clk, RN => n11385, Q 
                           => n8985, QN => n_1211);
   clk_r_REG3790_S7 : DFFR_X1 port map( D => n8985, CK => clk, RN => n11396, Q 
                           => n8984, QN => n_1212);
   clk_r_REG3859_S5 : DFFR_X1 port map( D => n4308, CK => clk, RN => n11396, Q 
                           => n8983, QN => n_1213);
   clk_r_REG3860_S6 : DFFR_X1 port map( D => n8983, CK => clk, RN => n11384, Q 
                           => n13174, QN => n11326);
   clk_r_REG3662_S5 : DFFR_X1 port map( D => n4303, CK => clk, RN => n11399, Q 
                           => n8981, QN => n_1214);
   clk_r_REG3663_S6 : DFFR_X1 port map( D => n8981, CK => clk, RN => n11397, Q 
                           => n8980, QN => n_1215);
   clk_r_REG4065_S5 : DFFR_X1 port map( D => n4302, CK => clk, RN => n11390, Q 
                           => n_1216, QN => n11328);
   clk_r_REG3535_S5 : DFFR_X1 port map( D => n4298, CK => clk, RN => n11377, Q 
                           => n8978, QN => n_1217);
   clk_r_REG4321_S5 : DFFR_X1 port map( D => n11331, CK => clk, RN => n11398, Q
                           => n_1218, QN => n8976);
   clk_r_REG4355_S4 : DFFR_X1 port map( D => n1870, CK => clk, RN => n11390, Q 
                           => n13183, QN => n8975);
   clk_r_REG4354_S4 : DFFS_X1 port map( D => n1870, CK => clk, SN => n11377, Q 
                           => n13156, QN => n8974);
   clk_r_REG4370_S4 : DFFS_X1 port map( D => n1874, CK => clk, SN => n11393, Q 
                           => n13165, QN => n8973);
   clk_r_REG4438_S4 : DFFS_X1 port map( D => n1868, CK => clk, SN => n11398, Q 
                           => n13192, QN => n8972);
   clk_r_REG3842_S5 : DFFR_X1 port map( D => n1808, CK => clk, RN => n11393, Q 
                           => n_1219, QN => n8971);
   clk_r_REG4477_S4 : DFFS_X1 port map( D => n1878, CK => clk, SN => n11384, Q 
                           => n_1220, QN => n8970);
   clk_r_REG4422_S4 : DFFR_X1 port map( D => n13223, CK => clk, RN => n11394, Q
                           => n_1221, QN => n8968);
   clk_r_REG4406_S4 : DFFR_X1 port map( D => n1865, CK => clk, RN => n11380, Q 
                           => n_1222, QN => n8967);
   clk_r_REG4405_S4 : DFFS_X1 port map( D => n1865, CK => clk, SN => n11380, Q 
                           => n_1223, QN => n8966);
   clk_r_REG4635_S5 : DFFR_X1 port map( D => n1802, CK => clk, RN => n11380, Q 
                           => n_1224, QN => n8965);
   clk_r_REG4654_S5 : DFFR_X1 port map( D => n1806, CK => clk, RN => n11389, Q 
                           => n_1225, QN => n8964);
   clk_r_REG3758_S5 : DFFR_X1 port map( D => n1805, CK => clk, RN => n11389, Q 
                           => n_1226, QN => n8963);
   clk_r_REG5999_S5 : DFFR_X1 port map( D => n1803, CK => clk, RN => n11383, Q 
                           => n_1227, QN => n8962);
   clk_r_REG5998_S5 : DFFS_X1 port map( D => n1803, CK => clk, SN => n11383, Q 
                           => n_1228, QN => n8961);
   clk_r_REG4389_S4 : DFFS_X1 port map( D => n13221, CK => clk, SN => n11384, Q
                           => n_1229, QN => n8960);
   clk_r_REG4147_S5 : DFFR_X1 port map( D => n4220, CK => clk, RN => n11390, Q 
                           => n8959, QN => n_1230);
   clk_r_REG4403_S4 : DFFS_X1 port map( D => n6338, CK => clk, SN => n11379, Q 
                           => n8958, QN => n_1231);
   clk_r_REG4333_S5 : DFFS_X1 port map( D => n6340, CK => clk, SN => n11386, Q 
                           => n8957, QN => n_1232);
   clk_r_REG4778_S5 : DFFS_X1 port map( D => n3892, CK => clk, SN => n11387, Q 
                           => n8956, QN => n_1233);
   clk_r_REG3680_S5 : DFFS_X1 port map( D => n4212, CK => clk, SN => n11400, Q 
                           => n8955, QN => n_1234);
   clk_r_REG3780_S4 : DFFR_X1 port map( D => n6502, CK => clk, RN => n11399, Q 
                           => n8954, QN => n_1235);
   clk_r_REG4435_S4 : DFFR_X1 port map( D => n6742, CK => clk, RN => n11391, Q 
                           => n8953, QN => n_1236);
   clk_r_REG3584_S5 : DFFS_X1 port map( D => n6749, CK => clk, SN => n11394, Q 
                           => n8952, QN => n_1237);
   clk_r_REG3681_S5 : DFFR_X1 port map( D => n6860, CK => clk, RN => n11382, Q 
                           => n8951, QN => n13210);
   clk_r_REG3576_S5 : DFFR_X1 port map( D => n6740, CK => clk, RN => n11392, Q 
                           => n8950, QN => n_1238);
   clk_r_REG4614_S4 : DFFS_X1 port map( D => n1836, CK => clk, SN => n11392, Q 
                           => n_1239, QN => n8949);
   clk_r_REG3682_S5 : DFFR_X1 port map( D => n6862, CK => clk, RN => n11378, Q 
                           => n_1240, QN => n13163);
   clk_r_REG3568_S5 : DFFR_X1 port map( D => n6876, CK => clk, RN => n11379, Q 
                           => n8947, QN => n_1241);
   clk_r_REG3773_S5 : DFFS_X1 port map( D => n6899, CK => clk, SN => n11392, Q 
                           => n8946, QN => n_1242);
   clk_r_REG3622_S5 : DFFS_X1 port map( D => n6908, CK => clk, SN => n11403, Q 
                           => n8945, QN => n_1243);
   clk_r_REG3807_S11 : DFFS_X1 port map( D => n6932, CK => clk, SN => n11398, Q
                           => n8944, QN => n_1244);
   clk_r_REG3847_S5 : DFFR_X1 port map( D => n7047, CK => clk, RN => n11388, Q 
                           => n8943, QN => n_1245);
   clk_r_REG3877_S4 : DFFR_X1 port map( D => n7086, CK => clk, RN => n11389, Q 
                           => n8942, QN => n_1246);
   clk_r_REG4084_S5 : DFFR_X1 port map( D => n4199, CK => clk, RN => n11387, Q 
                           => n8941, QN => n_1247);
   clk_r_REG3655_S14 : DFFS_X1 port map( D => n7153, CK => clk, SN => n11401, Q
                           => n8940, QN => n_1248);
   clk_r_REG4613_S4 : DFFS_X1 port map( D => n7325, CK => clk, SN => n11394, Q 
                           => n8939, QN => n_1249);
   clk_r_REG3593_S5 : DFFR_X1 port map( D => n4192, CK => clk, RN => n11388, Q 
                           => n8938, QN => n_1250);
   clk_r_REG3594_S6 : DFFR_X1 port map( D => n8938, CK => clk, RN => n11377, Q 
                           => n8937, QN => n_1251);
   clk_r_REG3595_S7 : DFFR_X1 port map( D => n8937, CK => clk, RN => n11394, Q 
                           => n8936, QN => n_1252);
   clk_r_REG3596_S8 : DFFR_X1 port map( D => n8936, CK => clk, RN => n11399, Q 
                           => n8935, QN => n_1253);
   clk_r_REG3597_S9 : DFFR_X1 port map( D => n8935, CK => clk, RN => n11397, Q 
                           => n8934, QN => n_1254);
   clk_r_REG3598_S10 : DFFR_X1 port map( D => n8934, CK => clk, RN => n11395, Q
                           => n8933, QN => n_1255);
   clk_r_REG3997_S5 : DFFS_X1 port map( D => n4055, CK => clk, SN => n11387, Q 
                           => n8932, QN => n_1256);
   clk_r_REG4132_S5 : DFFS_X1 port map( D => n11327, CK => clk, SN => n11380, Q
                           => n_1257, QN => n8930);
   clk_r_REG4134_S5 : DFFS_X1 port map( D => n7483, CK => clk, SN => n11399, Q 
                           => n8929, QN => n_1258);
   clk_r_REG4071_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_16_port, CK => clk, 
                           RN => n11385, Q => n8928, QN => n_1259);
   clk_r_REG4070_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_17_port, CK => clk, 
                           RN => n11382, Q => n8927, QN => n_1260);
   clk_r_REG4069_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_18_port, CK => clk, 
                           RN => n11386, Q => n8926, QN => n_1261);
   clk_r_REG4068_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_19_port, CK => clk, 
                           RN => n11381, Q => n8925, QN => n_1262);
   clk_r_REG4067_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_20_port, CK => clk, 
                           RN => n11398, Q => n8924, QN => n_1263);
   clk_r_REG3964_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_21_port, CK => clk, 
                           RN => n11390, Q => n8923, QN => n_1264);
   clk_r_REG3903_S5 : DFFR_X1 port map( D => n4186, CK => clk, RN => rst_BAR, Q
                           => n8922, QN => n_1265);
   clk_r_REG3904_S5 : DFFR_X1 port map( D => n4185, CK => clk, RN => n11378, Q 
                           => n8921, QN => n_1266);
   clk_r_REG3865_S7 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_23_port, CK => clk, 
                           RN => n11383, Q => n8920, QN => n_1267);
   clk_r_REG3864_S7 : DFFR_X1 port map( D => n4183, CK => clk, RN => n11389, Q 
                           => n8919, QN => n_1268);
   clk_r_REG3862_S7 : DFFR_X1 port map( D => n4182, CK => clk, RN => n11384, Q 
                           => n8918, QN => n_1269);
   clk_r_REG3801_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_25_port, CK => clk, 
                           RN => n11395, Q => n8917, QN => n_1270);
   clk_r_REG3800_S8 : DFFR_X1 port map( D => n4180, CK => clk, RN => n11389, Q 
                           => n8916, QN => n_1271);
   clk_r_REG3798_S8 : DFFR_X1 port map( D => n4179, CK => clk, RN => n11397, Q 
                           => n8915, QN => n_1272);
   clk_r_REG3841_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_27_port, CK => clk, 
                           RN => n11395, Q => n8914, QN => n_1273);
   clk_r_REG3840_S9 : DFFR_X1 port map( D => n4177, CK => clk, RN => n11384, Q 
                           => n8913, QN => n_1274);
   clk_r_REG3839_S9 : DFFR_X1 port map( D => n4176, CK => clk, RN => n11380, Q 
                           => n8912, QN => n_1275);
   clk_r_REG3838_S9 : DFFR_X1 port map( D => n4175, CK => clk, RN => n11380, Q 
                           => n8911, QN => n_1276);
   clk_r_REG4469_S4 : DFFR_X1 port map( D => n11324, CK => clk, RN => n11378, Q
                           => n_1277, QN => n8910);
   clk_r_REG4468_S4 : DFFS_X1 port map( D => n11324, CK => clk, SN => n11386, Q
                           => n_1278, QN => n8909);
   clk_r_REG4465_S4 : DFFS_X1 port map( D => n11313, CK => clk, SN => n11385, Q
                           => n_1279, QN => n8908);
   clk_r_REG4453_S4 : DFFS_X1 port map( D => n11312, CK => clk, SN => n11377, Q
                           => n13164, QN => n8906);
   clk_r_REG4359_S4 : DFFS_X1 port map( D => n11323, CK => clk, SN => n11402, Q
                           => n13148, QN => n8905);
   clk_r_REG4471_S4 : DFFR_X1 port map( D => n11311, CK => clk, RN => n11391, Q
                           => n_1280, QN => n8904);
   clk_r_REG3621_S5 : DFFS_X1 port map( D => n1804, CK => clk, SN => n11401, Q 
                           => n_1281, QN => n8903);
   clk_r_REG4479_S4 : DFFS_X1 port map( D => n1833, CK => clk, SN => n11400, Q 
                           => n13203, QN => n8902);
   clk_r_REG4630_S5 : DFFS_X1 port map( D => n4421, CK => clk, SN => n11400, Q 
                           => n8901, QN => n_1282);
   clk_r_REG4320_S5 : DFFS_X1 port map( D => n4111, CK => clk, SN => n11396, Q 
                           => n8900, QN => n_1283);
   clk_r_REG4462_S4 : DFFR_X1 port map( D => n11322, CK => clk, RN => n11377, Q
                           => n_1284, QN => n8899);
   clk_r_REG4461_S4 : DFFS_X1 port map( D => n11322, CK => clk, SN => n11401, Q
                           => n13181, QN => n8898);
   clk_r_REG4357_S4 : DFFS_X1 port map( D => n1876, CK => clk, SN => n11398, Q 
                           => n13184, QN => n8897);
   clk_r_REG4363_S4 : DFFS_X1 port map( D => n1875, CK => clk, SN => n11402, Q 
                           => n13159, QN => n8896);
   clk_r_REG4436_S4 : DFFS_X1 port map( D => n1867, CK => clk, SN => n11387, Q 
                           => n13151, QN => n8895);
   clk_r_REG4331_S5 : DFFS_X1 port map( D => n1429, CK => clk, SN => n11391, Q 
                           => n8894, QN => n_1285);
   clk_r_REG5915_S8 : DFFS_X1 port map( D => n1353, CK => clk, SN => n11400, Q 
                           => n8893, QN => n_1286);
   clk_r_REG4581_S4 : DFFR_X1 port map( D => n3862, CK => clk, RN => n11388, Q 
                           => n8892, QN => n_1287);
   clk_r_REG4421_S4 : DFFR_X1 port map( D => n13220, CK => clk, RN => n11391, Q
                           => n_1288, QN => n8891);
   clk_r_REG4420_S4 : DFFS_X1 port map( D => n13220, CK => clk, SN => n11378, Q
                           => n_1289, QN => n8890);
   clk_r_REG4402_S4 : DFFR_X1 port map( D => n13222, CK => clk, RN => n11388, Q
                           => n_1290, QN => n8889);
   clk_r_REG4319_S5 : DFFS_X1 port map( D => n2808, CK => clk, SN => n11392, Q 
                           => n8888, QN => n_1291);
   clk_r_REG4052_S5 : DFFR_X1 port map( D => n3933, CK => clk, RN => n11392, Q 
                           => n8887, QN => n_1292);
   clk_r_REG4705_S5 : DFFS_X1 port map( D => n7449, CK => clk, SN => n11391, Q 
                           => n8886, QN => n_1293);
   clk_r_REG3998_S6 : DFFR_X1 port map( D => n4274, CK => clk, RN => n11393, Q 
                           => n8885, QN => n_1294);
   clk_r_REG3999_S7 : DFFR_X1 port map( D => n8885, CK => clk, RN => n11399, Q 
                           => n8884, QN => n_1295);
   clk_r_REG4000_S8 : DFFR_X1 port map( D => n8884, CK => clk, RN => rst_BAR, Q
                           => n8883, QN => n_1296);
   clk_r_REG4001_S9 : DFFR_X1 port map( D => n8883, CK => clk, RN => n11388, Q 
                           => n8882, QN => n_1297);
   clk_r_REG4002_S10 : DFFR_X1 port map( D => n8882, CK => clk, RN => n11390, Q
                           => n8881, QN => n_1298);
   clk_r_REG4003_S11 : DFFS_X1 port map( D => n8881, CK => clk, SN => n11392, Q
                           => n8880, QN => n_1299);
   clk_r_REG3523_S6 : DFFR_X1 port map( D => n4270, CK => clk, RN => n11392, Q 
                           => n8879, QN => n_1300);
   clk_r_REG3524_S7 : DFFR_X1 port map( D => n8879, CK => clk, RN => n11399, Q 
                           => n8878, QN => n_1301);
   clk_r_REG3525_S8 : DFFR_X1 port map( D => n8878, CK => clk, RN => rst_BAR, Q
                           => n8877, QN => n_1302);
   clk_r_REG3526_S9 : DFFR_X1 port map( D => n8877, CK => clk, RN => n11391, Q 
                           => n8876, QN => n_1303);
   clk_r_REG3527_S10 : DFFR_X1 port map( D => n8876, CK => clk, RN => n11384, Q
                           => n8875, QN => n_1304);
   clk_r_REG3651_S10 : DFFR_X1 port map( D => n4266, CK => clk, RN => n11379, Q
                           => n8874, QN => n_1305);
   clk_r_REG3652_S11 : DFFR_X1 port map( D => n8874, CK => clk, RN => n11396, Q
                           => n8873, QN => n_1306);
   clk_r_REG3653_S12 : DFFR_X1 port map( D => n8873, CK => clk, RN => n11388, Q
                           => n8872, QN => n_1307);
   clk_r_REG3654_S13 : DFFR_X1 port map( D => n8872, CK => clk, RN => n11393, Q
                           => n8871, QN => n_1308);
   clk_r_REG4074_S8 : DFFR_X1 port map( D => n4263, CK => clk, RN => n11386, Q 
                           => n8870, QN => n_1309);
   clk_r_REG4075_S9 : DFFR_X1 port map( D => n8870, CK => clk, RN => n11390, Q 
                           => n8869, QN => n_1310);
   clk_r_REG4076_S10 : DFFR_X1 port map( D => n8869, CK => clk, RN => n11385, Q
                           => n8868, QN => n_1311);
   clk_r_REG4077_S11 : DFFS_X1 port map( D => n8868, CK => clk, SN => n11402, Q
                           => n8867, QN => n_1312);
   clk_r_REG4920_S5 : DFFR_X1 port map( D => n4257, CK => clk, RN => n11383, Q 
                           => n8866, QN => n_1313);
   clk_r_REG4921_S6 : DFFR_X1 port map( D => n8866, CK => clk, RN => n11387, Q 
                           => n8865, QN => n_1314);
   clk_r_REG4922_S7 : DFFR_X1 port map( D => n8865, CK => clk, RN => n11381, Q 
                           => n8864, QN => n_1315);
   clk_r_REG4923_S8 : DFFR_X1 port map( D => n8864, CK => clk, RN => n11395, Q 
                           => n8863, QN => n_1316);
   clk_r_REG4924_S9 : DFFR_X1 port map( D => n8863, CK => clk, RN => n11391, Q 
                           => n8862, QN => n_1317);
   clk_r_REG4925_S10 : DFFR_X1 port map( D => n8862, CK => clk, RN => n11396, Q
                           => n8861, QN => n_1318);
   clk_r_REG3975_S4 : DFFR_X1 port map( D => n1852, CK => clk, RN => n11395, Q 
                           => n_1319, QN => n8860);
   clk_r_REG4092_S4 : DFFS_X1 port map( D => n3918, CK => clk, SN => n11388, Q 
                           => n8859, QN => n_1320);
   clk_r_REG3781_S4 : DFFS_X1 port map( D => n6184, CK => clk, SN => n11377, Q 
                           => n13160, QN => n11337);
   clk_r_REG4044_S16 : DFFS_X1 port map( D => n6206, CK => clk, SN => n11402, Q
                           => n8857, QN => n_1321);
   clk_r_REG4415_S4 : DFFR_X1 port map( D => n1849, CK => clk, RN => n11390, Q 
                           => n_1322, QN => n8856);
   clk_r_REG4253_S4 : DFFS_X1 port map( D => n3910, CK => clk, SN => n11401, Q 
                           => n_1323, QN => n13214);
   clk_r_REG4449_S4 : DFFR_X1 port map( D => n1869, CK => clk, RN => n11393, Q 
                           => n_1324, QN => n8854);
   clk_r_REG4448_S4 : DFFS_X1 port map( D => n1869, CK => clk, SN => n11400, Q 
                           => n_1325, QN => n8853);
   clk_r_REG4377_S4 : DFFR_X1 port map( D => n11315, CK => clk, RN => n11383, Q
                           => n_1326, QN => n8852);
   clk_r_REG4376_S4 : DFFS_X1 port map( D => n11315, CK => clk, SN => n11402, Q
                           => n_1327, QN => n8851);
   clk_r_REG3930_S4 : DFFR_X1 port map( D => n6561, CK => clk, RN => n11397, Q 
                           => n8850, QN => n_1328);
   clk_r_REG4117_S4 : DFFS_X1 port map( D => n7114, CK => clk, SN => n11394, Q 
                           => n8849, QN => n13197);
   clk_r_REG3559_S5 : DFFS_X1 port map( D => n6869, CK => clk, SN => n11381, Q 
                           => n8848, QN => n_1329);
   clk_r_REG3632_S5 : DFFS_X1 port map( D => n6850, CK => clk, SN => n11377, Q 
                           => n8847, QN => n_1330);
   clk_r_REG3577_S5 : DFFS_X1 port map( D => n6733, CK => clk, SN => n11402, Q 
                           => n8846, QN => n_1331);
   clk_r_REG3567_S5 : DFFR_X1 port map( D => n6870, CK => clk, RN => n11381, Q 
                           => n8845, QN => n_1332);
   clk_r_REG3569_S5 : DFFS_X1 port map( D => n6858, CK => clk, SN => n11401, Q 
                           => n8844, QN => n_1333);
   clk_r_REG3624_S5 : DFFR_X1 port map( D => n6739, CK => clk, RN => n11385, Q 
                           => n8843, QN => n_1334);
   clk_r_REG6322_S4 : DFFR_X1 port map( D => n4078, CK => clk, RN => n11391, Q 
                           => n8842, QN => n_1335);
   clk_r_REG3691_S4 : DFFR_X1 port map( D => n6874, CK => clk, RN => n11385, Q 
                           => n8841, QN => n_1336);
   clk_r_REG3671_S11 : DFFS_X1 port map( D => n6871, CK => clk, SN => n11381, Q
                           => n8840, QN => n_1337);
   clk_r_REG3550_S5 : DFFR_X1 port map( D => n6888, CK => clk, RN => n11402, Q 
                           => n8839, QN => n_1338);
   clk_r_REG3774_S4 : DFFS_X1 port map( D => n3866, CK => clk, SN => n11400, Q 
                           => n8838, QN => n_1339);
   clk_r_REG3549_S5 : DFFS_X1 port map( D => n4075, CK => clk, SN => n11403, Q 
                           => n8837, QN => n_1340);
   clk_r_REG3623_S5 : DFFR_X1 port map( D => n6905, CK => clk, RN => n11395, Q 
                           => n8836, QN => n_1341);
   clk_r_REG3706_S4 : DFFR_X1 port map( D => n4074, CK => clk, RN => n11379, Q 
                           => n8835, QN => n_1342);
   clk_r_REG3705_S4 : DFFS_X1 port map( D => n4073, CK => clk, SN => n11383, Q 
                           => n8834, QN => n_1343);
   clk_r_REG3845_S5 : DFFR_X1 port map( D => n6957, CK => clk, RN => n11402, Q 
                           => n8833, QN => n_1344);
   clk_r_REG4434_S4 : DFFR_X1 port map( D => n4070, CK => clk, RN => n11403, Q 
                           => n8832, QN => n_1345);
   clk_r_REG4430_S4 : DFFS_X1 port map( D => n4069, CK => clk, SN => n11382, Q 
                           => n8831, QN => n_1346);
   clk_r_REG4658_S4 : DFFS_X1 port map( D => n4068, CK => clk, SN => n11402, Q 
                           => n8830, QN => n_1347);
   clk_r_REG5511_S4 : DFFR_X1 port map( D => n4067, CK => clk, RN => n11382, Q 
                           => n8829, QN => n_1348);
   clk_r_REG4666_S4 : DFFS_X1 port map( D => n3844, CK => clk, SN => n11401, Q 
                           => n8828, QN => n_1349);
   clk_r_REG6066_S4 : DFFR_X1 port map( D => n4066, CK => clk, RN => n11394, Q 
                           => n8827, QN => n_1350);
   clk_r_REG3888_S5 : DFFR_X1 port map( D => n4065, CK => clk, RN => n11381, Q 
                           => n8826, QN => n_1351);
   clk_r_REG3875_S9 : DFFR_X1 port map( D => n4200, CK => clk, RN => n11392, Q 
                           => n8825, QN => n_1352);
   clk_r_REG3876_S10 : DFFR_X1 port map( D => n8825, CK => clk, RN => n11382, Q
                           => n8824, QN => n_1353);
   clk_r_REG3958_S5 : DFFS_X1 port map( D => n3838, CK => clk, SN => n11398, Q 
                           => n8823, QN => n_1354);
   clk_r_REG3959_S4 : DFFR_X1 port map( D => n4064, CK => clk, RN => n11395, Q 
                           => n8822, QN => n_1355);
   clk_r_REG3957_S5 : DFFR_X1 port map( D => n4063, CK => clk, RN => n11387, Q 
                           => n8821, QN => n_1356);
   clk_r_REG4091_S5 : DFFS_X1 port map( D => n4061, CK => clk, SN => n11393, Q 
                           => n8820, QN => n_1357);
   clk_r_REG4086_S5 : DFFR_X1 port map( D => n7150, CK => clk, RN => n11386, Q 
                           => n8819, QN => n_1358);
   clk_r_REG4433_S4 : DFFS_X1 port map( D => n4060, CK => clk, SN => n11391, Q 
                           => n8818, QN => n_1359);
   clk_r_REG4606_S16 : DFFS_X1 port map( D => n7333, CK => clk, SN => n11402, Q
                           => n8817, QN => n_1360);
   clk_r_REG3637_S4 : DFFS_X1 port map( D => n7332, CK => clk, SN => n11379, Q 
                           => n8816, QN => n_1361);
   clk_r_REG3636_S4 : DFFS_X1 port map( D => n7339, CK => clk, SN => n11401, Q 
                           => n8815, QN => n_1362);
   clk_r_REG4142_S5 : DFFS_X1 port map( D => n7481, CK => clk, SN => n11397, Q 
                           => n8814, QN => n_1363);
   clk_r_REG4105_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_3_18_port, CK => clk, 
                           RN => n11379, Q => n8813, QN => n_1364);
   clk_r_REG3962_S5 : DFFR_X1 port map( D => n4190, CK => clk, RN => n11381, Q 
                           => n8812, QN => n_1365);
   clk_r_REG3898_S5 : DFFR_X1 port map( D => n4189, CK => clk, RN => n11390, Q 
                           => n8811, QN => n_1366);
   clk_r_REG3901_S6 : DFFR_X1 port map( D => n4188, CK => clk, RN => n11379, Q 
                           => n8810, QN => n_1367);
   clk_r_REG4373_S4 : DFFS_X1 port map( D => n11318, CK => clk, SN => n11378, Q
                           => n13142, QN => n8809);
   clk_r_REG4474_S4 : DFFS_X1 port map( D => n11316, CK => clk, SN => n11403, Q
                           => n13206, QN => n8808);
   clk_r_REG4340_S4 : DFFS_X1 port map( D => n11320, CK => clk, SN => n11397, Q
                           => n13150, QN => n8807);
   clk_r_REG4445_S4 : DFFS_X1 port map( D => n1866, CK => clk, SN => n11399, Q 
                           => n13139, QN => n8806);
   clk_r_REG4329_S4 : DFFS_X1 port map( D => n11317, CK => clk, SN => n11398, Q
                           => n_1368, QN => n8805);
   clk_r_REG4346_S4 : DFFR_X1 port map( D => n11319, CK => clk, RN => n11391, Q
                           => n_1369, QN => n8804);
   clk_r_REG3983_S5 : DFFS_X1 port map( D => n11330, CK => clk, SN => n11394, Q
                           => n_1370, QN => n8803);
   clk_r_REG4335_S4 : DFFR_X1 port map( D => n1877, CK => clk, RN => n11388, Q 
                           => n_1371, QN => n8802);
   clk_r_REG4343_S4 : DFFR_X1 port map( D => n1873, CK => clk, RN => n11388, Q 
                           => n13166, QN => n8801);
   clk_r_REG4777_S5 : DFFR_X1 port map( D => n4216, CK => clk, RN => n11387, Q 
                           => n8800, QN => n_1372);
   clk_r_REG3566_S5 : DFFR_X1 port map( D => n1800, CK => clk, RN => n11395, Q 
                           => n_1373, QN => n8799);
   clk_r_REG4770_S5 : DFFR_X1 port map( D => n4048, CK => clk, RN => n11396, Q 
                           => n8798, QN => n_1374);
   clk_r_REG4771_S6 : DFFR_X1 port map( D => n8798, CK => clk, RN => n11388, Q 
                           => n8797, QN => n_1375);
   clk_r_REG4772_S7 : DFFR_X1 port map( D => n8797, CK => clk, RN => n11381, Q 
                           => n8796, QN => n_1376);
   clk_r_REG4773_S8 : DFFR_X1 port map( D => n8796, CK => clk, RN => n11389, Q 
                           => n8795, QN => n_1377);
   clk_r_REG4774_S9 : DFFR_X1 port map( D => n8795, CK => clk, RN => n11398, Q 
                           => n8794, QN => n_1378);
   clk_r_REG4775_S10 : DFFR_X1 port map( D => n8794, CK => clk, RN => n11390, Q
                           => n8793, QN => n_1379);
   clk_r_REG4491_S5 : DFFR_X1 port map( D => n4046, CK => clk, RN => n11379, Q 
                           => n8792, QN => n_1380);
   clk_r_REG4492_S5 : DFFR_X1 port map( D => n4045, CK => clk, RN => n11398, Q 
                           => n8791, QN => n_1381);
   clk_r_REG4152_S5 : DFFR_X1 port map( D => n4044, CK => clk, RN => n11381, Q 
                           => n8790, QN => n_1382);
   clk_r_REG4151_S5 : DFFR_X1 port map( D => n4043, CK => clk, RN => n11399, Q 
                           => n8789, QN => n_1383);
   clk_r_REG4098_S5 : DFFR_X1 port map( D => n4042, CK => clk, RN => n11389, Q 
                           => n8788, QN => n_1384);
   clk_r_REG4096_S5 : DFFR_X1 port map( D => n4041, CK => clk, RN => n11387, Q 
                           => n8787, QN => n_1385);
   clk_r_REG4097_S5 : DFFR_X1 port map( D => n4040, CK => clk, RN => n11396, Q 
                           => n8786, QN => n_1386);
   clk_r_REG4095_S5 : DFFR_X1 port map( D => n4039, CK => clk, RN => n11385, Q 
                           => n8785, QN => n_1387);
   clk_r_REG3940_S5 : DFFR_X1 port map( D => n4038, CK => clk, RN => n11396, Q 
                           => n8784, QN => n_1388);
   clk_r_REG3899_S5 : DFFR_X1 port map( D => n4037, CK => clk, RN => n11398, Q 
                           => n8783, QN => n_1389);
   clk_r_REG3895_S5 : DFFR_X1 port map( D => n4036, CK => clk, RN => n11388, Q 
                           => n8782, QN => n_1390);
   clk_r_REG3600_S5 : DFFR_X1 port map( D => n4035, CK => clk, RN => n11383, Q 
                           => n8781, QN => n_1391);
   clk_r_REG3719_S5 : DFFR_X1 port map( D => n4034, CK => clk, RN => n11399, Q 
                           => n8780, QN => n_1392);
   clk_r_REG3907_S5 : DFFR_X1 port map( D => n4033, CK => clk, RN => n11398, Q 
                           => n8779, QN => n_1393);
   clk_r_REG3908_S6 : DFFR_X1 port map( D => n8779, CK => clk, RN => n11389, Q 
                           => n8778, QN => n_1394);
   clk_r_REG3985_S6 : DFFR_X1 port map( D => n4027, CK => clk, RN => n11396, Q 
                           => n8777, QN => n_1395);
   clk_r_REG3986_S7 : DFFR_X1 port map( D => n8777, CK => clk, RN => n11393, Q 
                           => n8776, QN => n_1396);
   clk_r_REG3987_S8 : DFFR_X1 port map( D => n8776, CK => clk, RN => n11386, Q 
                           => n8775, QN => n_1397);
   clk_r_REG3988_S9 : DFFR_X1 port map( D => n8775, CK => clk, RN => n11378, Q 
                           => n8774, QN => n_1398);
   clk_r_REG3989_S10 : DFFR_X1 port map( D => n8774, CK => clk, RN => n11391, Q
                           => n8773, QN => n_1399);
   clk_r_REG3891_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CK => clk, 
                           RN => rst_BAR, Q => n8772, QN => n_1400);
   clk_r_REG3893_S6 : DFFR_X1 port map( D => n4026, CK => clk, RN => n11382, Q 
                           => n8771, QN => n_1401);
   clk_r_REG3894_S6 : DFFR_X1 port map( D => n4025, CK => clk, RN => n11403, Q 
                           => n8770, QN => n_1402);
   clk_r_REG4135_S6 : DFFR_X1 port map( D => n4020, CK => clk, RN => n11397, Q 
                           => n8769, QN => n_1403);
   clk_r_REG4136_S7 : DFFR_X1 port map( D => n8769, CK => clk, RN => n11391, Q 
                           => n8768, QN => n_1404);
   clk_r_REG4137_S8 : DFFR_X1 port map( D => n8768, CK => clk, RN => n11393, Q 
                           => n8767, QN => n_1405);
   clk_r_REG4138_S9 : DFFR_X1 port map( D => n8767, CK => clk, RN => n11386, Q 
                           => n8766, QN => n_1406);
   clk_r_REG4139_S10 : DFFR_X1 port map( D => n8766, CK => clk, RN => n11383, Q
                           => n8765, QN => n_1407);
   clk_r_REG3601_S6 : DFFR_X1 port map( D => n4011, CK => clk, RN => n11386, Q 
                           => n8764, QN => n_1408);
   clk_r_REG3720_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CK => clk, RN => n11391, Q => n8763, QN => n_1409);
   clk_r_REG3721_S6 : DFFR_X1 port map( D => n4010, CK => clk, RN => n11402, Q 
                           => n8762, QN => n_1410);
   clk_r_REG4053_S6 : DFFR_X1 port map( D => n4003, CK => clk, RN => n11385, Q 
                           => n8761, QN => n_1411);
   clk_r_REG4054_S7 : DFFR_X1 port map( D => n8761, CK => clk, RN => n11385, Q 
                           => n8760, QN => n_1412);
   clk_r_REG4055_S8 : DFFR_X1 port map( D => n8760, CK => clk, RN => n11386, Q 
                           => n8759, QN => n_1413);
   clk_r_REG4056_S9 : DFFR_X1 port map( D => n8759, CK => clk, RN => rst_BAR, Q
                           => n8758, QN => n_1414);
   clk_r_REG4057_S10 : DFFR_X1 port map( D => n8758, CK => clk, RN => n11382, Q
                           => n8757, QN => n_1415);
   clk_r_REG3650_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_10_port, CK => clk, 
                           RN => n11379, Q => n_1416, QN => n11333);
   clk_r_REG4078_S9 : DFFR_X1 port map( D => n4001, CK => clk, RN => n11387, Q 
                           => n8755, QN => n_1417);
   clk_r_REG4072_S6 : DFFR_X1 port map( D => n4000, CK => clk, RN => n11380, Q 
                           => n8754, QN => n_1418);
   clk_r_REG3941_S6 : DFFR_X1 port map( D => n3999, CK => clk, RN => n11398, Q 
                           => n8753, QN => n_1419);
   clk_r_REG3900_S6 : DFFR_X1 port map( D => n3998, CK => clk, RN => n11384, Q 
                           => n8752, QN => n_1420);
   clk_r_REG3896_S6 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CK => clk, RN => n11389, Q => n8751, QN => n_1421);
   clk_r_REG3897_S6 : DFFR_X1 port map( D => n3997, CK => clk, RN => n11384, Q 
                           => n8750, QN => n_1422);
   clk_r_REG3892_S7 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CK => clk, 
                           RN => n11395, Q => n8749, QN => n_1423);
   clk_r_REG3537_S7 : DFFR_X1 port map( D => n3989, CK => clk, RN => n11390, Q 
                           => n8748, QN => n_1424);
   clk_r_REG4079_S10 : DFFR_X1 port map( D => n3986, CK => clk, RN => rst_BAR, 
                           Q => n8747, QN => n_1425);
   clk_r_REG4080_S11 : DFFR_X1 port map( D => n8747, CK => clk, RN => n11394, Q
                           => n8746, QN => n_1426);
   clk_r_REG4081_S12 : DFFR_X1 port map( D => n8746, CK => clk, RN => n11403, Q
                           => n8745, QN => n_1427);
   clk_r_REG4082_S13 : DFFR_X1 port map( D => n8745, CK => clk, RN => n11391, Q
                           => n8744, QN => n_1428);
   clk_r_REG4073_S7 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_12_port, CK => clk, 
                           RN => n11399, Q => n_1429, QN => n11334);
   clk_r_REG3942_S7 : DFFR_X1 port map( D => n3984, CK => clk, RN => n11394, Q 
                           => n8742, QN => n_1430);
   clk_r_REG3873_S7 : DFFR_X1 port map( D => n3983, CK => clk, RN => n11380, Q 
                           => n8741, QN => n_1431);
   clk_r_REG3872_S7 : DFFR_X1 port map( D => n3982, CK => clk, RN => n11377, Q 
                           => n8740, QN => n_1432);
   clk_r_REG3602_S7 : DFFR_X1 port map( D => n3981, CK => clk, RN => n11383, Q 
                           => n8739, QN => n_1433);
   clk_r_REG3722_S7 : DFFR_X1 port map( D => n3980, CK => clk, RN => n11393, Q 
                           => n8738, QN => n_1434);
   clk_r_REG3871_S7 : DFFR_X1 port map( D => n3979, CK => clk, RN => n11385, Q 
                           => n8737, QN => n_1435);
   clk_r_REG3870_S7 : DFFR_X1 port map( D => n3978, CK => clk, RN => n11392, Q 
                           => n8736, QN => n_1436);
   clk_r_REG3869_S7 : DFFR_X1 port map( D => n3977, CK => clk, RN => n11383, Q 
                           => n8735, QN => n_1437);
   clk_r_REG3868_S7 : DFFR_X1 port map( D => n3976, CK => clk, RN => n11390, Q 
                           => n8734, QN => n_1438);
   clk_r_REG3866_S7 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CK => clk, RN => n11398, Q => n8733, QN => n_1439);
   clk_r_REG3867_S7 : DFFR_X1 port map( D => n3975, CK => clk, RN => n11389, Q 
                           => n8732, QN => n_1440);
   clk_r_REG3863_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CK => clk, 
                           RN => n11400, Q => n8731, QN => n_1441);
   clk_r_REG3665_S8 : DFFR_X1 port map( D => n3972, CK => clk, RN => n11395, Q 
                           => n8730, QN => n_1442);
   clk_r_REG3943_S8 : DFFR_X1 port map( D => n3970, CK => clk, RN => n11382, Q 
                           => n8729, QN => n_1443);
   clk_r_REG3944_S9 : DFFR_X1 port map( D => n8729, CK => clk, RN => n11385, Q 
                           => n8728, QN => n_1444);
   clk_r_REG3945_S10 : DFFR_X1 port map( D => n8728, CK => clk, RN => n11388, Q
                           => n8727, QN => n_1445);
   clk_r_REG3874_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_14_port, CK => clk, 
                           RN => n11396, Q => n_1446, QN => n11340);
   clk_r_REG3824_S8 : DFFR_X1 port map( D => n3968, CK => clk, RN => n11391, Q 
                           => n8725, QN => n_1447);
   clk_r_REG3603_S8 : DFFR_X1 port map( D => n3967, CK => clk, RN => n11383, Q 
                           => n8724, QN => n_1448);
   clk_r_REG3723_S8 : DFFR_X1 port map( D => n3966, CK => clk, RN => n11393, Q 
                           => n8723, QN => n_1449);
   clk_r_REG3823_S8 : DFFR_X1 port map( D => n3965, CK => clk, RN => n11398, Q 
                           => n8722, QN => n_1450);
   clk_r_REG3819_S8 : DFFR_X1 port map( D => n3964, CK => clk, RN => n11394, Q 
                           => n8721, QN => n_1451);
   clk_r_REG3815_S8 : DFFR_X1 port map( D => n3963, CK => clk, RN => n11397, Q 
                           => n8720, QN => n_1452);
   clk_r_REG3812_S8 : DFFR_X1 port map( D => n3962, CK => clk, RN => n11380, Q 
                           => n8719, QN => n_1453);
   clk_r_REG3808_S8 : DFFR_X1 port map( D => n3961, CK => clk, RN => n11396, Q 
                           => n8718, QN => n_1454);
   clk_r_REG3804_S8 : DFFR_X1 port map( D => n3960, CK => clk, RN => n11389, Q 
                           => n8717, QN => n_1455);
   clk_r_REG3538_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CK => clk, RN => n11389, Q => n8716, QN => n_1456);
   clk_r_REG3539_S8 : DFFR_X1 port map( D => n3959, CK => clk, RN => n11398, Q 
                           => n8715, QN => n_1457);
   clk_r_REG3799_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CK => clk, 
                           RN => n11401, Q => n8714, QN => n_1458);
   clk_r_REG3792_S9 : DFFR_X1 port map( D => n3956, CK => clk, RN => n11400, Q 
                           => n8713, QN => n_1459);
   clk_r_REG3825_S9 : DFFR_X1 port map( D => n3954, CK => clk, RN => n11384, Q 
                           => n8712, QN => n_1460);
   clk_r_REG3826_S10 : DFFR_X1 port map( D => n8712, CK => clk, RN => n11384, Q
                           => n8711, QN => n_1461);
   clk_r_REG3827_S11 : DFFS_X1 port map( D => n8711, CK => clk, SN => n11399, Q
                           => n8710, QN => n_1462);
   clk_r_REG3604_S9 : DFFR_X1 port map( D => n3953, CK => clk, RN => n11394, Q 
                           => n8709, QN => n_1463);
   clk_r_REG3605_S10 : DFFR_X1 port map( D => n8709, CK => clk, RN => n11402, Q
                           => n8708, QN => n_1464);
   clk_r_REG3724_S9 : DFFR_X1 port map( D => n3952, CK => clk, RN => n11387, Q 
                           => n8707, QN => n_1465);
   clk_r_REG3725_S10 : DFFR_X1 port map( D => n8707, CK => clk, RN => n11384, Q
                           => n8706, QN => n_1466);
   clk_r_REG3727_S9 : DFFR_X1 port map( D => n3951, CK => clk, RN => n11382, Q 
                           => n8705, QN => n_1467);
   clk_r_REG3728_S10 : DFFR_X1 port map( D => n8705, CK => clk, RN => n11383, Q
                           => n8704, QN => n_1468);
   clk_r_REG3820_S9 : DFFR_X1 port map( D => n3950, CK => clk, RN => n11389, Q 
                           => n8703, QN => n_1469);
   clk_r_REG3821_S10 : DFFR_X1 port map( D => n8703, CK => clk, RN => n11381, Q
                           => n8702, QN => n_1470);
   clk_r_REG3816_S9 : DFFR_X1 port map( D => n3949, CK => clk, RN => n11393, Q 
                           => n8701, QN => n_1471);
   clk_r_REG3817_S10 : DFFR_X1 port map( D => n8701, CK => clk, RN => n11379, Q
                           => n8700, QN => n_1472);
   clk_r_REG3813_S9 : DFFR_X1 port map( D => n3948, CK => clk, RN => n11393, Q 
                           => n8699, QN => n_1473);
   clk_r_REG3814_S10 : DFFR_X1 port map( D => n8699, CK => clk, RN => n11396, Q
                           => n8698, QN => n_1474);
   clk_r_REG3809_S9 : DFFR_X1 port map( D => n3947, CK => clk, RN => n11386, Q 
                           => n8697, QN => n_1475);
   clk_r_REG3810_S10 : DFFR_X1 port map( D => n8697, CK => clk, RN => n11391, Q
                           => n8696, QN => n_1476);
   clk_r_REG3805_S9 : DFFR_X1 port map( D => n3945, CK => clk, RN => n11397, Q 
                           => n8695, QN => n_1477);
   clk_r_REG3806_S10 : DFFR_X1 port map( D => n8695, CK => clk, RN => n11384, Q
                           => n8694, QN => n_1478);
   clk_r_REG3540_S9 : DFFR_X1 port map( D => n3944, CK => clk, RN => n11387, Q 
                           => n8693, QN => n_1479);
   clk_r_REG3541_S10 : DFFR_X1 port map( D => n8693, CK => clk, RN => n11394, Q
                           => n8692, QN => n_1480);
   clk_r_REG3802_S9 : DFFR_X1 port map( D => n3943, CK => clk, RN => n11382, Q 
                           => n8691, QN => n_1481);
   clk_r_REG3803_S10 : DFFR_X1 port map( D => n8691, CK => clk, RN => n11403, Q
                           => n8690, QN => n_1482);
   clk_r_REG3666_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CK => clk, RN => n11388, Q => n8689, QN => n_1483);
   clk_r_REG3667_S9 : DFFR_X1 port map( D => n3941, CK => clk, RN => n11390, Q 
                           => n8688, QN => n_1484);
   clk_r_REG3668_S10 : DFFR_X1 port map( D => n8688, CK => clk, RN => n11403, Q
                           => n8687, QN => n_1485);
   clk_r_REG3669_S11 : DFFR_X1 port map( D => n8687, CK => clk, RN => n11380, Q
                           => n8686, QN => n_1486);
   clk_r_REG3670_S10 : DFFR_X1 port map( D => n3938, CK => clk, RN => n11395, Q
                           => n8685, QN => n_1487);
   clk_r_REG3672_S10 : DFFR_X1 port map( D => n3937, CK => clk, RN => n11392, Q
                           => n8684, QN => n_1488);
   clk_r_REG3673_S11 : DFFR_X1 port map( D => n8684, CK => clk, RN => n11387, Q
                           => n8683, QN => n_1489);
   clk_r_REG3793_S10 : DFFR_X1 port map( D => n3936, CK => clk, RN => n11400, Q
                           => n8682, QN => n_1490);
   clk_r_REG3794_S10 : DFFR_X1 port map( D => n3935, CK => clk, RN => n11393, Q
                           => n8681, QN => n_1491);
   clk_r_REG3796_S10 : DFFR_X1 port map( D => n3934, CK => clk, RN => n11397, Q
                           => n8680, QN => n_1492);
   clk_r_REG3797_S11 : DFFS_X1 port map( D => n8680, CK => clk, SN => n11383, Q
                           => n8679, QN => n_1493);
   clk_r_REG4352_S4 : DFFR_X1 port map( D => n11321, CK => clk, RN => rst_BAR, 
                           Q => n13178, QN => n8678);
   clk_r_REG4351_S4 : DFFS_X1 port map( D => n11321, CK => clk, SN => n11380, Q
                           => n13202, QN => n8677);
   clk_r_REG4457_S4 : DFFR_X1 port map( D => n1872, CK => clk, RN => n11381, Q 
                           => n_1494, QN => n8676);
   clk_r_REG4058_S4 : DFFS_X1 port map( D => n3932, CK => clk, SN => n11400, Q 
                           => n8675, QN => n_1495);
   clk_r_REG4090_S5 : DFFR_X1 port map( D => n3920, CK => clk, RN => n11381, Q 
                           => n8674, QN => n_1496);
   clk_r_REG4089_S5 : DFFR_X1 port map( D => n3919, CK => clk, RN => n11402, Q 
                           => n8673, QN => n_1497);
   clk_r_REG4431_S4 : DFFR_X1 port map( D => n6880, CK => clk, RN => n11398, Q 
                           => n8672, QN => n_1498);
   clk_r_REG4429_S4 : DFFS_X1 port map( D => n6179, CK => clk, SN => n11403, Q 
                           => n8671, QN => n_1499);
   clk_r_REG4401_S4 : DFFS_X1 port map( D => n6174, CK => clk, SN => n11378, Q 
                           => n8670, QN => n_1500);
   clk_r_REG4387_S4 : DFFR_X1 port map( D => n6177, CK => clk, RN => n11388, Q 
                           => n8669, QN => n_1501);
   clk_r_REG3690_S4 : DFFS_X1 port map( D => n6881, CK => clk, SN => n11403, Q 
                           => n8668, QN => n_1502);
   clk_r_REG4386_S4 : DFFR_X1 port map( D => n6192, CK => clk, RN => n11382, Q 
                           => n8667, QN => n_1503);
   clk_r_REG4412_S16 : DFFR_X1 port map( D => n6191, CK => clk, RN => n11391, Q
                           => n8666, QN => n_1504);
   clk_r_REG4383_S4 : DFFR_X1 port map( D => n6197, CK => clk, RN => n11401, Q 
                           => n8665, QN => n_1505);
   clk_r_REG3712_S4 : DFFR_X1 port map( D => n6196, CK => clk, RN => n11395, Q 
                           => n8664, QN => n_1506);
   clk_r_REG4396_S4 : DFFS_X1 port map( D => n6205, CK => clk, SN => n11380, Q 
                           => n8663, QN => n_1507);
   clk_r_REG4380_S4 : DFFS_X1 port map( D => n6204, CK => clk, SN => n11377, Q 
                           => n8662, QN => n_1508);
   clk_r_REG4391_S4 : DFFR_X1 port map( D => n6208, CK => clk, RN => n11385, Q 
                           => n8661, QN => n_1509);
   clk_r_REG4045_S16 : DFFR_X1 port map( D => n6207, CK => clk, RN => n11394, Q
                           => n8660, QN => n_1510);
   clk_r_REG4379_S4 : DFFS_X1 port map( D => n6213, CK => clk, SN => n11400, Q 
                           => n8659, QN => n_1511);
   clk_r_REG4395_S4 : DFFS_X1 port map( D => n6212, CK => clk, SN => n11395, Q 
                           => n8658, QN => n_1512);
   clk_r_REG4388_S4 : DFFR_X1 port map( D => n6215, CK => clk, RN => n11379, Q 
                           => n8657, QN => n_1513);
   clk_r_REG4399_S4 : DFFS_X1 port map( D => n6214, CK => clk, SN => n11387, Q 
                           => n8656, QN => n_1514);
   clk_r_REG4394_S4 : DFFS_X1 port map( D => n6238, CK => clk, SN => n11397, Q 
                           => n8655, QN => n_1515);
   clk_r_REG4381_S4 : DFFS_X1 port map( D => n6237, CK => clk, SN => n11401, Q 
                           => n8654, QN => n_1516);
   clk_r_REG4393_S4 : DFFS_X1 port map( D => n6241, CK => clk, SN => n11400, Q 
                           => n8653, QN => n_1517);
   clk_r_REG4378_S4 : DFFS_X1 port map( D => n6240, CK => clk, SN => n11395, Q 
                           => n8652, QN => n_1518);
   clk_r_REG4168_S4 : DFFR_X1 port map( D => n6261, CK => clk, RN => n11393, Q 
                           => n8651, QN => n_1519);
   clk_r_REG4165_S4 : DFFR_X1 port map( D => n6260, CK => clk, RN => n11386, Q 
                           => n8650, QN => n_1520);
   clk_r_REG3528_S11 : DFFS_X1 port map( D => n3911, CK => clk, SN => n11396, Q
                           => n8649, QN => n_1521);
   clk_r_REG4145_S5 : DFFR_X1 port map( D => n6267, CK => clk, RN => n11397, Q 
                           => n8648, QN => n_1522);
   clk_r_REG4125_S4 : DFFR_X1 port map( D => n6381, CK => clk, RN => n11382, Q 
                           => n8647, QN => n_1523);
   clk_r_REG4148_S5 : DFFS_X1 port map( D => n6314, CK => clk, SN => n11381, Q 
                           => n8646, QN => n_1524);
   clk_r_REG4167_S4 : DFFR_X1 port map( D => n6294, CK => clk, RN => n11393, Q 
                           => n8645, QN => n_1525);
   clk_r_REG3976_S4 : DFFS_X1 port map( D => n6422, CK => clk, SN => n11398, Q 
                           => n8644, QN => n13188);
   clk_r_REG4334_S5 : DFFS_X1 port map( D => n3905, CK => clk, SN => n11399, Q 
                           => n8643, QN => n_1526);
   clk_r_REG5914_S8 : DFFR_X1 port map( D => n3904, CK => clk, RN => n11385, Q 
                           => n8642, QN => n_1527);
   clk_r_REG4121_S4 : DFFR_X1 port map( D => n1854, CK => clk, RN => n11386, Q 
                           => n_1528, QN => n8641);
   clk_r_REG4409_S4 : DFFS_X1 port map( D => n3902, CK => clk, SN => n11393, Q 
                           => n8640, QN => n_1529);
   clk_r_REG3990_S4 : DFFS_X1 port map( D => n3900, CK => clk, SN => n11395, Q 
                           => n8639, QN => n_1530);
   clk_r_REG4332_S5 : DFFS_X1 port map( D => n6367, CK => clk, SN => n11396, Q 
                           => n8638, QN => n_1531);
   clk_r_REG4120_S4 : DFFS_X1 port map( D => n6980, CK => clk, SN => n11403, Q 
                           => n8637, QN => n13187);
   clk_r_REG4780_S5 : DFFS_X1 port map( D => n3897, CK => clk, SN => n11377, Q 
                           => n8636, QN => n_1532);
   clk_r_REG4328_S4 : DFFS_X1 port map( D => n3896, CK => clk, SN => n11377, Q 
                           => n8635, QN => n_1533);
   clk_r_REG4779_S5 : DFFR_X1 port map( D => n3895, CK => clk, RN => n11390, Q 
                           => n8634, QN => n_1534);
   clk_r_REG3932_S4 : DFFS_X1 port map( D => n1858, CK => clk, SN => n11379, Q 
                           => n13158, QN => n8633);
   clk_r_REG4428_S4 : DFFS_X1 port map( D => n3894, CK => clk, SN => n11378, Q 
                           => n8632, QN => n_1535);
   clk_r_REG4776_S4 : DFFS_X1 port map( D => n3893, CK => clk, SN => n11395, Q 
                           => n8631, QN => n_1536);
   clk_r_REG4119_S4 : DFFR_X1 port map( D => n7287, CK => clk, RN => n11389, Q 
                           => n8630, QN => n13198);
   clk_r_REG4384_S4 : DFFS_X1 port map( D => n3888, CK => clk, SN => n11393, Q 
                           => n8629, QN => n_1537);
   clk_r_REG4385_S4 : DFFS_X1 port map( D => n3885, CK => clk, SN => n11378, Q 
                           => n8628, QN => n_1538);
   clk_r_REG3687_S4 : DFFR_X1 port map( D => n11335, CK => clk, RN => rst_BAR, 
                           Q => n_1539, QN => n8627);
   clk_r_REG4478_S4 : DFFS_X1 port map( D => n4205, CK => clk, SN => n11403, Q 
                           => n8626, QN => n_1540);
   clk_r_REG3931_S4 : DFFR_X1 port map( D => n6533, CK => clk, RN => n11386, Q 
                           => n_1541, QN => n11339);
   clk_r_REG3970_S4 : DFFS_X1 port map( D => n6523, CK => clk, SN => n11388, Q 
                           => n_1542, QN => n11338);
   clk_r_REG4398_S4 : DFFS_X1 port map( D => n6505, CK => clk, SN => n11377, Q 
                           => n8623, QN => n_1543);
   clk_r_REG3765_S4 : DFFR_X1 port map( D => n6506, CK => clk, RN => n11380, Q 
                           => n8622, QN => n_1544);
   clk_r_REG3710_S4 : DFFR_X1 port map( D => n6510, CK => clk, RN => n11393, Q 
                           => n8621, QN => n_1545);
   clk_r_REG3763_S4 : DFFS_X1 port map( D => n6517, CK => clk, SN => n11396, Q 
                           => n8620, QN => n_1546);
   clk_r_REG4390_S4 : DFFS_X1 port map( D => n6525, CK => clk, SN => n11382, Q 
                           => n8619, QN => n_1547);
   clk_r_REG3929_S4 : DFFR_X1 port map( D => n6524, CK => clk, RN => n11384, Q 
                           => n8618, QN => n_1548);
   clk_r_REG3971_S4 : DFFR_X1 port map( D => n6530, CK => clk, RN => n11380, Q 
                           => n8617, QN => n_1549);
   clk_r_REG3928_S4 : DFFR_X1 port map( D => n6529, CK => clk, RN => n11396, Q 
                           => n8616, QN => n_1550);
   clk_r_REG3689_S4 : DFFS_X1 port map( D => n6677, CK => clk, SN => n11377, Q 
                           => n8615, QN => n_1551);
   clk_r_REG3762_S4 : DFFS_X1 port map( D => n6541, CK => clk, SN => n11401, Q 
                           => n8614, QN => n_1552);
   clk_r_REG3926_S4 : DFFS_X1 port map( D => n1850, CK => clk, SN => n11385, Q 
                           => n13186, QN => n8613);
   clk_r_REG3925_S4 : DFFS_X1 port map( D => n6618, CK => clk, SN => n11395, Q 
                           => n8612, QN => n_1553);
   clk_r_REG4432_S4 : DFFS_X1 port map( D => n6675, CK => clk, SN => n11380, Q 
                           => n8611, QN => n_1554);
   clk_r_REG3923_S4 : DFFS_X1 port map( D => n1851, CK => clk, SN => n11402, Q 
                           => n13194, QN => n8610);
   clk_r_REG3920_S4 : DFFR_X1 port map( D => n1855, CK => clk, RN => n11385, Q 
                           => n_1555, QN => n8609);
   clk_r_REG3973_S4 : DFFR_X1 port map( D => n1856, CK => clk, RN => n11381, Q 
                           => n_1556, QN => n8608);
   clk_r_REG3921_S4 : DFFS_X1 port map( D => n6617, CK => clk, SN => n11401, Q 
                           => n8607, QN => n_1557);
   clk_r_REG4118_S4 : DFFR_X1 port map( D => n7097, CK => clk, RN => n11381, Q 
                           => n8606, QN => n13154);
   clk_r_REG4426_S4 : DFFS_X1 port map( D => n6676, CK => clk, SN => n11382, Q 
                           => n8605, QN => n_1558);
   clk_r_REG4116_S4 : DFFS_X1 port map( D => n7134, CK => clk, SN => n11400, Q 
                           => n8604, QN => n_1559);
   clk_r_REG4115_S4 : DFFR_X1 port map( D => n6763, CK => clk, RN => n11379, Q 
                           => n8603, QN => n_1560);
   clk_r_REG4166_S4 : DFFR_X1 port map( D => n6762, CK => clk, RN => n11390, Q 
                           => n8602, QN => n_1561);
   clk_r_REG3795_S11 : DFFR_X1 port map( D => n6793, CK => clk, RN => n11392, Q
                           => n8601, QN => n_1562);
   clk_r_REG4427_S4 : DFFS_X1 port map( D => n3875, CK => clk, SN => n11385, Q 
                           => n8600, QN => n_1563);
   clk_r_REG4926_S4 : DFFS_X1 port map( D => n6837, CK => clk, SN => n11395, Q 
                           => n8599, QN => n_1564);
   clk_r_REG4123_S4 : DFFR_X1 port map( D => n7284, CK => clk, RN => n11382, Q 
                           => n8598, QN => n13200);
   clk_r_REG3634_S4 : DFFS_X1 port map( D => n1838, CK => clk, SN => n11403, Q 
                           => n_1565, QN => n8597);
   clk_r_REG3635_S4 : DFFS_X1 port map( D => n6853, CK => clk, SN => n11402, Q 
                           => n8596, QN => n_1566);
   clk_r_REG3638_S4 : DFFS_X1 port map( D => n6852, CK => clk, SN => n11401, Q 
                           => n8595, QN => n_1567);
   clk_r_REG3683_S4 : DFFR_X1 port map( D => n6865, CK => clk, RN => n11384, Q 
                           => n8594, QN => n_1568);
   clk_r_REG3558_S5 : DFFR_X1 port map( D => n6889, CK => clk, RN => n11392, Q 
                           => n8593, QN => n_1569);
   clk_r_REG3775_S4 : DFFS_X1 port map( D => n3867, CK => clk, SN => n11382, Q 
                           => n_1570, QN => n13215);
   clk_r_REG3772_S5 : DFFR_X1 port map( D => n6896, CK => clk, RN => n11386, Q 
                           => n8591, QN => n_1571);
   clk_r_REG3542_S11 : DFFS_X1 port map( D => n3865, CK => clk, SN => n11397, Q
                           => n_1572, QN => n13216);
   clk_r_REG3698_S5 : DFFS_X1 port map( D => n3863, CK => clk, SN => n11397, Q 
                           => n8589, QN => n_1573);
   clk_r_REG3811_S11 : DFFS_X1 port map( D => n3861, CK => clk, SN => n11402, Q
                           => n8588, QN => n_1574);
   clk_r_REG3757_S5 : DFFR_X1 port map( D => n6935, CK => clk, RN => n11384, Q 
                           => n8587, QN => n_1575);
   clk_r_REG3844_S5 : DFFS_X1 port map( D => n3860, CK => clk, SN => n11382, Q 
                           => n8586, QN => n_1576);
   clk_r_REG3759_S4 : DFFS_X1 port map( D => n3859, CK => clk, SN => n11385, Q 
                           => n_1577, QN => n13217);
   clk_r_REG3750_S5 : DFFR_X1 port map( D => n6949, CK => clk, RN => n11396, Q 
                           => n8584, QN => n_1578);
   clk_r_REG3743_S5 : DFFS_X1 port map( D => n3858, CK => clk, SN => n11384, Q 
                           => n8583, QN => n_1579);
   clk_r_REG3818_S11 : DFFS_X1 port map( D => n3856, CK => clk, SN => n11383, Q
                           => n8582, QN => n_1580);
   clk_r_REG5129_S4 : DFFS_X1 port map( D => n3854, CK => clk, SN => n11377, Q 
                           => n8581, QN => n_1581);
   clk_r_REG4162_S4 : DFFR_X1 port map( D => n7286, CK => clk, RN => n11402, Q 
                           => n8580, QN => n_1582);
   clk_r_REG3822_S11 : DFFS_X1 port map( D => n3851, CK => clk, SN => n11394, Q
                           => n8579, QN => n_1583);
   clk_r_REG3736_S5 : DFFR_X1 port map( D => n7007, CK => clk, RN => n11380, Q 
                           => n8578, QN => n_1584);
   clk_r_REG3843_S5 : DFFR_X1 port map( D => n3850, CK => clk, RN => n11387, Q 
                           => n8577, QN => n_1585);
   clk_r_REG3729_S11 : DFFS_X1 port map( D => n3849, CK => clk, SN => n11393, Q
                           => n8576, QN => n_1586);
   clk_r_REG3846_S5 : DFFS_X1 port map( D => n3848, CK => clk, SN => n11400, Q 
                           => n8575, QN => n_1587);
   clk_r_REG3726_S11 : DFFS_X1 port map( D => n3847, CK => clk, SN => n11377, Q
                           => n8574, QN => n_1588);
   clk_r_REG3620_S5 : DFFR_X1 port map( D => n3846, CK => clk, RN => rst_BAR, Q
                           => n8573, QN => n_1589);
   clk_r_REG3613_S5 : DFFR_X1 port map( D => n3845, CK => clk, RN => n11387, Q 
                           => n8572, QN => n_1590);
   clk_r_REG3606_S11 : DFFS_X1 port map( D => n3843, CK => clk, SN => n11388, Q
                           => n8571, QN => n_1591);
   clk_r_REG3849_S5 : DFFR_X1 port map( D => n3842, CK => clk, RN => n11394, Q 
                           => n8570, QN => n_1592);
   clk_r_REG3946_S4 : DFFS_X1 port map( D => n3837, CK => clk, SN => n11400, Q 
                           => n_1593, QN => n13219);
   clk_r_REG4085_S5 : DFFR_X1 port map( D => n3836, CK => clk, RN => n11386, Q 
                           => n_1594, QN => n13213);
   clk_r_REG3852_S4 : DFFS_X1 port map( D => n4062, CK => clk, SN => n11380, Q 
                           => n8567, QN => n_1595);
   clk_r_REG4083_S5 : DFFR_X1 port map( D => n3834, CK => clk, RN => n11387, Q 
                           => n8566, QN => n_1596);
   clk_r_REG3599_S11 : DFFS_X1 port map( D => n3831, CK => clk, SN => n11397, Q
                           => n8565, QN => n_1597);
   clk_r_REG4163_S4 : DFFR_X1 port map( D => n7285, CK => clk, RN => n11396, Q 
                           => n8564, QN => n_1598);
   clk_r_REG3684_S4 : DFFR_X1 port map( D => n7326, CK => clk, RN => n11395, Q 
                           => n8563, QN => n_1599);
   clk_r_REG3586_S4 : DFFR_X1 port map( D => n7340, CK => clk, RN => n11394, Q 
                           => n8562, QN => n_1600);
   clk_r_REG4337_S4 : DFFR_X1 port map( D => n1871, CK => clk, RN => n11391, Q 
                           => n13155, QN => n8561);
   clk_r_REG3709_S4 : DFFR_X1 port map( D => n1840, CK => clk, RN => n11400, Q 
                           => n_1601, QN => n8560);
   clk_r_REG4323_S6 : DFFR_X1 port map( D => n4280, CK => clk, RN => n11390, Q 
                           => n8559, QN => n_1602);
   clk_r_REG4324_S7 : DFFR_X1 port map( D => n8559, CK => clk, RN => rst_BAR, Q
                           => n8558, QN => n_1603);
   clk_r_REG4325_S8 : DFFR_X1 port map( D => n8558, CK => clk, RN => n11391, Q 
                           => n8557, QN => n_1604);
   clk_r_REG4326_S9 : DFFR_X1 port map( D => n8557, CK => clk, RN => n11397, Q 
                           => n8556, QN => n_1605);
   clk_r_REG4327_S10 : DFFR_X1 port map( D => n8556, CK => clk, RN => n11393, Q
                           => n8555, QN => n_1606);
   clk_r_REG4611_S16 : DFFR_X1 port map( D => n6744, CK => clk, RN => n11392, Q
                           => n8554, QN => n_1607);
   clk_r_REG5582_S5 : DFFS_X1 port map( D => n3822, CK => clk, SN => n11401, Q 
                           => n8553, QN => n_1608);
   clk_r_REG3848_S5 : DFFS_X1 port map( D => n3821, CK => clk, SN => n11379, Q 
                           => n_1609, QN => n13218);
   clk_r_REG4088_S5 : DFFS_X1 port map( D => n3835, CK => clk, SN => n11403, Q 
                           => n8551, QN => n_1610);
   clk_r_REG4087_S5 : DFFR_X1 port map( D => n3820, CK => clk, RN => n11379, Q 
                           => n8550, QN => n_1611);
   clk_r_REG3536_S6 : DFFR_X1 port map( D => n4184, CK => clk, RN => n11378, Q 
                           => n8549, QN => n_1612);
   clk_r_REG3664_S7 : DFFR_X1 port map( D => n4181, CK => clk, RN => n11392, Q 
                           => n8548, QN => n_1613);
   clk_r_REG3791_S8 : DFFR_X1 port map( D => n4178, CK => clk, RN => n11383, Q 
                           => n8547, QN => n_1614);
   clk_r_REG4414_S4 : DFFS_X1 port map( D => n6198, CK => clk, SN => n11380, Q 
                           => n8546, QN => n_1615);
   clk_r_REG4410_S4 : DFFR_X1 port map( D => n6187, CK => clk, RN => n11378, Q 
                           => n8545, QN => n_1616);
   clk_r_REG4411_S4 : DFFR_X1 port map( D => n6938, CK => clk, RN => n11384, Q 
                           => n8544, QN => n13191);
   clk_r_REG3711_S4 : DFFS_X1 port map( D => n1845, CK => clk, SN => n11378, Q 
                           => n_1617, QN => n8543);
   clk_r_REG4124_S4 : DFFR_X1 port map( D => n6351, CK => clk, RN => n11396, Q 
                           => n8542, QN => n_1618);
   clk_r_REG4419_S4 : DFFR_X1 port map( D => n1853, CK => clk, RN => n11391, Q 
                           => n_1619, QN => n8541);
   clk_r_REG4413_S4 : DFFS_X1 port map( D => n1830, CK => clk, SN => n11403, Q 
                           => n_1620, QN => n8540);
   clk_r_REG4164_S4 : DFFR_X1 port map( D => n6268, CK => clk, RN => rst_BAR, Q
                           => n8539, QN => n_1621);
   clk_r_REG4417_S4 : DFFS_X1 port map( D => n6516, CK => clk, SN => n11389, Q 
                           => n8538, QN => n_1622);
   clk_r_REG3778_S4 : DFFS_X1 port map( D => n1842, CK => clk, SN => n11390, Q 
                           => n_1623, QN => n8537);
   clk_r_REG3688_S4 : DFFR_X1 port map( D => n6671, CK => clk, RN => n11382, Q 
                           => n13176, QN => n11304);
   clk_r_REG3910_S5 : DFFR_X1 port map( D => n3800, CK => clk, RN => n11389, Q 
                           => n8535, QN => n_1624);
   clk_r_REG3909_S6 : DFFR_X1 port map( D => n4187, CK => clk, RN => n11392, Q 
                           => n8534, QN => n_1625);
   clk_r_REG5576_S5 : DFFR_X1 port map( D => n3794, CK => clk, RN => n11390, Q 
                           => n8533, QN => n_1626);
   clk_r_REG5577_S6 : DFFR_X1 port map( D => n8533, CK => clk, RN => n11397, Q 
                           => n8532, QN => n_1627);
   clk_r_REG5578_S7 : DFFR_X1 port map( D => n8532, CK => clk, RN => n11386, Q 
                           => n8531, QN => n_1628);
   clk_r_REG5579_S8 : DFFR_X1 port map( D => n8531, CK => clk, RN => n11395, Q 
                           => n8530, QN => n_1629);
   clk_r_REG5580_S9 : DFFR_X1 port map( D => n8530, CK => clk, RN => n11395, Q 
                           => n8529, QN => n_1630);
   clk_r_REG5581_S10 : DFFR_X1 port map( D => n8529, CK => clk, RN => n11388, Q
                           => n8528, QN => n_1631);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n554, Q => n4395);
   clk_r_REG4482_S4 : DFFS_X1 port map( D => n1834, CK => clk, SN => n11394, Q 
                           => n13205, QN => n8969);
   clk_r_REG3522_S5 : DFFS_X1 port map( D => n7485, CK => clk, SN => n11394, Q 
                           => n8931, QN => n_1632);
   clk_r_REG4143_S5 : DFFS_X1 port map( D => n11305, CK => clk, SN => n11394, Q
                           => n_1633, QN => n8977);
   clk_r_REG4367_S4 : DFFS_X1 port map( D => n11314, CK => clk, SN => n11397, Q
                           => n_1634, QN => n8907);
   U3 : CLKBUF_X1 port map( A => n11378, Z => n11377);
   U4 : CLKBUF_X1 port map( A => rst_BAR, Z => n11378);
   U5 : CLKBUF_X1 port map( A => n11403, Z => n11379);
   U6 : CLKBUF_X1 port map( A => n11403, Z => n11380);
   U7 : CLKBUF_X1 port map( A => n11402, Z => n11381);
   U8 : CLKBUF_X1 port map( A => n11402, Z => n11382);
   U9 : CLKBUF_X1 port map( A => n11402, Z => n11383);
   U10 : CLKBUF_X1 port map( A => n11401, Z => n11384);
   U11 : CLKBUF_X1 port map( A => n11401, Z => n11385);
   U12 : CLKBUF_X1 port map( A => n11401, Z => n11386);
   U13 : CLKBUF_X1 port map( A => n11400, Z => n11387);
   U14 : CLKBUF_X1 port map( A => n11400, Z => n11388);
   U15 : CLKBUF_X1 port map( A => n11400, Z => n11389);
   U16 : CLKBUF_X1 port map( A => n11382, Z => n11390);
   U17 : CLKBUF_X1 port map( A => n11399, Z => n11391);
   U18 : CLKBUF_X1 port map( A => n11399, Z => n11392);
   U19 : CLKBUF_X1 port map( A => n11383, Z => n11393);
   U20 : CLKBUF_X1 port map( A => n11386, Z => n11394);
   U21 : CLKBUF_X1 port map( A => n11386, Z => n11395);
   U22 : CLKBUF_X1 port map( A => n11399, Z => n11396);
   U23 : CLKBUF_X1 port map( A => n11382, Z => n11397);
   U24 : CLKBUF_X1 port map( A => n11400, Z => n11398);
   U25 : CLKBUF_X1 port map( A => n11384, Z => n11399);
   U26 : CLKBUF_X1 port map( A => n11377, Z => n11400);
   U27 : CLKBUF_X1 port map( A => n11377, Z => n11401);
   U28 : CLKBUF_X1 port map( A => n11377, Z => n11402);
   U29 : CLKBUF_X1 port map( A => n11377, Z => n11403);
   U30 : INV_X2 port map( A => n12341, ZN => n12541);
   U31 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , A2 => n12790, ZN => n12819);
   U32 : NOR2_X2 port map( A1 => n13174, A2 => n12930, ZN => n12959);
   U33 : NOR2_X2 port map( A1 => n13175, A2 => n12969, ZN => n12998);
   U34 : NOR2_X2 port map( A1 => n11325, A2 => n13007, ZN => n13041);
   U35 : NOR2_X2 port map( A1 => n11328, A2 => n12891, ZN => n12924);
   U36 : NOR2_X2 port map( A1 => n13182, A2 => n13007, ZN => n13040);
   U37 : NOR2_X2 port map( A1 => n11326, A2 => n12930, ZN => n12963);
   U38 : NOR2_X2 port map( A1 => n11329, A2 => n12969, ZN => n13002);
   U39 : NOR2_X2 port map( A1 => n12790, A2 => n12823, ZN => n12825);
   U40 : NOR2_X2 port map( A1 => n12890, A2 => n11328, ZN => n12925);
   U41 : NOR3_X4 port map( A1 => n13121, A2 => n13092, A3 => n11553, ZN => 
                           n13123);
   U42 : OAI21_X2 port map( B1 => n13078, B2 => n13088, A => n13072, ZN => 
                           n13121);
   U43 : NOR3_X4 port map( A1 => n11325, A2 => n11309, A3 => n8990, ZN => 
                           n13042);
   U44 : INV_X2 port map( A => n11917, ZN => n11895);
   U45 : OR2_X1 port map( A1 => n11532, A2 => n11781, ZN => n12237);
   U46 : NOR2_X1 port map( A1 => DATA2(3), A2 => n1870, ZN => n11553);
   U47 : NAND2_X1 port map( A1 => n11553, A2 => n13077, ZN => n11917);
   U48 : INV_X1 port map( A => n12163, ZN => n12332);
   U49 : NOR2_X1 port map( A1 => n1835, A2 => FUNC(3), ZN => n12518);
   U50 : INV_X1 port map( A => n13220, ZN => n11781);
   U51 : AOI21_X1 port map( B1 => n13082, B2 => n11553, A => n13220, ZN => 
                           n13108);
   U52 : INV_X1 port map( A => data1_mul_0_port, ZN => n1826);
   U53 : INV_X1 port map( A => data1_mul_15_port, ZN => n1810);
   U54 : INV_X1 port map( A => n12545, ZN => n12216);
   U55 : INV_X1 port map( A => n554, ZN => n12756);
   U56 : CLKBUF_X1 port map( A => n12786, Z => n12781);
   U57 : INV_X1 port map( A => n11906, ZN => n1865);
   U58 : INV_X1 port map( A => n13133, ZN => n1872);
   U59 : AOI211_X1 port map( C1 => n12541, C2 => n11544, A => n11543, B => 
                           n7822, ZN => n6095);
   U60 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n4295, ZN => n11404);
   U61 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, B2 
                           => n4295, A => n11404, ZN => n7449);
   U62 : INV_X1 port map( A => n7769, ZN => n1827);
   U63 : INV_X1 port map( A => n7449, ZN => n13070);
   U64 : NAND2_X1 port map( A1 => n13070, A2 => n1827, ZN => n11327);
   U65 : OR2_X1 port map( A1 => n7769, A2 => n11404, ZN => n7481);
   U66 : AND2_X1 port map( A1 => n11327, A2 => n7481, ZN => n7483);
   U67 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_2_4_port, ZN => 
                           n1821);
   U68 : XOR2_X1 port map( A => n1810, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => n1809);
   U69 : INV_X1 port map( A => DATA2(3), ZN => n13078);
   U70 : NOR2_X1 port map( A1 => DATA2(5), A2 => DATA2(4), ZN => n13099);
   U71 : NOR2_X1 port map( A1 => n13078, A2 => n13099, ZN => n13096);
   U72 : INV_X1 port map( A => n13096, ZN => n1874);
   U73 : INV_X1 port map( A => n13099, ZN => n1870);
   U74 : INV_X1 port map( A => DATA2(1), ZN => n13088);
   U75 : INV_X1 port map( A => DATA2(0), ZN => n13082);
   U76 : NOR2_X1 port map( A1 => n13088, A2 => n13082, ZN => n13091);
   U77 : INV_X1 port map( A => n13091, ZN => n13075);
   U78 : NOR2_X1 port map( A1 => n13078, A2 => n13075, ZN => n13073);
   U79 : AOI21_X1 port map( B1 => DATA2(2), B2 => n13073, A => n1870, ZN => 
                           n1875);
   U80 : INV_X1 port map( A => n1875, ZN => n4506);
   U81 : NOR2_X1 port map( A1 => DATA2(2), A2 => n1870, ZN => n13074);
   U82 : OR2_X1 port map( A1 => n11553, A2 => n13074, ZN => n13072);
   U83 : AOI21_X1 port map( B1 => n13088, B2 => n13099, A => n13072, ZN => 
                           n1867);
   U84 : INV_X1 port map( A => DATA2(2), ZN => n13077);
   U85 : NOR2_X1 port map( A1 => n13077, A2 => n13082, ZN => n11532);
   U86 : AND2_X1 port map( A1 => DATA2(3), A2 => n11532, ZN => n11644);
   U87 : NOR3_X1 port map( A1 => n13072, A2 => n1867, A3 => n11644, ZN => 
                           n11927);
   U88 : INV_X1 port map( A => n11927, ZN => n1866);
   U89 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n12409);
   U90 : OAI21_X1 port map( B1 => DATA1(16), B2 => DATA2_I_16_port, A => n12409
                           , ZN => n1807);
   U91 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n11650);
   U92 : INV_X1 port map( A => FUNC(2), ZN => n11536);
   U93 : NAND2_X1 port map( A1 => n11650, A2 => n11536, ZN => n554);
   U94 : INV_X1 port map( A => n12756, ZN => n13225);
   U95 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n11736)
                           ;
   U96 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n11736, 
                           ZN => n1429);
   U97 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n11738)
                           ;
   U98 : OAI21_X1 port map( B1 => DATA1(6), B2 => DATA2_I_6_port, A => n11738, 
                           ZN => n1353);
   U99 : XOR2_X1 port map( A => DATA2_I_15_port, B => DATA1(15), Z => n12442);
   U100 : XOR2_X1 port map( A => DATA2_I_7_port, B => DATA1(7), Z => n11743);
   U101 : INV_X1 port map( A => DATA1(5), ZN => n11764);
   U102 : XOR2_X1 port map( A => n11764, B => DATA2_I_5_port, Z => n11769);
   U103 : INV_X1 port map( A => n11769, ZN => n11772);
   U104 : XOR2_X1 port map( A => DATA2_I_3_port, B => n9225, Z => n11732);
   U105 : NAND2_X1 port map( A1 => n9223, A2 => DATA2_I_2_port, ZN => n11730);
   U106 : OAI21_X1 port map( B1 => n9223, B2 => DATA2_I_2_port, A => n11730, ZN
                           => n12171);
   U107 : NAND2_X1 port map( A1 => DATA2_I_1_port, A2 => n9222, ZN => n11733);
   U108 : NAND2_X1 port map( A1 => n9221, A2 => DATA2_I_0_port, ZN => n12334);
   U109 : INV_X1 port map( A => n12334, ZN => n12532);
   U110 : NOR2_X1 port map( A1 => n9221, A2 => DATA2_I_0_port, ZN => n12531);
   U111 : OAI21_X1 port map( B1 => DATA2_I_1_port, B2 => n9222, A => n11733, ZN
                           => n12333);
   U112 : NOR2_X1 port map( A1 => n12531, A2 => n12333, ZN => n12328);
   U113 : OAI21_X1 port map( B1 => n12532, B2 => n9220, A => n12328, ZN => 
                           n11405);
   U114 : OAI221_X1 port map( B1 => n12171, B2 => n11733, C1 => n12171, C2 => 
                           n11405, A => n11730, ZN => n11406);
   U115 : AND2_X1 port map( A1 => n9225, A2 => DATA2_I_3_port, ZN => n11735);
   U116 : AOI21_X1 port map( B1 => n11732, B2 => n11406, A => n11735, ZN => 
                           n11407);
   U117 : OAI21_X1 port map( B1 => n11407, B2 => n1429, A => n11736, ZN => 
                           n11408);
   U118 : AND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n11737)
                           ;
   U119 : AOI21_X1 port map( B1 => n11772, B2 => n11408, A => n11737, ZN => 
                           n11409);
   U120 : OAI21_X1 port map( B1 => n11409, B2 => n1353, A => n11738, ZN => 
                           n11410);
   U121 : AOI22_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, B1 => n11743
                           , B2 => n11410, ZN => n11661);
   U122 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n12448);
   U123 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => 
                           n12448, ZN => n12468);
   U124 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n12469);
   U125 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => 
                           n12469, ZN => n12485);
   U126 : NOR2_X1 port map( A1 => n12468, A2 => n12485, ZN => n12431);
   U127 : NOR2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n11660)
                           ;
   U128 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => DATA1(8), A => n11660,
                           ZN => n11717);
   U129 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n12514
                           );
   U130 : OAI21_X1 port map( B1 => DATA1(9), B2 => DATA2_I_9_port, A => n12514,
                           ZN => n11664);
   U131 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n12427);
   U132 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n12427, ZN => n12515);
   U133 : NAND2_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, ZN => 
                           n12432);
   U134 : OAI21_X1 port map( B1 => DATA1(14), B2 => DATA2_I_14_port, A => 
                           n12432, ZN => n12451);
   U135 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n12429);
   U136 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => 
                           n12429, ZN => n12504);
   U137 : NOR4_X1 port map( A1 => n11664, A2 => n12515, A3 => n12451, A4 => 
                           n12504, ZN => n11411);
   U138 : NAND3_X1 port map( A1 => n12431, A2 => n11717, A3 => n11411, ZN => 
                           n11414);
   U139 : INV_X1 port map( A => n12451, ZN => n12459);
   U140 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n11413);
   U141 : INV_X1 port map( A => DATA1(8), ZN => n12656);
   U142 : INV_X1 port map( A => DATA2_I_8_port, ZN => n11412);
   U143 : NOR3_X1 port map( A1 => n12656, A2 => n11664, A3 => n11412, ZN => 
                           n11662);
   U144 : INV_X1 port map( A => n11662, ZN => n12522);
   U145 : AOI21_X1 port map( B1 => n12514, B2 => n12522, A => n12515, ZN => 
                           n12511);
   U146 : AOI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n12511, ZN => n12505);
   U147 : OAI21_X1 port map( B1 => n11413, B2 => n12505, A => n12429, ZN => 
                           n12484);
   U148 : NOR2_X1 port map( A1 => n12469, A2 => n12468, ZN => n12430);
   U149 : AOI21_X1 port map( B1 => n12431, B2 => n12484, A => n12430, ZN => 
                           n12450);
   U150 : NAND2_X1 port map( A1 => n12450, A2 => n12448, ZN => n12454);
   U151 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n12459, B2 => n12454, ZN => n12439);
   U152 : OAI21_X1 port map( B1 => n11661, B2 => n11414, A => n12439, ZN => 
                           n11415);
   U153 : AOI22_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, B1 => 
                           n12442, B2 => n11415, ZN => n11427);
   U154 : NOR2_X1 port map( A1 => n13225, A2 => n11427, ZN => n12388);
   U155 : AND2_X1 port map( A1 => n1807, A2 => n12388, ZN => n7047);
   U156 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n11420);
   U157 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => 
                           n11420, ZN => n1806);
   U158 : INV_X1 port map( A => n12388, ZN => n12403);
   U159 : INV_X1 port map( A => n1806, ZN => n11423);
   U160 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n11421);
   U161 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n11418);
   U162 : INV_X1 port map( A => n11418, ZN => n11419);
   U163 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n11416);
   U164 : INV_X1 port map( A => n11416, ZN => n11417);
   U165 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n12405);
   U166 : OAI21_X1 port map( B1 => DATA1(17), B2 => DATA2_I_17_port, A => 
                           n11416, ZN => n12408);
   U167 : NOR2_X1 port map( A1 => n12405, A2 => n12408, ZN => n12404);
   U168 : NOR2_X1 port map( A1 => n11417, A2 => n12404, ZN => n12385);
   U169 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => 
                           n11418, ZN => n12386);
   U170 : NOR2_X1 port map( A1 => n12385, A2 => n12386, ZN => n12384);
   U171 : NOR2_X1 port map( A1 => n11419, A2 => n12384, ZN => n12367);
   U172 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n11425);
   U173 : OAI21_X1 port map( B1 => n11421, B2 => n12367, A => n11425, ZN => 
                           n12316);
   U174 : INV_X1 port map( A => n11420, ZN => n11422);
   U175 : AOI21_X1 port map( B1 => n11423, B2 => n12316, A => n11422, ZN => 
                           n12307);
   U176 : NAND2_X1 port map( A1 => n12756, A2 => n11427, ZN => n12406);
   U177 : NOR2_X1 port map( A1 => n12409, A2 => n12408, ZN => n12407);
   U178 : AOI21_X1 port map( B1 => DATA2_I_17_port, B2 => DATA1(17), A => 
                           n12407, ZN => n12383);
   U179 : NOR2_X1 port map( A1 => n12383, A2 => n12386, ZN => n12382);
   U180 : AOI21_X1 port map( B1 => DATA2_I_18_port, B2 => DATA1(18), A => 
                           n12382, ZN => n12366);
   U181 : OAI21_X1 port map( B1 => n12366, B2 => n11421, A => n11425, ZN => 
                           n12317);
   U182 : AOI21_X1 port map( B1 => n11423, B2 => n12317, A => n11422, ZN => 
                           n12308);
   U183 : OAI22_X1 port map( A1 => n12403, A2 => n12307, B1 => n12406, B2 => 
                           n12308, ZN => n11424);
   U184 : INV_X1 port map( A => n11424, ZN => n3860);
   U185 : INV_X1 port map( A => n12406, ZN => n1808);
   U186 : INV_X1 port map( A => DATA1(2), ZN => n1860);
   U187 : NAND2_X1 port map( A1 => DATA1(29), A2 => n4395, ZN => n11944);
   U188 : INV_X1 port map( A => n11944, ZN => n1799);
   U189 : INV_X1 port map( A => DATA2(31), ZN => n12757);
   U190 : NOR2_X1 port map( A1 => n12757, A2 => DATA1(31), ZN => n12632);
   U191 : INV_X1 port map( A => n12632, ZN => n7325);
   U192 : NAND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n12275);
   U193 : OAI21_X1 port map( B1 => DATA1(21), B2 => DATA2_I_21_port, A => 
                           n12275, ZN => n1805);
   U194 : NAND2_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, ZN => 
                           n11429);
   U195 : OAI21_X1 port map( B1 => DATA1(23), B2 => DATA2_I_23_port, A => 
                           n11429, ZN => n12283);
   U196 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n12282);
   U197 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => 
                           n11425, ZN => n12369);
   U198 : OR4_X1 port map( A1 => n12386, A2 => n12408, A3 => n1807, A4 => 
                           n12369, ZN => n11426);
   U199 : NOR4_X1 port map( A1 => n11427, A2 => n1806, A3 => n1805, A4 => 
                           n11426, ZN => n11428);
   U200 : OAI21_X1 port map( B1 => n12308, B2 => n1805, A => n12275, ZN => 
                           n12279);
   U201 : XOR2_X1 port map( A => DATA2_I_22_port, B => DATA1(22), Z => n12281);
   U202 : OAI21_X1 port map( B1 => n11428, B2 => n12279, A => n12281, ZN => 
                           n11430);
   U203 : OAI221_X1 port map( B1 => n12283, B2 => n12282, C1 => n12283, C2 => 
                           n11430, A => n11429, ZN => n11431);
   U204 : NOR2_X1 port map( A1 => n13225, A2 => n11431, ZN => n1803);
   U205 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n11943);
   U206 : INV_X1 port map( A => n11943, ZN => n4421);
   U207 : NAND2_X1 port map( A1 => n12756, A2 => n11431, ZN => n1804);
   U208 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n1802);
   U209 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n11432);
   U210 : INV_X1 port map( A => n11432, ZN => n11647);
   U211 : OAI21_X1 port map( B1 => DATA1(25), B2 => DATA2_I_25_port, A => 
                           n11432, ZN => n12259);
   U212 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n12265);
   U213 : NOR2_X1 port map( A1 => n12259, A2 => n12265, ZN => n12258);
   U214 : OR2_X1 port map( A1 => n11647, A2 => n12258, ZN => n11645);
   U215 : OAI21_X1 port map( B1 => DATA1(26), B2 => DATA2_I_26_port, A => n1802
                           , ZN => n12248);
   U216 : INV_X1 port map( A => n12248, ZN => n11646);
   U217 : NAND2_X1 port map( A1 => n11645, A2 => n11646, ZN => n11945);
   U218 : INV_X1 port map( A => n11945, ZN => n1801);
   U219 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n6740);
   U220 : OAI21_X1 port map( B1 => DATA1(30), B2 => DATA2_I_30_port, A => n6740
                           , ZN => n11946);
   U221 : INV_X1 port map( A => n11946, ZN => n1828);
   U222 : INV_X1 port map( A => DATA1(3), ZN => n1859);
   U223 : INV_X1 port map( A => DATA1(31), ZN => n1837);
   U224 : NOR2_X1 port map( A1 => n1837, A2 => DATA2(31), ZN => n12585);
   U225 : INV_X1 port map( A => n12585, ZN => n1836);
   U226 : OAI22_X1 port map( A1 => n9109, A2 => n8958, B1 => n8893, B2 => n8643
                           , ZN => n11526);
   U227 : AOI211_X1 port map( C1 => n8543, C2 => n8853, A => n8661, B => n8660,
                           ZN => n11446);
   U228 : OAI211_X1 port map( C1 => n8889, C2 => n8541, A => n8653, B => n8652,
                           ZN => n11455);
   U229 : OAI211_X1 port map( C1 => n8860, C2 => n8889, A => n8659, B => n8658,
                           ZN => n11473);
   U230 : AOI22_X1 port map( A1 => n8906, A2 => n11455, B1 => n8809, B2 => 
                           n11473, ZN => n11434);
   U231 : OAI211_X1 port map( C1 => n9012, C2 => n8857, A => n8663, B => n8662,
                           ZN => n11457);
   U232 : OAI211_X1 port map( C1 => n8856, C2 => n9094, A => n8657, B => n8656,
                           ZN => n11456);
   U233 : AOI22_X1 port map( A1 => n9105, A2 => n11457, B1 => n11456, B2 => 
                           n13170, ZN => n11433);
   U234 : OAI211_X1 port map( C1 => n11446, C2 => n13190, A => n11434, B => 
                           n11433, ZN => n11476);
   U235 : AOI211_X1 port map( C1 => n9202, C2 => n9187, A => n8667, B => n8666,
                           ZN => n11449);
   U236 : INV_X1 port map( A => n11446, ZN => n11454);
   U237 : AOI22_X1 port map( A1 => n8906, A2 => n11473, B1 => n11454, B2 => 
                           n13192, ZN => n11436);
   U238 : AOI22_X1 port map( A1 => n11456, A2 => n13144, B1 => n11457, B2 => 
                           n13153, ZN => n11435);
   U239 : OAI211_X1 port map( C1 => n9019, C2 => n11449, A => n11436, B => 
                           n11435, ZN => n11465);
   U240 : AOI211_X1 port map( C1 => n8546, C2 => n8853, A => n8665, B => n8664,
                           ZN => n11450);
   U241 : INV_X1 port map( A => n11456, ZN => n11470);
   U242 : OAI22_X1 port map( A1 => n8895, A2 => n11450, B1 => n11470, B2 => 
                           n13164, ZN => n11438);
   U243 : OAI22_X1 port map( A1 => n9022, A2 => n11446, B1 => n11449, B2 => 
                           n8972, ZN => n11437);
   U244 : AOI211_X1 port map( C1 => n11457, C2 => n13144, A => n11438, B => 
                           n11437, ZN => n11463);
   U245 : INV_X1 port map( A => n11463, ZN => n11439);
   U246 : AOI222_X1 port map( A1 => n9011, A2 => n11476, B1 => n8907, B2 => 
                           n11465, C1 => n9008, C2 => n11439, ZN => n11503);
   U247 : INV_X1 port map( A => n11503, ZN => n11494);
   U248 : AOI22_X1 port map( A1 => n8546, A2 => n9016, B1 => n8545, B2 => n8852
                           , ZN => n11440);
   U249 : OAI211_X1 port map( C1 => n9094, C2 => n13160, A => n8670, B => 
                           n11440, ZN => n11510);
   U250 : OAI22_X1 port map( A1 => n9104, A2 => n11450, B1 => n9182, B2 => 
                           n11449, ZN => n11444);
   U251 : AOI22_X1 port map( A1 => n8853, A2 => n8545, B1 => n8543, B2 => n9186
                           , ZN => n11441);
   U252 : OAI211_X1 port map( C1 => n8857, C2 => n8889, A => n8669, B => n11441
                           , ZN => n11513);
   U253 : INV_X1 port map( A => n11513, ZN => n11451);
   U254 : OAI22_X1 port map( A1 => n9094, A2 => n13191, B1 => n9180, B2 => 
                           n13160, ZN => n11442);
   U255 : AOI211_X1 port map( C1 => n8545, C2 => n9185, A => n9203, B => n11442
                           , ZN => n12395);
   U256 : OAI22_X1 port map( A1 => n9022, A2 => n11451, B1 => n8895, B2 => 
                           n12395, ZN => n11443);
   U257 : AOI211_X1 port map( C1 => n9216, C2 => n11510, A => n11444, B => 
                           n11443, ZN => n11495);
   U258 : INV_X1 port map( A => n11450, ZN => n11496);
   U259 : AOI22_X1 port map( A1 => n11457, A2 => n13141, B1 => n11496, B2 => 
                           n13146, ZN => n11445);
   U260 : INV_X1 port map( A => n11445, ZN => n11448);
   U261 : OAI22_X1 port map( A1 => n11446, A2 => n9104, B1 => n9165, B2 => 
                           n11449, ZN => n11447);
   U262 : AOI211_X1 port map( C1 => n9215, C2 => n11513, A => n11448, B => 
                           n11447, ZN => n11462);
   U263 : OAI22_X1 port map( A1 => n13139, A2 => n11450, B1 => n9181, B2 => 
                           n11449, ZN => n11453);
   U264 : INV_X1 port map( A => n11510, ZN => n12396);
   U265 : OAI22_X1 port map( A1 => n13145, A2 => n11451, B1 => n13140, B2 => 
                           n12396, ZN => n11452);
   U266 : AOI211_X1 port map( C1 => n11454, C2 => n8906, A => n11453, B => 
                           n11452, ZN => n11460);
   U267 : OAI222_X1 port map( A1 => n8975, A2 => n11495, B1 => n11462, B2 => 
                           n8896, C1 => n9103, C2 => n11460, ZN => n11520);
   U268 : INV_X1 port map( A => n11520, ZN => n12490);
   U269 : INV_X1 port map( A => n11455, ZN => n11482);
   U270 : OAI211_X1 port map( C1 => n8889, C2 => n8542, A => n8655, B => n8654,
                           ZN => n11788);
   U271 : AOI22_X1 port map( A1 => n9216, A2 => n11456, B1 => n11788, B2 => 
                           n13141, ZN => n11459);
   U272 : AOI22_X1 port map( A1 => n8806, A2 => n11473, B1 => n9215, B2 => 
                           n11457, ZN => n11458);
   U273 : OAI211_X1 port map( C1 => n11482, C2 => n13142, A => n11459, B => 
                           n11458, ZN => n11475);
   U274 : AOI222_X1 port map( A1 => n11465, A2 => n9008, B1 => n11476, B2 => 
                           n8907, C1 => n11475, C2 => n9011, ZN => n11786);
   U275 : OAI22_X1 port map( A1 => n13196, A2 => n12490, B1 => n11786, B2 => 
                           n8897, ZN => n11467);
   U276 : INV_X1 port map( A => n11460, ZN => n11502);
   U277 : OAI22_X1 port map( A1 => n11463, A2 => n8896, B1 => n11462, B2 => 
                           n9103, ZN => n11461);
   U278 : AOI21_X1 port map( B1 => n13183, B2 => n11502, A => n11461, ZN => 
                           n12491);
   U279 : OAI22_X1 port map( A1 => n11463, A2 => n9103, B1 => n8975, B2 => 
                           n11462, ZN => n11464);
   U280 : AOI21_X1 port map( B1 => n11465, B2 => n13159, A => n11464, ZN => 
                           n11509);
   U281 : OAI22_X1 port map( A1 => n9107, A2 => n12491, B1 => n11509, B2 => 
                           n8561, ZN => n11466);
   U282 : AOI211_X1 port map( C1 => n11494, C2 => n13167, A => n11467, B => 
                           n11466, ZN => n11796);
   U283 : INV_X1 port map( A => n11796, ZN => n11508);
   U284 : INV_X1 port map( A => n11509, ZN => n11481);
   U285 : OAI22_X1 port map( A1 => n9104, A2 => n8647, B1 => n8644, B2 => 
                           n13164, ZN => n11469);
   U286 : INV_X1 port map( A => n11788, ZN => n11483);
   U287 : OAI22_X1 port map( A1 => n11483, A2 => n13139, B1 => n11482, B2 => 
                           n13145, ZN => n11468);
   U288 : AOI211_X1 port map( C1 => n9017, C2 => n11473, A => n11469, B => 
                           n11468, ZN => n11487);
   U289 : OAI22_X1 port map( A1 => n11470, A2 => n13140, B1 => n8647, B2 => 
                           n13164, ZN => n11472);
   U290 : OAI22_X1 port map( A1 => n11483, A2 => n9104, B1 => n11482, B2 => 
                           n13139, ZN => n11471);
   U291 : AOI211_X1 port map( C1 => n9216, C2 => n11473, A => n11472, B => 
                           n11471, ZN => n11478);
   U292 : INV_X1 port map( A => n11478, ZN => n11488);
   U293 : AOI22_X1 port map( A1 => n9008, A2 => n11475, B1 => n8907, B2 => 
                           n11488, ZN => n11474);
   U294 : OAI21_X1 port map( B1 => n11487, B2 => n13185, A => n11474, ZN => 
                           n11853);
   U295 : INV_X1 port map( A => n11853, ZN => n11813);
   U296 : OAI22_X1 port map( A1 => n11786, A2 => n13180, B1 => n11813, B2 => 
                           n13143, ZN => n11480);
   U297 : AOI22_X1 port map( A1 => n9008, A2 => n11476, B1 => n8907, B2 => 
                           n11475, ZN => n11477);
   U298 : OAI21_X1 port map( B1 => n11478, B2 => n13185, A => n11477, ZN => 
                           n11489);
   U299 : INV_X1 port map( A => n11489, ZN => n11814);
   U300 : OAI22_X1 port map( A1 => n11503, A2 => n9107, B1 => n11814, B2 => 
                           n13148, ZN => n11479);
   U301 : AOI211_X1 port map( C1 => n9102, C2 => n11481, A => n11480, B => 
                           n11479, ZN => n11817);
   U302 : OAI22_X1 port map( A1 => n8647, A2 => n9165, B1 => n8644, B2 => 
                           n13142, ZN => n11485);
   U303 : OAI22_X1 port map( A1 => n11483, A2 => n13145, B1 => n11482, B2 => 
                           n13140, ZN => n11484);
   U304 : AOI211_X1 port map( C1 => n8906, C2 => n9201, A => n11485, B => 
                           n11484, ZN => n11486);
   U305 : INV_X1 port map( A => n11486, ZN => n11812);
   U306 : INV_X1 port map( A => n11487, ZN => n11791);
   U307 : AOI222_X1 port map( A1 => n9011, A2 => n11812, B1 => n8907, B2 => 
                           n11791, C1 => n9008, C2 => n11488, ZN => n11792);
   U308 : INV_X1 port map( A => n11792, ZN => n12191);
   U309 : AOI22_X1 port map( A1 => n9183, A2 => n12191, B1 => n11853, B2 => 
                           n13167, ZN => n11491);
   U310 : AOI22_X1 port map( A1 => n9162, A2 => n11489, B1 => n9102, B2 => 
                           n11494, ZN => n11490);
   U311 : OAI211_X1 port map( C1 => n11786, C2 => n13150, A => n11491, B => 
                           n11490, ZN => n11856);
   U312 : INV_X1 port map( A => n11856, ZN => n12197);
   U313 : OAI22_X1 port map( A1 => n11817, A2 => n13181, B1 => n12197, B2 => 
                           n8801, ZN => n11507);
   U314 : OAI22_X1 port map( A1 => n11814, A2 => n8897, B1 => n9217, B2 => 
                           n12491, ZN => n11493);
   U315 : OAI22_X1 port map( A1 => n11786, A2 => n9106, B1 => n9107, B2 => 
                           n11509, ZN => n11492);
   U316 : AOI211_X1 port map( C1 => n9162, C2 => n11494, A => n11493, B => 
                           n11492, ZN => n11818);
   U317 : INV_X1 port map( A => n11495, ZN => n11517);
   U318 : AOI22_X1 port map( A1 => n8809, A2 => n11513, B1 => n8906, B2 => 
                           n11496, ZN => n11501);
   U319 : OAI222_X1 port map( A1 => n8671, A2 => n8966, B1 => n9204, B2 => 
                           n8968, C1 => n9184, C2 => n8672, ZN => n11497);
   U320 : INV_X1 port map( A => n11497, ZN => n12300);
   U321 : AOI22_X1 port map( A1 => n9016, A2 => n11337, B1 => n8544, B2 => 
                           n8851, ZN => n11499);
   U322 : AOI22_X1 port map( A1 => n8546, A2 => n9014, B1 => n9186, B2 => n8545
                           , ZN => n11498);
   U323 : OAI211_X1 port map( C1 => n9028, C2 => n12300, A => n11499, B => 
                           n11498, ZN => n12393);
   U324 : AOI22_X1 port map( A1 => n8806, A2 => n11510, B1 => n13151, B2 => 
                           n12393, ZN => n11500);
   U325 : OAI211_X1 port map( C1 => n12395, C2 => n13179, A => n11501, B => 
                           n11500, ZN => n12416);
   U326 : AOI222_X1 port map( A1 => n11517, A2 => n8907, B1 => n11502, B2 => 
                           n9218, C1 => n12416, C2 => n9098, ZN => n12489);
   U327 : OAI22_X1 port map( A1 => n11503, A2 => n8897, B1 => n9217, B2 => 
                           n12489, ZN => n11505);
   U328 : OAI22_X1 port map( A1 => n11509, A2 => n9031, B1 => n12491, B2 => 
                           n8561, ZN => n11504);
   U329 : AOI211_X1 port map( C1 => n8807, C2 => n11520, A => n11505, B => 
                           n11504, ZN => n12524);
   U330 : OAI22_X1 port map( A1 => n8677, A2 => n11818, B1 => n9027, B2 => 
                           n12524, ZN => n11506);
   U331 : AOI211_X1 port map( C1 => n13172, C2 => n11508, A => n11507, B => 
                           n11506, ZN => n11823);
   U332 : INV_X1 port map( A => n11817, ZN => n11857);
   U333 : OAI22_X1 port map( A1 => n11509, A2 => n13143, B1 => n12491, B2 => 
                           n13148, ZN => n11519);
   U334 : INV_X1 port map( A => n12393, ZN => n11516);
   U335 : INV_X1 port map( A => n12395, ZN => n12373);
   U336 : AOI22_X1 port map( A1 => n8809, A2 => n11510, B1 => n8806, B2 => 
                           n12373, ZN => n11515);
   U337 : AOI22_X1 port map( A1 => n8545, A2 => n9014, B1 => n9016, B2 => n8544
                           , ZN => n11512);
   U338 : OAI222_X1 port map( A1 => n8671, A2 => n8968, B1 => n8966, B2 => 
                           n8672, C1 => n9184, C2 => n8668, ZN => n12302);
   U339 : AOI22_X1 port map( A1 => n9186, A2 => n11337, B1 => n8854, B2 => 
                           n12302, ZN => n11511);
   U340 : OAI211_X1 port map( C1 => n9180, C2 => n12300, A => n11512, B => 
                           n11511, ZN => n12392);
   U341 : AOI22_X1 port map( A1 => n8906, A2 => n11513, B1 => n9215, B2 => 
                           n12392, ZN => n11514);
   U342 : OAI211_X1 port map( C1 => n9020, C2 => n11516, A => n11515, B => 
                           n11514, ZN => n12417);
   U343 : AOI222_X1 port map( A1 => n12416, A2 => n8907, B1 => n12417, B2 => 
                           n9098, C1 => n11517, C2 => n9218, ZN => n12488);
   U344 : OAI22_X1 port map( A1 => n9217, A2 => n12488, B1 => n12489, B2 => 
                           n13150, ZN => n11518);
   U345 : AOI211_X1 port map( C1 => n9162, C2 => n11520, A => n11519, B => 
                           n11518, ZN => n12523);
   U346 : OAI22_X1 port map( A1 => n8677, A2 => n11796, B1 => n12523, B2 => 
                           n13165, ZN => n11522);
   U347 : OAI22_X1 port map( A1 => n11818, A2 => n9166, B1 => n9167, B2 => 
                           n12524, ZN => n11521);
   U348 : AOI211_X1 port map( C1 => n11857, C2 => n13166, A => n11522, B => 
                           n11521, ZN => n11800);
   U349 : OAI22_X1 port map( A1 => n11823, A2 => n9163, B1 => n8908, B2 => 
                           n11800, ZN => n11523);
   U350 : AOI21_X1 port map( B1 => n13204, B2 => n11523, A => n8642, ZN => 
                           n11524);
   U351 : NAND2_X1 port map( A1 => n8957, A2 => n11524, ZN => n11525);
   U352 : AOI211_X1 port map( C1 => n9210, C2 => n8880, A => n11526, B => 
                           n11525, ZN => n11527);
   U353 : INV_X1 port map( A => n11527, ZN => OUTALU(6));
   U354 : NOR2_X1 port map( A1 => n9220, A2 => n13225, ZN => n7166);
   U355 : NOR2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n13092);
   U356 : INV_X1 port map( A => n13123, ZN => n11315);
   U357 : OAI21_X1 port map( B1 => n13088, B2 => n13077, A => n11553, ZN => 
                           n11528);
   U358 : INV_X1 port map( A => n11528, ZN => n13220);
   U359 : NOR2_X1 port map( A1 => n13082, A2 => DATA2(1), ZN => n13081);
   U360 : NAND2_X1 port map( A1 => n11895, A2 => n13081, ZN => n12163);
   U361 : INV_X1 port map( A => DATA1(24), ZN => n12700);
   U362 : NAND2_X1 port map( A1 => n11895, A2 => n13091, ZN => n12232);
   U363 : INV_X1 port map( A => n12232, ZN => n12215);
   U364 : INV_X1 port map( A => DATA1(25), ZN => n12256);
   U365 : NAND2_X1 port map( A1 => n13092, A2 => n11895, ZN => n12341);
   U366 : NOR2_X1 port map( A1 => n12256, A2 => n12341, ZN => n11676);
   U367 : INV_X1 port map( A => DATA1(21), ZN => n12692);
   U368 : NOR2_X1 port map( A1 => n11895, A2 => n12692, ZN => n11563);
   U369 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(22), A => n11676, B => 
                           n11563, ZN => n11529);
   U370 : NAND3_X1 port map( A1 => n13082, A2 => DATA2(1), A3 => n11895, ZN => 
                           n12545);
   U371 : NAND2_X1 port map( A1 => DATA1(23), A2 => n12216, ZN => n11578);
   U372 : OAI211_X1 port map( C1 => n12163, C2 => n12700, A => n11529, B => 
                           n11578, ZN => n1843);
   U373 : NAND3_X1 port map( A1 => n13088, A2 => n11553, A3 => n11532, ZN => 
                           n11906);
   U374 : INV_X1 port map( A => DATA1(22), ZN => n12554);
   U375 : NOR2_X1 port map( A1 => n12554, A2 => n12545, ZN => n11575);
   U376 : INV_X1 port map( A => DATA1(20), ZN => n12319);
   U377 : NOR2_X1 port map( A1 => n11895, A2 => n12319, ZN => n11558);
   U378 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(21), A => n11575, B => 
                           n11558, ZN => n11530);
   U379 : NAND2_X1 port map( A1 => DATA1(23), A2 => n12332, ZN => n11581);
   U380 : OAI211_X1 port map( C1 => n12341, C2 => n12700, A => n11530, B => 
                           n11581, ZN => n11887);
   U381 : INV_X1 port map( A => DATA1(26), ZN => n12572);
   U382 : NOR2_X1 port map( A1 => n12572, A2 => n12341, ZN => n11667);
   U383 : NOR2_X1 port map( A1 => n11895, A2 => n12554, ZN => n11568);
   U384 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(23), A => n11667, B => 
                           n11568, ZN => n11531);
   U385 : NAND2_X1 port map( A1 => DATA1(25), A2 => n12332, ZN => n11672);
   U386 : OAI211_X1 port map( C1 => n12545, C2 => n12700, A => n11531, B => 
                           n11672, ZN => n11894);
   U387 : INV_X1 port map( A => n12237, ZN => n12182);
   U388 : AOI222_X1 port map( A1 => n11887, A2 => n11781, B1 => n11894, B2 => 
                           n12182, C1 => n1843, C2 => n1865, ZN => n1842);
   U389 : INV_X1 port map( A => n13121, ZN => n1869);
   U390 : INV_X1 port map( A => DATA1(23), ZN => n1846);
   U391 : NOR2_X1 port map( A1 => n1846, A2 => n12341, ZN => n11670);
   U392 : NOR2_X1 port map( A1 => n12692, A2 => n12545, ZN => n11583);
   U393 : AOI211_X1 port map( C1 => DATA1(19), C2 => n11917, A => n11670, B => 
                           n11583, ZN => n11534);
   U394 : NOR2_X1 port map( A1 => n12319, A2 => n12232, ZN => n11564);
   U395 : INV_X1 port map( A => n11564, ZN => n11533);
   U396 : OAI211_X1 port map( C1 => n12163, C2 => n12554, A => n11534, B => 
                           n11533, ZN => n11886);
   U397 : CLKBUF_X1 port map( A => n1865, Z => n11844);
   U398 : AOI222_X1 port map( A1 => n11886, A2 => n11528, B1 => n1843, B2 => 
                           n12182, C1 => n11887, C2 => n11844, ZN => n13134);
   U399 : OAI22_X1 port map( A1 => n11315, A2 => n1842, B1 => n1869, B2 => 
                           n13134, ZN => n11535);
   U400 : INV_X1 port map( A => n11535, ZN => n6541);
   U401 : INV_X1 port map( A => FUNC(0), ZN => n1832);
   U402 : NAND3_X1 port map( A1 => FUNC(1), A2 => n1832, A3 => n11536, ZN => 
                           n1835);
   U403 : INV_X1 port map( A => FUNC(3), ZN => n12755);
   U404 : NAND3_X1 port map( A1 => FUNC(2), A2 => n11650, A3 => n12755, ZN => 
                           n7822);
   U405 : INV_X1 port map( A => DATA2(7), ZN => n12783);
   U406 : INV_X1 port map( A => DATA2(6), ZN => n12784);
   U407 : INV_X1 port map( A => DATA2(11), ZN => n12777);
   U408 : INV_X1 port map( A => DATA2(13), ZN => n12775);
   U409 : NAND4_X1 port map( A1 => n12783, A2 => n12784, A3 => n12777, A4 => 
                           n12775, ZN => n11538);
   U410 : INV_X1 port map( A => DATA2(14), ZN => n12774);
   U411 : INV_X1 port map( A => DATA2(12), ZN => n12776);
   U412 : INV_X1 port map( A => DATA2(10), ZN => n12778);
   U413 : INV_X1 port map( A => DATA2(15), ZN => n12773);
   U414 : NAND4_X1 port map( A1 => n12774, A2 => n12776, A3 => n12778, A4 => 
                           n12773, ZN => n11537);
   U415 : NOR4_X1 port map( A1 => DATA2(8), A2 => DATA2(9), A3 => n11538, A4 =>
                           n11537, ZN => n11544);
   U416 : OR4_X1 port map( A1 => DATA1(7), A2 => n9223, A3 => DATA1(11), A4 => 
                           DATA1(13), ZN => n11542);
   U417 : INV_X1 port map( A => DATA1(14), ZN => n12675);
   U418 : INV_X1 port map( A => DATA1(12), ZN => n12668);
   U419 : INV_X1 port map( A => DATA1(10), ZN => n12571);
   U420 : INV_X1 port map( A => DATA1(15), ZN => n12424);
   U421 : NAND4_X1 port map( A1 => n12675, A2 => n12668, A3 => n12571, A4 => 
                           n12424, ZN => n11541);
   U422 : INV_X1 port map( A => DATA1(4), ZN => n11803);
   U423 : NAND4_X1 port map( A1 => n11764, A2 => n13173, A3 => n13149, A4 => 
                           n11803, ZN => n11540);
   U424 : INV_X1 port map( A => DATA1(6), ZN => n12651);
   U425 : INV_X1 port map( A => DATA1(9), ZN => n11659);
   U426 : NAND4_X1 port map( A1 => n11332, A2 => n12656, A3 => n12651, A4 => 
                           n11659, ZN => n11539);
   U427 : NOR4_X1 port map( A1 => n11542, A2 => n11541, A3 => n11540, A4 => 
                           n11539, ZN => n11543);
   U428 : CLKBUF_X1 port map( A => n6095, Z => n13224);
   U429 : NAND2_X1 port map( A1 => n12783, A2 => DATA1(7), ZN => n12567);
   U430 : INV_X1 port map( A => n12567, ZN => n12653);
   U431 : INV_X1 port map( A => n1835, ZN => n12535);
   U432 : AOI22_X1 port map( A1 => n12653, A2 => n12535, B1 => n13224, B2 => 
                           n8765, ZN => n11545);
   U433 : INV_X1 port map( A => n11545, ZN => n1829);
   U434 : INV_X1 port map( A => n12237, ZN => n13223);
   U435 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(4), ZN => n13089);
   U436 : NOR2_X1 port map( A1 => n13077, A2 => n13089, ZN => n13086);
   U437 : NAND2_X1 port map( A1 => n13091, A2 => n13086, ZN => n11870);
   U438 : INV_X1 port map( A => n11870, ZN => n11546);
   U439 : INV_X1 port map( A => DATA2(5), ZN => n12785);
   U440 : NAND4_X1 port map( A1 => FUNC(1), A2 => FUNC(2), A3 => n12785, A4 => 
                           n1832, ZN => n11869);
   U441 : NOR2_X1 port map( A1 => n11546, A2 => n11869, ZN => n11547);
   U442 : NAND2_X1 port map( A1 => n11547, A2 => n12755, ZN => n1834);
   U443 : NAND2_X1 port map( A1 => FUNC(3), A2 => n11547, ZN => n1833);
   U444 : INV_X1 port map( A => n11661, ZN => n12465);
   U445 : NAND2_X1 port map( A1 => n12465, A2 => n12756, ZN => n12434);
   U446 : INV_X1 port map( A => n12434, ZN => n7147);
   U447 : NOR2_X1 port map( A1 => n9205, A2 => n12545, ZN => n11548);
   U448 : NOR2_X1 port map( A1 => n13149, A2 => n12163, ZN => n12177);
   U449 : AOI211_X1 port map( C1 => n12215, C2 => n9222, A => n11548, B => 
                           n12177, ZN => n11549);
   U450 : NAND2_X1 port map( A1 => DATA1(4), A2 => n12541, ZN => n11838);
   U451 : OAI211_X1 port map( C1 => n11895, C2 => n13173, A => n11549, B => 
                           n11838, ZN => n11802);
   U452 : NOR2_X1 port map( A1 => n11764, A2 => n12163, ZN => n11841);
   U453 : NOR2_X1 port map( A1 => n12651, A2 => n12341, ZN => n11777);
   U454 : AOI211_X1 port map( C1 => n13177, C2 => n11917, A => n11841, B => 
                           n11777, ZN => n11551);
   U455 : NOR2_X1 port map( A1 => n13149, A2 => n12232, ZN => n12539);
   U456 : INV_X1 port map( A => n12539, ZN => n11550);
   U457 : OAI211_X1 port map( C1 => n12545, C2 => n11803, A => n11551, B => 
                           n11550, ZN => n11711);
   U458 : NOR2_X1 port map( A1 => n11803, A2 => n12163, ZN => n11836);
   U459 : NOR2_X1 port map( A1 => n13149, A2 => n12545, ZN => n12337);
   U460 : AOI211_X1 port map( C1 => n12215, C2 => n9223, A => n11836, B => 
                           n12337, ZN => n11552);
   U461 : NAND2_X1 port map( A1 => DATA1(5), A2 => n12541, ZN => n11775);
   U462 : OAI211_X1 port map( C1 => n11332, C2 => n11895, A => n11552, B => 
                           n11775, ZN => n11760);
   U463 : AOI222_X1 port map( A1 => n11802, A2 => n11781, B1 => n11711, B2 => 
                           n13223, C1 => n11760, C2 => n11844, ZN => n1830);
   U464 : OR2_X1 port map( A1 => n13108, A2 => n1830, ZN => n6338);
   U465 : INV_X1 port map( A => n13108, ZN => n13222);
   U466 : INV_X1 port map( A => n13222, ZN => n13138);
   U467 : NAND2_X1 port map( A1 => n11553, A2 => n13138, ZN => n13135);
   U468 : INV_X1 port map( A => n13135, ZN => n13221);
   U469 : AOI22_X1 port map( A1 => DATA1(16), A2 => n12332, B1 => DATA1(17), B2
                           => n12216, ZN => n11557);
   U470 : NAND2_X1 port map( A1 => DATA1(15), A2 => n12541, ZN => n11556);
   U471 : CLKBUF_X1 port map( A => n12215, Z => n12179);
   U472 : NAND2_X1 port map( A1 => DATA1(18), A2 => n12179, ZN => n11555);
   U473 : NAND2_X1 port map( A1 => DATA1(19), A2 => n11917, ZN => n11554);
   U474 : NAND4_X1 port map( A1 => n11557, A2 => n11556, A3 => n11555, A4 => 
                           n11554, ZN => n11566);
   U475 : INV_X1 port map( A => n11566, ZN => n11689);
   U476 : INV_X1 port map( A => DATA1(16), ZN => n12613);
   U477 : INV_X1 port map( A => DATA1(18), ZN => n12687);
   U478 : NOR2_X1 port map( A1 => n12687, A2 => n12545, ZN => n11559);
   U479 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(19), A => n11559, B => 
                           n11558, ZN => n11560);
   U480 : NAND2_X1 port map( A1 => DATA1(17), A2 => n12332, ZN => n11864);
   U481 : OAI211_X1 port map( C1 => n12341, C2 => n12613, A => n11560, B => 
                           n11864, ZN => n11572);
   U482 : AOI22_X1 port map( A1 => DATA1(16), A2 => n12216, B1 => DATA1(17), B2
                           => n12215, ZN => n11561);
   U483 : NAND2_X1 port map( A1 => DATA1(14), A2 => n12541, ZN => n11616);
   U484 : NAND2_X1 port map( A1 => DATA1(15), A2 => n12332, ZN => n11632);
   U485 : NAND2_X1 port map( A1 => DATA1(18), A2 => n11917, ZN => n11596);
   U486 : NAND4_X1 port map( A1 => n11561, A2 => n11616, A3 => n11632, A4 => 
                           n11596, ZN => n11693);
   U487 : AOI22_X1 port map( A1 => n11781, A2 => n11572, B1 => n13223, B2 => 
                           n11693, ZN => n11562);
   U488 : OAI21_X1 port map( B1 => n11689, B2 => n11906, A => n11562, ZN => 
                           n11699);
   U489 : INV_X1 port map( A => DATA1(17), ZN => n12402);
   U490 : NOR2_X1 port map( A1 => n12687, A2 => n12163, ZN => n11604);
   U491 : NOR3_X1 port map( A1 => n11604, A2 => n11564, A3 => n11563, ZN => 
                           n11565);
   U492 : NAND2_X1 port map( A1 => DATA1(19), A2 => n12216, ZN => n11592);
   U493 : OAI211_X1 port map( C1 => n12341, C2 => n12402, A => n11565, B => 
                           n11592, ZN => n11684);
   U494 : AOI222_X1 port map( A1 => n11684, A2 => n11781, B1 => n11566, B2 => 
                           n13223, C1 => n11572, C2 => n11844, ZN => n11682);
   U495 : INV_X1 port map( A => n11682, ZN => n11694);
   U496 : AOI22_X1 port map( A1 => n13222, A2 => n11699, B1 => n11694, B2 => 
                           n13221, ZN => n11567);
   U497 : INV_X1 port map( A => n11567, ZN => n6208);
   U498 : NOR2_X1 port map( A1 => n12319, A2 => n12545, ZN => n11569);
   U499 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(21), A => n11569, B => 
                           n11568, ZN => n11571);
   U500 : NAND2_X1 port map( A1 => DATA1(19), A2 => n12332, ZN => n11570);
   U501 : OAI211_X1 port map( C1 => n12341, C2 => n12687, A => n11571, B => 
                           n11570, ZN => n11683);
   U502 : INV_X1 port map( A => n11683, ZN => n11574);
   U503 : AOI22_X1 port map( A1 => n12182, A2 => n11572, B1 => n1865, B2 => 
                           n11684, ZN => n11573);
   U504 : OAI21_X1 port map( B1 => n11574, B2 => n13220, A => n11573, ZN => 
                           n1849);
   U505 : NOR2_X1 port map( A1 => n12319, A2 => n12341, ZN => n11598);
   U506 : AOI211_X1 port map( C1 => DATA1(24), C2 => n11917, A => n11598, B => 
                           n11575, ZN => n11576);
   U507 : NAND2_X1 port map( A1 => DATA1(21), A2 => n12332, ZN => n11594);
   U508 : OAI211_X1 port map( C1 => n12232, C2 => n1846, A => n11576, B => 
                           n11594, ZN => n11586);
   U509 : INV_X1 port map( A => n11586, ZN => n11587);
   U510 : NOR2_X1 port map( A1 => n12692, A2 => n12341, ZN => n11580);
   U511 : NOR2_X1 port map( A1 => n12256, A2 => n11895, ZN => n11910);
   U512 : INV_X1 port map( A => n11910, ZN => n11577);
   U513 : OAI211_X1 port map( C1 => n12163, C2 => n12554, A => n11578, B => 
                           n11577, ZN => n11579);
   U514 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(24), A => n11580, B => 
                           n11579, ZN => n11671);
   U515 : NOR2_X1 port map( A1 => n12256, A2 => n12232, ZN => n11898);
   U516 : NAND2_X1 port map( A1 => DATA1(22), A2 => n12541, ZN => n11595);
   U517 : OAI211_X1 port map( C1 => n11895, C2 => n12572, A => n11595, B => 
                           n11581, ZN => n11582);
   U518 : AOI211_X1 port map( C1 => n12216, C2 => DATA1(24), A => n11898, B => 
                           n11582, ZN => n11678);
   U519 : OAI222_X1 port map( A1 => n12237, A2 => n11587, B1 => n11906, B2 => 
                           n11671, C1 => n13220, C2 => n11678, ZN => n6198);
   U520 : NOR2_X1 port map( A1 => n12319, A2 => n12163, ZN => n11590);
   U521 : NOR2_X1 port map( A1 => n11590, A2 => n11583, ZN => n11585);
   U522 : NAND2_X1 port map( A1 => DATA1(19), A2 => n12541, ZN => n11602);
   U523 : NAND2_X1 port map( A1 => DATA1(22), A2 => n12179, ZN => n11584);
   U524 : NAND2_X1 port map( A1 => DATA1(23), A2 => n11917, ZN => n11892);
   U525 : NAND4_X1 port map( A1 => n11585, A2 => n11602, A3 => n11584, A4 => 
                           n11892, ZN => n11685);
   U526 : AOI222_X1 port map( A1 => n11586, A2 => n11781, B1 => n11683, B2 => 
                           n13223, C1 => n11685, C2 => n1865, ZN => n1845);
   U527 : INV_X1 port map( A => n11685, ZN => n11588);
   U528 : OAI222_X1 port map( A1 => n12237, A2 => n11588, B1 => n11906, B2 => 
                           n11587, C1 => n13220, C2 => n11671, ZN => n11681);
   U529 : INV_X1 port map( A => n11681, ZN => n13137);
   U530 : OAI22_X1 port map( A1 => n13135, A2 => n13137, B1 => n13138, B2 => 
                           n1845, ZN => n11589);
   U531 : INV_X1 port map( A => n11589, ZN => n6174);
   U532 : NOR2_X1 port map( A1 => n11895, A2 => n12402, ZN => n11591);
   U533 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(18), A => n11591, B => 
                           n11590, ZN => n11593);
   U534 : OAI211_X1 port map( C1 => n12341, C2 => n12692, A => n11593, B => 
                           n11592, ZN => n11605);
   U535 : AOI22_X1 port map( A1 => DATA1(20), A2 => n12216, B1 => DATA1(19), B2
                           => n12215, ZN => n11597);
   U536 : NAND4_X1 port map( A1 => n11597, A2 => n11596, A3 => n11595, A4 => 
                           n11594, ZN => n11885);
   U537 : AOI222_X1 port map( A1 => n11605, A2 => n11781, B1 => n11886, B2 => 
                           n12182, C1 => n11885, C2 => n1865, ZN => n1847);
   U538 : NOR2_X1 port map( A1 => n11895, A2 => n12613, ZN => n11599);
   U539 : AOI211_X1 port map( C1 => n12332, C2 => DATA1(19), A => n11599, B => 
                           n11598, ZN => n11601);
   U540 : NAND2_X1 port map( A1 => DATA1(17), A2 => n12179, ZN => n11600);
   U541 : OAI211_X1 port map( C1 => n12545, C2 => n12687, A => n11601, B => 
                           n11600, ZN => n11863);
   U542 : AOI222_X1 port map( A1 => n11863, A2 => n11781, B1 => n11885, B2 => 
                           n12182, C1 => n11605, C2 => n11844, ZN => n1848);
   U543 : NAND2_X1 port map( A1 => DATA1(15), A2 => n11917, ZN => n11610);
   U544 : OAI211_X1 port map( C1 => n12545, C2 => n12402, A => n11610, B => 
                           n11602, ZN => n11603);
   U545 : AOI211_X1 port map( C1 => n12179, C2 => DATA1(16), A => n11604, B => 
                           n11603, ZN => n11879);
   U546 : AOI22_X1 port map( A1 => n13223, A2 => n11605, B1 => n11844, B2 => 
                           n11863, ZN => n11606);
   U547 : OAI21_X1 port map( B1 => n11879, B2 => n13220, A => n11606, ZN => 
                           n11882);
   U548 : INV_X1 port map( A => n11882, ZN => n11903);
   U549 : OAI22_X1 port map( A1 => n11315, A2 => n1848, B1 => n1869, B2 => 
                           n11903, ZN => n11607);
   U550 : INV_X1 port map( A => n11607, ZN => n3888);
   U551 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12179, ZN => n11631);
   U552 : NAND2_X1 port map( A1 => DATA1(11), A2 => n12332, ZN => n11622);
   U553 : NAND2_X1 port map( A1 => DATA1(10), A2 => n12541, ZN => n11608);
   U554 : AND3_X1 port map( A1 => n11631, A2 => n11622, A3 => n11608, ZN => 
                           n11609);
   U555 : NAND2_X1 port map( A1 => DATA1(12), A2 => n12216, ZN => n11617);
   U556 : OAI211_X1 port map( C1 => n11895, C2 => n12675, A => n11609, B => 
                           n11617, ZN => n11723);
   U557 : AOI22_X1 port map( A1 => DATA1(12), A2 => n12332, B1 => DATA1(11), B2
                           => n12541, ZN => n11611);
   U558 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12216, ZN => n11636);
   U559 : NAND2_X1 port map( A1 => DATA1(14), A2 => n12179, ZN => n11874);
   U560 : NAND4_X1 port map( A1 => n11611, A2 => n11636, A3 => n11874, A4 => 
                           n11610, ZN => n11695);
   U561 : NOR2_X1 port map( A1 => n12668, A2 => n12341, ZN => n11613);
   U562 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12332, ZN => n11618);
   U563 : NAND2_X1 port map( A1 => DATA1(14), A2 => n12216, ZN => n11630);
   U564 : OAI211_X1 port map( C1 => n11895, C2 => n12613, A => n11618, B => 
                           n11630, ZN => n11612);
   U565 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(15), A => n11613, B => 
                           n11612, ZN => n11697);
   U566 : INV_X1 port map( A => n11697, ZN => n11614);
   U567 : AOI222_X1 port map( A1 => n13223, A2 => n11723, B1 => n1865, B2 => 
                           n11695, C1 => n11781, C2 => n11614, ZN => n11751);
   U568 : INV_X1 port map( A => n11751, ZN => n1853);
   U569 : NOR2_X1 port map( A1 => n12668, A2 => n12232, ZN => n11634);
   U570 : INV_X1 port map( A => DATA1(13), ZN => n12470);
   U571 : NOR2_X1 port map( A1 => n11895, A2 => n12470, ZN => n11876);
   U572 : AOI211_X1 port map( C1 => n12541, C2 => DATA1(9), A => n11634, B => 
                           n11876, ZN => n11615);
   U573 : NAND2_X1 port map( A1 => DATA1(11), A2 => n12216, ZN => n11620);
   U574 : NAND2_X1 port map( A1 => DATA1(10), A2 => n12332, ZN => n11625);
   U575 : NAND3_X1 port map( A1 => n11615, A2 => n11620, A3 => n11625, ZN => 
                           n11750);
   U576 : AOI222_X1 port map( A1 => n11695, A2 => n11781, B1 => n11750, B2 => 
                           n12182, C1 => n11723, C2 => n11844, ZN => n6351);
   U577 : NAND3_X1 port map( A1 => DATA2(3), A2 => n13092, A3 => n13074, ZN => 
                           n13133);
   U578 : AOI22_X1 port map( A1 => DATA1(10), A2 => n11917, B1 => DATA1(11), B2
                           => n12179, ZN => n11619);
   U579 : NAND4_X1 port map( A1 => n11619, A2 => n11618, A3 => n11617, A4 => 
                           n11616, ZN => n11638);
   U580 : INV_X1 port map( A => n11638, ZN => n11641);
   U581 : NOR2_X1 port map( A1 => n11895, A2 => n11659, ZN => n11774);
   U582 : NAND2_X1 port map( A1 => DATA1(10), A2 => n12179, ZN => n11748);
   U583 : OAI211_X1 port map( C1 => n12163, C2 => n12668, A => n11748, B => 
                           n11620, ZN => n11621);
   U584 : AOI211_X1 port map( C1 => n12541, C2 => DATA1(13), A => n11774, B => 
                           n11621, ZN => n11640);
   U585 : NOR2_X1 port map( A1 => n12571, A2 => n12545, ZN => n11719);
   U586 : NAND2_X1 port map( A1 => DATA1(9), A2 => n12179, ZN => n11779);
   U587 : OAI211_X1 port map( C1 => n11895, C2 => n12656, A => n11779, B => 
                           n11622, ZN => n11623);
   U588 : AOI211_X1 port map( C1 => n12541, C2 => DATA1(12), A => n11719, B => 
                           n11623, ZN => n11629);
   U589 : OAI222_X1 port map( A1 => n12237, A2 => n11641, B1 => n11906, B2 => 
                           n11640, C1 => n13220, C2 => n11629, ZN => n11921);
   U590 : NOR2_X1 port map( A1 => n12656, A2 => n12545, ZN => n11778);
   U591 : NOR2_X1 port map( A1 => n11895, A2 => n12651, ZN => n12178);
   U592 : AOI211_X1 port map( C1 => n12541, C2 => DATA1(10), A => n11778, B => 
                           n12178, ZN => n11624);
   U593 : NAND2_X1 port map( A1 => DATA1(7), A2 => n12179, ZN => n11839);
   U594 : OAI211_X1 port map( C1 => n12163, C2 => n11659, A => n11624, B => 
                           n11839, ZN => n11931);
   U595 : NOR2_X1 port map( A1 => n11659, A2 => n12545, ZN => n11747);
   U596 : INV_X1 port map( A => DATA1(7), ZN => n12588);
   U597 : NOR2_X1 port map( A1 => n12656, A2 => n12232, ZN => n11773);
   U598 : INV_X1 port map( A => n11773, ZN => n11626);
   U599 : OAI211_X1 port map( C1 => n11895, C2 => n12588, A => n11626, B => 
                           n11625, ZN => n11627);
   U600 : AOI211_X1 port map( C1 => n12541, C2 => DATA1(11), A => n11747, B => 
                           n11627, ZN => n11929);
   U601 : OAI22_X1 port map( A1 => n11629, A2 => n12237, B1 => n11929, B2 => 
                           n11906, ZN => n11628);
   U602 : AOI21_X1 port map( B1 => n11781, B2 => n11931, A => n11628, ZN => 
                           n13112);
   U603 : OAI222_X1 port map( A1 => n12237, A2 => n11640, B1 => n11906, B2 => 
                           n11629, C1 => n13220, C2 => n11929, ZN => n13117);
   U604 : INV_X1 port map( A => n13117, ZN => n13107);
   U605 : OAI22_X1 port map( A1 => n1869, A2 => n13112, B1 => n13107, B2 => 
                           n11315, ZN => n11643);
   U606 : AOI22_X1 port map( A1 => DATA1(16), A2 => n12541, B1 => DATA1(12), B2
                           => n11917, ZN => n11633);
   U607 : NAND4_X1 port map( A1 => n11633, A2 => n11632, A3 => n11631, A4 => 
                           n11630, ZN => n11877);
   U608 : AOI22_X1 port map( A1 => DATA1(11), A2 => n11917, B1 => DATA1(15), B2
                           => n12541, ZN => n11637);
   U609 : INV_X1 port map( A => n11634, ZN => n11635);
   U610 : NAND2_X1 port map( A1 => DATA1(14), A2 => n12332, ZN => n11686);
   U611 : NAND4_X1 port map( A1 => n11637, A2 => n11636, A3 => n11635, A4 => 
                           n11686, ZN => n11639);
   U612 : AOI222_X1 port map( A1 => n11638, A2 => n11781, B1 => n11877, B2 => 
                           n12182, C1 => n11639, C2 => n11844, ZN => n13130);
   U613 : INV_X1 port map( A => n11639, ZN => n11904);
   U614 : OAI222_X1 port map( A1 => n12237, A2 => n11904, B1 => n11906, B2 => 
                           n11641, C1 => n13220, C2 => n11640, ZN => n11923);
   U615 : INV_X1 port map( A => n11923, ZN => n13128);
   U616 : INV_X1 port map( A => n13221, ZN => n13100);
   U617 : OAI22_X1 port map( A1 => n13138, A2 => n13130, B1 => n13128, B2 => 
                           n13100, ZN => n11642);
   U618 : AOI211_X1 port map( C1 => n1872, C2 => n11921, A => n11643, B => 
                           n11642, ZN => n1855);
   U619 : INV_X1 port map( A => n1867, ZN => n4476);
   U620 : NAND2_X1 port map( A1 => n4476, A2 => n11644, ZN => n7759);
   U621 : INV_X1 port map( A => n7759, ZN => n1868);
   U622 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_64_port, ZN => 
                           n1825);
   U623 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_63_port, ZN => 
                           n1824);
   U624 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_62_port, ZN => 
                           n1823);
   U625 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_61_port, ZN => 
                           n1822);
   U626 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_60_port, ZN => 
                           n1820);
   U627 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_59_port, ZN => 
                           n1819);
   U628 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_34_port, ZN => 
                           n1818);
   U629 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_33_port, ZN => 
                           n1817);
   U630 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_32_port, ZN => 
                           n1816);
   U631 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_31_port, ZN => 
                           n1815);
   U632 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_30_port, ZN => 
                           n1814);
   U633 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_29_port, ZN => 
                           n1813);
   U634 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_28_port, ZN => 
                           n1812);
   U635 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_27_port, ZN => 
                           n1811);
   U636 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n12268);
   U637 : NOR2_X1 port map( A1 => n12268, A2 => n12259, ZN => n12257);
   U638 : OAI21_X1 port map( B1 => n11647, B2 => n12257, A => n11646, ZN => 
                           n6106);
   U639 : OAI21_X1 port map( B1 => n11646, B2 => n11645, A => n1803, ZN => 
                           n11649);
   U640 : INV_X1 port map( A => n1804, ZN => n12269);
   U641 : OAI211_X1 port map( C1 => n11647, C2 => n11646, A => n12269, B => 
                           n6106, ZN => n11648);
   U642 : OAI21_X1 port map( B1 => n1801, B2 => n11649, A => n11648, ZN => 
                           n6888);
   U643 : NAND3_X1 port map( A1 => n11650, A2 => FUNC(2), A3 => FUNC(3), ZN => 
                           n12530);
   U644 : INV_X1 port map( A => n12530, ZN => n12519);
   U645 : NOR2_X1 port map( A1 => n12519, A2 => n12518, ZN => n12496);
   U646 : INV_X1 port map( A => DATA2(22), ZN => n12766);
   U647 : NOR3_X1 port map( A1 => n12496, A2 => n12766, A3 => n12554, ZN => 
                           n3862);
   U648 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_5_port,
                           ZN => n13085);
   U649 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n13085, ZN => n2808);
   U650 : AOI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n2808, ZN => n3933);
   U651 : NOR3_X1 port map( A1 => n9172, A2 => n8900, A3 => n1826, ZN => n3026)
                           ;
   U652 : AOI221_X1 port map( B1 => n8900, B2 => n9172, C1 => n1826, C2 => 
                           n9172, A => n3026, ZN => n4280);
   U653 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_3_6_port, ZN => 
                           n11651);
   U654 : NOR3_X1 port map( A1 => n8886, A2 => n1826, A3 => n11651, ZN => n3030
                           );
   U655 : AOI221_X1 port map( B1 => n8886, B2 => n11651, C1 => n1826, C2 => 
                           n11651, A => n3030, ZN => n4274);
   U656 : NAND2_X1 port map( A1 => n8978, A2 => n11306, ZN => n11652);
   U657 : OAI21_X1 port map( B1 => n8978, B2 => n11306, A => n11652, ZN => 
                           n12891);
   U658 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_4_8_port, ZN => 
                           n11653);
   U659 : NOR3_X1 port map( A1 => n1826, A2 => n12891, A3 => n11653, ZN => 
                           n3029);
   U660 : INV_X1 port map( A => n12891, ZN => n12892);
   U661 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n12892, ZN => n11654
                           );
   U662 : AOI21_X1 port map( B1 => n11654, B2 => n11653, A => n3029, ZN => 
                           n4270);
   U663 : NAND2_X1 port map( A1 => n8980, A2 => n11307, ZN => n11655);
   U664 : OAI21_X1 port map( B1 => n8980, B2 => n11307, A => n11655, ZN => 
                           n12930);
   U665 : NOR3_X1 port map( A1 => n11310, A2 => n11333, A3 => n12930, ZN => 
                           n3028);
   U666 : AOI221_X1 port map( B1 => n11310, B2 => n11333, C1 => n12930, C2 => 
                           n11333, A => n3028, ZN => n4266);
   U667 : NAND2_X1 port map( A1 => n8984, A2 => n11308, ZN => n11656);
   U668 : OAI21_X1 port map( B1 => n8984, B2 => n11308, A => n11656, ZN => 
                           n12969);
   U669 : NOR3_X1 port map( A1 => n11300, A2 => n11334, A3 => n12969, ZN => 
                           n3027);
   U670 : AOI221_X1 port map( B1 => n11300, B2 => n11334, C1 => n12969, C2 => 
                           n11334, A => n3027, ZN => n4263);
   U671 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n13060);
   U672 : INV_X1 port map( A => n13060, ZN => n13064);
   U673 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN 
                           => n12788);
   U674 : NAND2_X1 port map( A1 => n12788, A2 => data2_mul_1_port, ZN => n13058
                           );
   U675 : INV_X1 port map( A => n13058, ZN => n13063);
   U676 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => n12788, ZN => n13045)
                           ;
   U677 : AOI222_X1 port map( A1 => n13064, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           n13063, B2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, C1 => 
                           n13045, C2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, ZN => 
                           n11658);
   U678 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n12827);
   U679 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n12827, ZN => n12789);
   U680 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n12789, ZN => n11657
                           );
   U681 : NOR2_X1 port map( A1 => n11658, A2 => n11657, ZN => n3036);
   U682 : AOI21_X1 port map( B1 => n11658, B2 => n11657, A => n3036, ZN => 
                           n4257);
   U683 : INV_X1 port map( A => DATA2(9), ZN => n12779);
   U684 : NAND2_X1 port map( A1 => n12779, A2 => DATA1(9), ZN => n12636);
   U685 : NAND2_X1 port map( A1 => DATA2(9), A2 => n11659, ZN => n12659);
   U686 : NAND2_X1 port map( A1 => n12636, A2 => n12659, ZN => n12561);
   U687 : AOI22_X1 port map( A1 => n12535, A2 => n12561, B1 => n13224, B2 => 
                           n8757, ZN => n3932);
   U688 : NOR2_X1 port map( A1 => n11660, A2 => n11664, ZN => n12516);
   U689 : AOI211_X1 port map( C1 => n11660, C2 => n11664, A => n12516, B => 
                           n12434, ZN => n3920);
   U690 : NAND2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n11663
                           );
   U691 : NAND2_X1 port map( A1 => n12756, A2 => n11661, ZN => n12510);
   U692 : AOI211_X1 port map( C1 => n11664, C2 => n11663, A => n11662, B => 
                           n12510, ZN => n3919);
   U693 : INV_X1 port map( A => n12496, ZN => n12477);
   U694 : NAND3_X1 port map( A1 => DATA1(9), A2 => DATA2(9), A3 => n12477, ZN 
                           => n3918);
   U695 : INV_X1 port map( A => DATA1(30), ZN => n12586);
   U696 : NAND2_X1 port map( A1 => DATA1(27), A2 => n12332, ZN => n11665);
   U697 : NAND2_X1 port map( A1 => DATA1(28), A2 => n12216, ZN => n11918);
   U698 : OAI211_X1 port map( C1 => n11895, C2 => n12586, A => n11665, B => 
                           n11918, ZN => n11666);
   U699 : AOI211_X1 port map( C1 => n12179, C2 => DATA1(29), A => n11667, B => 
                           n11666, ZN => n6880);
   U700 : NAND2_X1 port map( A1 => DATA1(26), A2 => n12179, ZN => n11912);
   U701 : INV_X1 port map( A => DATA1(27), ZN => n12239);
   U702 : NOR2_X1 port map( A1 => n12239, A2 => n11895, ZN => n11938);
   U703 : INV_X1 port map( A => n11938, ZN => n11668);
   U704 : OAI211_X1 port map( C1 => n12163, C2 => n12700, A => n11912, B => 
                           n11668, ZN => n11669);
   U705 : AOI211_X1 port map( C1 => n12216, C2 => DATA1(25), A => n11670, B => 
                           n11669, ZN => n11677);
   U706 : OAI222_X1 port map( A1 => n12237, A2 => n11671, B1 => n11906, B2 => 
                           n11678, C1 => n13220, C2 => n11677, ZN => n6187);
   U707 : NOR2_X1 port map( A1 => n12239, A2 => n12232, ZN => n11916);
   U708 : INV_X1 port map( A => DATA1(28), ZN => n12710);
   U709 : NAND2_X1 port map( A1 => DATA1(24), A2 => n12541, ZN => n11673);
   U710 : OAI211_X1 port map( C1 => n11895, C2 => n12710, A => n11673, B => 
                           n11672, ZN => n11674);
   U711 : AOI211_X1 port map( C1 => n12216, C2 => DATA1(26), A => n11916, B => 
                           n11674, ZN => n1839);
   U712 : NAND2_X1 port map( A1 => DATA1(27), A2 => n12216, ZN => n11911);
   U713 : NAND2_X1 port map( A1 => DATA1(26), A2 => n12332, ZN => n11891);
   U714 : OAI211_X1 port map( C1 => n12232, C2 => n12710, A => n11911, B => 
                           n11891, ZN => n11675);
   U715 : AOI211_X1 port map( C1 => DATA1(29), C2 => n11917, A => n11676, B => 
                           n11675, ZN => n6179);
   U716 : OAI222_X1 port map( A1 => n12237, A2 => n11677, B1 => n11906, B2 => 
                           n1839, C1 => n13220, C2 => n6179, ZN => n6938);
   U717 : INV_X1 port map( A => n11677, ZN => n11680);
   U718 : OAI22_X1 port map( A1 => n11678, A2 => n12237, B1 => n1839, B2 => 
                           n13220, ZN => n11679);
   U719 : AOI21_X1 port map( B1 => n1865, B2 => n11680, A => n11679, ZN => 
                           n6184);
   U720 : AOI22_X1 port map( A1 => n1872, A2 => n11681, B1 => n13123, B2 => 
                           n6198, ZN => n6177);
   U721 : OAI22_X1 port map( A1 => n13138, A2 => n11682, B1 => n1845, B2 => 
                           n11315, ZN => n6192);
   U722 : AOI222_X1 port map( A1 => n11685, A2 => n11781, B1 => n11684, B2 => 
                           n13223, C1 => n11683, C2 => n11844, ZN => n6206);
   U723 : OAI22_X1 port map( A1 => n1869, A2 => n13137, B1 => n6206, B2 => 
                           n13133, ZN => n6191);
   U724 : INV_X1 port map( A => n1849, ZN => n11691);
   U725 : OAI22_X1 port map( A1 => n13138, A2 => n11691, B1 => n13137, B2 => 
                           n11315, ZN => n6197);
   U726 : OAI22_X1 port map( A1 => n1845, A2 => n13133, B1 => n6206, B2 => 
                           n13135, ZN => n6196);
   U727 : AOI22_X1 port map( A1 => n1872, A2 => n11694, B1 => n13221, B2 => 
                           n11699, ZN => n6205);
   U728 : NOR2_X1 port map( A1 => n12470, A2 => n12341, ZN => n11688);
   U729 : NAND2_X1 port map( A1 => DATA1(15), A2 => n12216, ZN => n11873);
   U730 : OAI211_X1 port map( C1 => n11895, C2 => n12402, A => n11686, B => 
                           n11873, ZN => n11687);
   U731 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(16), A => n11688, B => 
                           n11687, ZN => n11696);
   U732 : INV_X1 port map( A => n11693, ZN => n11690);
   U733 : OAI222_X1 port map( A1 => n12237, A2 => n11696, B1 => n11906, B2 => 
                           n11690, C1 => n13220, C2 => n11689, ZN => n11700);
   U734 : AOI22_X1 port map( A1 => n13123, A2 => n1849, B1 => n13222, B2 => 
                           n11700, ZN => n6204);
   U735 : OAI22_X1 port map( A1 => n6206, A2 => n11315, B1 => n11691, B2 => 
                           n13133, ZN => n6207);
   U736 : AOI22_X1 port map( A1 => n13123, A2 => n11699, B1 => n13121, B2 => 
                           n11694, ZN => n6213);
   U737 : OAI22_X1 port map( A1 => n11696, A2 => n11906, B1 => n11697, B2 => 
                           n12237, ZN => n11692);
   U738 : AOI21_X1 port map( B1 => n11781, B2 => n11693, A => n11692, ZN => 
                           n11718);
   U739 : INV_X1 port map( A => n11718, ZN => n11701);
   U740 : AOI22_X1 port map( A1 => n1872, A2 => n11700, B1 => n13221, B2 => 
                           n11701, ZN => n6212);
   U741 : AOI22_X1 port map( A1 => n1872, A2 => n11699, B1 => n13123, B2 => 
                           n11694, ZN => n6215);
   U742 : AOI22_X1 port map( A1 => n13221, A2 => n11700, B1 => n13222, B2 => 
                           n11701, ZN => n6214);
   U743 : INV_X1 port map( A => n11695, ZN => n11698);
   U744 : OAI222_X1 port map( A1 => n12237, A2 => n11698, B1 => n11906, B2 => 
                           n11697, C1 => n13220, C2 => n11696, ZN => n1852);
   U745 : AOI22_X1 port map( A1 => n1872, A2 => n1852, B1 => n13221, B2 => 
                           n1853, ZN => n6238);
   U746 : AOI22_X1 port map( A1 => n13123, A2 => n11701, B1 => n13121, B2 => 
                           n11700, ZN => n6237);
   U747 : AOI22_X1 port map( A1 => n13221, A2 => n1852, B1 => n13121, B2 => 
                           n11699, ZN => n6241);
   U748 : AOI22_X1 port map( A1 => n1872, A2 => n11701, B1 => n13123, B2 => 
                           n11700, ZN => n6240);
   U749 : NOR2_X1 port map( A1 => n12588, A2 => n12545, ZN => n11702);
   U750 : NOR2_X1 port map( A1 => n11895, A2 => n11764, ZN => n12339);
   U751 : AOI211_X1 port map( C1 => n12541, C2 => DATA1(9), A => n11702, B => 
                           n12339, ZN => n11703);
   U752 : NAND2_X1 port map( A1 => DATA1(6), A2 => n12179, ZN => n11833);
   U753 : OAI211_X1 port map( C1 => n12163, C2 => n12656, A => n11703, B => 
                           n11833, ZN => n11930);
   U754 : NOR2_X1 port map( A1 => n12656, A2 => n12341, ZN => n11704);
   U755 : NOR2_X1 port map( A1 => n11895, A2 => n11803, ZN => n12540);
   U756 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(5), A => n11704, B => 
                           n12540, ZN => n11706);
   U757 : NAND2_X1 port map( A1 => DATA1(6), A2 => n12216, ZN => n11705);
   U758 : OAI211_X1 port map( C1 => n12163, C2 => n12588, A => n11706, B => 
                           n11705, ZN => n11928);
   U759 : NOR2_X1 port map( A1 => n11764, A2 => n12545, ZN => n11709);
   U760 : NOR2_X1 port map( A1 => n11803, A2 => n12232, ZN => n12338);
   U761 : INV_X1 port map( A => n12338, ZN => n11707);
   U762 : NAND2_X1 port map( A1 => DATA1(7), A2 => n12541, ZN => n11745);
   U763 : OAI211_X1 port map( C1 => n11895, C2 => n9206, A => n11707, B => 
                           n11745, ZN => n11708);
   U764 : AOI211_X1 port map( C1 => n12332, C2 => DATA1(6), A => n11709, B => 
                           n11708, ZN => n11710);
   U765 : INV_X1 port map( A => n11710, ZN => n11712);
   U766 : AOI222_X1 port map( A1 => n13223, A2 => n11930, B1 => n1865, B2 => 
                           n11928, C1 => n11781, C2 => n11712, ZN => n11949);
   U767 : OAI22_X1 port map( A1 => n13138, A2 => n11949, B1 => n1830, B2 => 
                           n11315, ZN => n6261);
   U768 : AOI222_X1 port map( A1 => n11711, A2 => n11781, B1 => n11928, B2 => 
                           n13223, C1 => n11712, C2 => n11844, ZN => n11947);
   U769 : AOI222_X1 port map( A1 => n11760, A2 => n11781, B1 => n11712, B2 => 
                           n13223, C1 => n11711, C2 => n11844, ZN => n11948);
   U770 : OAI22_X1 port map( A1 => n11947, A2 => n13100, B1 => n11948, B2 => 
                           n13133, ZN => n6260);
   U771 : OAI222_X1 port map( A1 => n8677, A2 => n12523, B1 => n8801, B2 => 
                           n11796, C1 => n9166, C2 => n12524, ZN => n11713);
   U772 : AOI211_X1 port map( C1 => n8902, C2 => n11713, A => n8674, B => n8673
                           , ZN => n11715);
   U773 : OAI21_X1 port map( B1 => n8651, B2 => n8650, A => n8969, ZN => n11714
                           );
   U774 : NAND4_X1 port map( A1 => n8675, A2 => n8859, A3 => n11715, A4 => 
                           n11714, ZN => OUTALU(9));
   U775 : INV_X1 port map( A => DATA2(8), ZN => n12780);
   U776 : OAI22_X1 port map( A1 => n12780, A2 => DATA1(8), B1 => n12656, B2 => 
                           DATA2(8), ZN => n12599);
   U777 : AOI22_X1 port map( A1 => n8875, A2 => n13224, B1 => n12535, B2 => 
                           n12599, ZN => n3911);
   U778 : NAND3_X1 port map( A1 => DATA1(8), A2 => DATA2(8), A3 => n12477, ZN 
                           => n3910);
   U779 : OAI222_X1 port map( A1 => n13100, A2 => n11948, B1 => n13133, B2 => 
                           n1830, C1 => n11947, C2 => n13108, ZN => n6268);
   U780 : INV_X1 port map( A => n11717, ZN => n11716);
   U781 : AOI22_X1 port map( A1 => n11717, A2 => n12510, B1 => n12434, B2 => 
                           n11716, ZN => n6267);
   U782 : OAI22_X1 port map( A1 => n1869, A2 => n11718, B1 => n11751, B2 => 
                           n13133, ZN => n11725);
   U783 : NOR2_X1 port map( A1 => n11895, A2 => n12668, ZN => n11720);
   U784 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(11), A => n11720, B => 
                           n11719, ZN => n11722);
   U785 : NAND2_X1 port map( A1 => DATA1(9), A2 => n12332, ZN => n11721);
   U786 : OAI211_X1 port map( C1 => n12341, C2 => n12656, A => n11722, B => 
                           n11721, ZN => n11783);
   U787 : AOI222_X1 port map( A1 => n11723, A2 => n11781, B1 => n11783, B2 => 
                           n12182, C1 => n11750, C2 => n11844, ZN => n13119);
   U788 : OAI22_X1 port map( A1 => n13138, A2 => n13119, B1 => n6351, B2 => 
                           n13135, ZN => n11724);
   U789 : AOI211_X1 port map( C1 => n13123, C2 => n1852, A => n11725, B => 
                           n11724, ZN => n6381);
   U790 : AOI211_X1 port map( C1 => n8539, C2 => n8969, A => n8648, B => n13214
                           , ZN => n11729);
   U791 : OAI22_X1 port map( A1 => n8677, A2 => n12524, B1 => n9166, B2 => 
                           n11796, ZN => n11727);
   U792 : OAI22_X1 port map( A1 => n11818, A2 => n8801, B1 => n9167, B2 => 
                           n12523, ZN => n11726);
   U793 : OAI21_X1 port map( B1 => n11727, B2 => n11726, A => n8902, ZN => 
                           n11728);
   U794 : NAND3_X1 port map( A1 => n8649, A2 => n11729, A3 => n11728, ZN => 
                           OUTALU(8));
   U795 : NAND2_X1 port map( A1 => n12756, A2 => n9220, ZN => n12327);
   U796 : INV_X1 port map( A => n12327, ZN => n12533);
   U797 : INV_X1 port map( A => n11730, ZN => n11734);
   U798 : INV_X1 port map( A => n12328, ZN => n11731);
   U799 : AOI21_X1 port map( B1 => n11733, B2 => n11731, A => n12171, ZN => 
                           n12169);
   U800 : NOR2_X1 port map( A1 => n11734, A2 => n12169, ZN => n11831);
   U801 : INV_X1 port map( A => n11732, ZN => n13068);
   U802 : NOR2_X1 port map( A1 => n11831, A2 => n13068, ZN => n11830);
   U803 : NOR2_X1 port map( A1 => n11735, A2 => n11830, ZN => n11808);
   U804 : OAI21_X1 port map( B1 => n11808, B2 => n1429, A => n11736, ZN => 
                           n11767);
   U805 : AOI21_X1 port map( B1 => n11772, B2 => n11767, A => n11737, ZN => 
                           n11758);
   U806 : OAI21_X1 port map( B1 => n11758, B2 => n1353, A => n11738, ZN => 
                           n11741);
   U807 : INV_X1 port map( A => n12333, ZN => n12335);
   U808 : INV_X1 port map( A => n11733, ZN => n12168);
   U809 : AOI21_X1 port map( B1 => n12532, B2 => n12335, A => n12168, ZN => 
                           n12167);
   U810 : NOR2_X1 port map( A1 => n12167, A2 => n12171, ZN => n12166);
   U811 : NOR2_X1 port map( A1 => n11734, A2 => n12166, ZN => n13069);
   U812 : NOR2_X1 port map( A1 => n13069, A2 => n13068, ZN => n13067);
   U813 : NOR2_X1 port map( A1 => n11735, A2 => n13067, ZN => n11807);
   U814 : OAI21_X1 port map( B1 => n11807, B2 => n1429, A => n11736, ZN => 
                           n11766);
   U815 : AOI21_X1 port map( B1 => n11772, B2 => n11766, A => n11737, ZN => 
                           n11757);
   U816 : OAI21_X1 port map( B1 => n11757, B2 => n1353, A => n11738, ZN => 
                           n11740);
   U817 : AOI22_X1 port map( A1 => n12533, A2 => n11741, B1 => n7166, B2 => 
                           n11740, ZN => n11739);
   U818 : NOR2_X1 port map( A1 => n11743, A2 => n11739, ZN => n4220);
   U819 : INV_X1 port map( A => n12518, ZN => n12466);
   U820 : OAI221_X1 port map( B1 => DATA1(7), B2 => n1835, C1 => n12588, C2 => 
                           n12530, A => n12466, ZN => n11744);
   U821 : INV_X1 port map( A => n7166, ZN => n12165);
   U822 : OAI22_X1 port map( A1 => n12327, A2 => n11741, B1 => n12165, B2 => 
                           n11740, ZN => n11742);
   U823 : AOI22_X1 port map( A1 => DATA2(7), A2 => n11744, B1 => n11743, B2 => 
                           n11742, ZN => n6314);
   U824 : OAI22_X1 port map( A1 => n13138, A2 => n11948, B1 => n1830, B2 => 
                           n13135, ZN => n6294);
   U825 : INV_X1 port map( A => DATA1(11), ZN => n12497);
   U826 : INV_X1 port map( A => n11745, ZN => n11746);
   U827 : AOI211_X1 port map( C1 => n12332, C2 => DATA1(8), A => n11747, B => 
                           n11746, ZN => n11749);
   U828 : OAI211_X1 port map( C1 => n11895, C2 => n12497, A => n11749, B => 
                           n11748, ZN => n11782);
   U829 : AOI222_X1 port map( A1 => n11750, A2 => n11781, B1 => n11782, B2 => 
                           n12182, C1 => n11783, C2 => n11844, ZN => n13126);
   U830 : OAI22_X1 port map( A1 => n13138, A2 => n13126, B1 => n6351, B2 => 
                           n13133, ZN => n11753);
   U831 : OAI22_X1 port map( A1 => n13119, A2 => n13100, B1 => n11751, B2 => 
                           n11315, ZN => n11752);
   U832 : AOI211_X1 port map( C1 => n13121, C2 => n1852, A => n11753, B => 
                           n11752, ZN => n6422);
   U833 : OR2_X1 port map( A1 => n9163, A2 => n9100, ZN => n11755);
   U834 : AOI211_X1 port map( C1 => n8645, C2 => n8969, A => n8959, B => n9174,
                           ZN => n11754);
   U835 : OAI211_X1 port map( C1 => n11800, C2 => n11755, A => n8646, B => 
                           n11754, ZN => OUTALU(7));
   U836 : AOI22_X1 port map( A1 => n12533, A2 => n11758, B1 => n7166, B2 => 
                           n11757, ZN => n3905);
   U837 : AOI22_X1 port map( A1 => DATA2(6), A2 => n12651, B1 => DATA1(6), B2 
                           => n12784, ZN => n12655);
   U838 : AOI21_X1 port map( B1 => n12519, B2 => DATA1(6), A => n12518, ZN => 
                           n11756);
   U839 : OAI22_X1 port map( A1 => n12655, A2 => n1835, B1 => n11756, B2 => 
                           n12784, ZN => n3904);
   U840 : OAI22_X1 port map( A1 => n11758, A2 => n12327, B1 => n11757, B2 => 
                           n12165, ZN => n11759);
   U841 : NAND2_X1 port map( A1 => n1353, A2 => n11759, ZN => n6340);
   U842 : OAI21_X1 port map( B1 => n12530, B2 => n11764, A => n12466, ZN => 
                           n11763);
   U843 : INV_X1 port map( A => n1834, ZN => n12331);
   U844 : AOI22_X1 port map( A1 => n11760, A2 => n13223, B1 => n11802, B2 => 
                           n1865, ZN => n11761);
   U845 : INV_X1 port map( A => n11761, ZN => n11762);
   U846 : AOI22_X1 port map( A1 => DATA2(5), A2 => n11763, B1 => n12331, B2 => 
                           n11762, ZN => n3902);
   U847 : NOR2_X1 port map( A1 => n11764, A2 => DATA2(5), ZN => n12597);
   U848 : NOR2_X1 port map( A1 => DATA1(5), A2 => n12785, ZN => n12650);
   U849 : NOR2_X1 port map( A1 => n12597, A2 => n12650, ZN => n12573);
   U850 : INV_X1 port map( A => n12573, ZN => n11765);
   U851 : AOI22_X1 port map( A1 => n12535, A2 => n11765, B1 => n13224, B2 => 
                           n8773, ZN => n3900);
   U852 : OAI22_X1 port map( A1 => n12327, A2 => n11767, B1 => n12165, B2 => 
                           n11766, ZN => n11771);
   U853 : AOI22_X1 port map( A1 => n11767, A2 => n12533, B1 => n11766, B2 => 
                           n7166, ZN => n11768);
   U854 : INV_X1 port map( A => n11768, ZN => n11770);
   U855 : AOI22_X1 port map( A1 => n11772, A2 => n11771, B1 => n11770, B2 => 
                           n11769, ZN => n6367);
   U856 : INV_X1 port map( A => n6351, ZN => n13122);
   U857 : AOI211_X1 port map( C1 => n12332, C2 => DATA1(6), A => n11774, B => 
                           n11773, ZN => n11776);
   U858 : OAI211_X1 port map( C1 => n12545, C2 => n12588, A => n11776, B => 
                           n11775, ZN => n11845);
   U859 : AOI211_X1 port map( C1 => DATA1(10), C2 => n11917, A => n11778, B => 
                           n11777, ZN => n11780);
   U860 : OAI211_X1 port map( C1 => n12163, C2 => n12588, A => n11780, B => 
                           n11779, ZN => n11846);
   U861 : AOI222_X1 port map( A1 => n11782, A2 => n11781, B1 => n11845, B2 => 
                           n12182, C1 => n11846, C2 => n11844, ZN => n13101);
   U862 : AOI222_X1 port map( A1 => n11783, A2 => n11781, B1 => n11846, B2 => 
                           n12182, C1 => n11782, C2 => n1865, ZN => n13118);
   U863 : OAI22_X1 port map( A1 => n13138, A2 => n13101, B1 => n13118, B2 => 
                           n13135, ZN => n11785);
   U864 : OAI22_X1 port map( A1 => n13119, A2 => n11315, B1 => n13126, B2 => 
                           n13133, ZN => n11784);
   U865 : AOI211_X1 port map( C1 => n13121, C2 => n13122, A => n11785, B => 
                           n11784, ZN => n6980);
   U866 : INV_X1 port map( A => n11786, ZN => n11795);
   U867 : OAI22_X1 port map( A1 => n13139, A2 => n8644, B1 => n8647, B2 => 
                           n9021, ZN => n11787);
   U868 : INV_X1 port map( A => n11787, ZN => n11790);
   U869 : AOI22_X1 port map( A1 => n11788, A2 => n13151, B1 => n13141, B2 => 
                           n13187, ZN => n11789);
   U870 : OAI211_X1 port map( C1 => n9104, C2 => n8641, A => n11790, B => 
                           n11789, ZN => n11852);
   U871 : AOI222_X1 port map( A1 => n11791, A2 => n9008, B1 => n11852, B2 => 
                           n9011, C1 => n11812, C2 => n8907, ZN => n12349);
   U872 : OAI22_X1 port map( A1 => n11792, A2 => n13148, B1 => n12349, B2 => 
                           n13143, ZN => n11794);
   U873 : OAI22_X1 port map( A1 => n11813, A2 => n8561, B1 => n11814, B2 => 
                           n13150, ZN => n11793);
   U874 : AOI211_X1 port map( C1 => n9102, C2 => n11795, A => n11794, B => 
                           n11793, ZN => n12357);
   U875 : INV_X1 port map( A => n12357, ZN => n12194);
   U876 : AOI22_X1 port map( A1 => n12194, A2 => n9010, B1 => n11857, B2 => 
                           n13178, ZN => n11799);
   U877 : OAI22_X1 port map( A1 => n11818, A2 => n9167, B1 => n9101, B2 => 
                           n11796, ZN => n11797);
   U878 : INV_X1 port map( A => n11797, ZN => n11798);
   U879 : OAI211_X1 port map( C1 => n12197, C2 => n9166, A => n11799, B => 
                           n11798, ZN => n11860);
   U880 : INV_X1 port map( A => n11860, ZN => n11822);
   U881 : OAI222_X1 port map( A1 => n9219, A2 => n11800, B1 => n11823, B2 => 
                           n8908, C1 => n9163, C2 => n11822, ZN => n12362);
   U882 : INV_X1 port map( A => n12362, ZN => n12186);
   U883 : OR3_X1 port map( A1 => n12186, A2 => n8802, A3 => n9100, ZN => n11801
                           );
   U884 : NAND4_X1 port map( A1 => n8638, A2 => n8640, A3 => n8639, A4 => 
                           n11801, ZN => OUTALU(5));
   U885 : AOI22_X1 port map( A1 => n12533, A2 => n11808, B1 => n7166, B2 => 
                           n11807, ZN => n3897);
   U886 : AND3_X1 port map( A1 => n11802, A2 => n13223, A3 => n12331, ZN => 
                           n11806);
   U887 : AOI21_X1 port map( B1 => n12519, B2 => DATA1(4), A => n12518, ZN => 
                           n11804);
   U888 : INV_X1 port map( A => DATA2(4), ZN => n13076);
   U889 : NAND2_X1 port map( A1 => DATA2(4), A2 => n11803, ZN => n12644);
   U890 : NAND2_X1 port map( A1 => DATA1(4), A2 => n13076, ZN => n12648);
   U891 : AND2_X1 port map( A1 => n12644, A2 => n12648, ZN => n12565);
   U892 : OAI22_X1 port map( A1 => n11804, A2 => n13076, B1 => n12565, B2 => 
                           n1835, ZN => n11805);
   U893 : AOI211_X1 port map( C1 => n13224, C2 => n8555, A => n11806, B => 
                           n11805, ZN => n3896);
   U894 : OAI22_X1 port map( A1 => n11808, A2 => n12327, B1 => n11807, B2 => 
                           n12165, ZN => n3895);
   U895 : AOI22_X1 port map( A1 => n8906, A2 => n8633, B1 => n13188, B2 => 
                           n13146, ZN => n11811);
   U896 : OAI22_X1 port map( A1 => n8647, A2 => n8895, B1 => n9181, B2 => n8637
                           , ZN => n11809);
   U897 : INV_X1 port map( A => n11809, ZN => n11810);
   U898 : OAI211_X1 port map( C1 => n9165, C2 => n8641, A => n11811, B => 
                           n11810, ZN => n12187);
   U899 : AOI222_X1 port map( A1 => n11812, A2 => n9008, B1 => n12187, B2 => 
                           n9011, C1 => n11852, C2 => n8907, ZN => n12353);
   U900 : OAI22_X1 port map( A1 => n12353, A2 => n13189, B1 => n12349, B2 => 
                           n13148, ZN => n11816);
   U901 : OAI22_X1 port map( A1 => n11814, A2 => n9217, B1 => n11813, B2 => 
                           n13150, ZN => n11815);
   U902 : AOI211_X1 port map( C1 => n9025, C2 => n12191, A => n11816, B => 
                           n11815, ZN => n12737);
   U903 : INV_X1 port map( A => n12737, ZN => n12354);
   U904 : AOI22_X1 port map( A1 => n12194, A2 => n8899, B1 => n12354, B2 => 
                           n13166, ZN => n11821);
   U905 : OAI22_X1 port map( A1 => n11818, A2 => n9101, B1 => n11817, B2 => 
                           n9167, ZN => n11819);
   U906 : INV_X1 port map( A => n11819, ZN => n11820);
   U907 : OAI211_X1 port map( C1 => n12197, C2 => n8677, A => n11821, B => 
                           n11820, ZN => n12198);
   U908 : INV_X1 port map( A => n12198, ZN => n11824);
   U909 : OAI222_X1 port map( A1 => n11824, A2 => n9163, B1 => n9219, B2 => 
                           n11823, C1 => n11822, C2 => n8908, ZN => n12747);
   U910 : INV_X1 port map( A => n12747, ZN => n12359);
   U911 : OAI22_X1 port map( A1 => n8805, A2 => n12186, B1 => n12359, B2 => 
                           n8802, ZN => n11825);
   U912 : AOI22_X1 port map( A1 => n8902, A2 => n11825, B1 => n8634, B2 => 
                           n8894, ZN => n11826);
   U913 : OAI211_X1 port map( C1 => n8894, C2 => n8636, A => n8635, B => n11826
                           , ZN => OUTALU(4));
   U914 : NAND2_X1 port map( A1 => n13078, A2 => n9225, ZN => n12589);
   U915 : NAND2_X1 port map( A1 => DATA2(3), A2 => n13149, ZN => n12643);
   U916 : NAND2_X1 port map( A1 => n12589, A2 => n12643, ZN => n12557);
   U917 : NOR2_X1 port map( A1 => n9205, A2 => n12163, ZN => n12336);
   U918 : AOI21_X1 port map( B1 => n12215, B2 => n9221, A => n12336, ZN => 
                           n11827);
   U919 : NAND2_X1 port map( A1 => n9225, A2 => n12541, ZN => n11834);
   U920 : OAI211_X1 port map( C1 => n11332, C2 => n12545, A => n11827, B => 
                           n11834, ZN => n11828);
   U921 : AOI22_X1 port map( A1 => n12535, A2 => n12557, B1 => n12331, B2 => 
                           n11828, ZN => n3894);
   U922 : OAI21_X1 port map( B1 => n9206, B2 => n12530, A => n12466, ZN => 
                           n11829);
   U923 : AOI22_X1 port map( A1 => DATA2(3), A2 => n11829, B1 => n13224, B2 => 
                           n8793, ZN => n3893);
   U924 : AOI21_X1 port map( B1 => n13068, B2 => n11831, A => n11830, ZN => 
                           n11832);
   U925 : NAND2_X1 port map( A1 => n12533, A2 => n11832, ZN => n3892);
   U926 : OAI211_X1 port map( C1 => n11895, C2 => n12588, A => n11834, B => 
                           n11833, ZN => n11835);
   U927 : AOI211_X1 port map( C1 => n12216, C2 => DATA1(5), A => n11836, B => 
                           n11835, ZN => n11837);
   U928 : INV_X1 port map( A => n11837, ZN => n12342);
   U929 : OAI211_X1 port map( C1 => n11895, C2 => n12656, A => n11839, B => 
                           n11838, ZN => n11840);
   U930 : AOI211_X1 port map( C1 => n12216, C2 => DATA1(6), A => n11841, B => 
                           n11840, ZN => n11842);
   U931 : INV_X1 port map( A => n11842, ZN => n12183);
   U932 : AOI222_X1 port map( A1 => n12182, A2 => n12342, B1 => n1865, B2 => 
                           n12183, C1 => n11781, C2 => n11845, ZN => n11843);
   U933 : INV_X1 port map( A => n11843, ZN => n12553);
   U934 : AOI222_X1 port map( A1 => n11846, A2 => n11781, B1 => n12183, B2 => 
                           n12182, C1 => n11845, C2 => n11844, ZN => n13102);
   U935 : OAI22_X1 port map( A1 => n13118, A2 => n11315, B1 => n13102, B2 => 
                           n13135, ZN => n11848);
   U936 : OAI22_X1 port map( A1 => n1869, A2 => n13126, B1 => n13101, B2 => 
                           n13133, ZN => n11847);
   U937 : AOI211_X1 port map( C1 => n13222, C2 => n12553, A => n11848, B => 
                           n11847, ZN => n7287);
   U938 : OAI22_X1 port map( A1 => n9020, A2 => n8641, B1 => n13142, B2 => 
                           n13158, ZN => n11850);
   U939 : OAI22_X1 port map( A1 => n9182, A2 => n8630, B1 => n9165, B2 => n8637
                           , ZN => n11849);
   U940 : AOI211_X1 port map( C1 => n13151, C2 => n13188, A => n11850, B => 
                           n11849, ZN => n12347);
   U941 : INV_X1 port map( A => n12347, ZN => n11851);
   U942 : AOI222_X1 port map( A1 => n8907, A2 => n12187, B1 => n13183, B2 => 
                           n11852, C1 => n11851, C2 => n13159, ZN => n12730);
   U943 : INV_X1 port map( A => n12730, ZN => n12348);
   U944 : INV_X1 port map( A => n12353, ZN => n12727);
   U945 : AOI22_X1 port map( A1 => n9183, A2 => n12348, B1 => n8905, B2 => 
                           n12727, ZN => n11855);
   U946 : AOI22_X1 port map( A1 => n8807, A2 => n12191, B1 => n9026, B2 => 
                           n11853, ZN => n11854);
   U947 : OAI211_X1 port map( C1 => n12349, C2 => n8561, A => n11855, B => 
                           n11854, ZN => n12733);
   U948 : AOI22_X1 port map( A1 => n9164, A2 => n12733, B1 => n9173, B2 => 
                           n12194, ZN => n11859);
   U949 : AOI22_X1 port map( A1 => n8973, A2 => n11857, B1 => n8804, B2 => 
                           n11856, ZN => n11858);
   U950 : OAI211_X1 port map( C1 => n12737, C2 => n9166, A => n11859, B => 
                           n11858, ZN => n12358);
   U951 : AOI222_X1 port map( A1 => n11860, A2 => n9034, B1 => n12198, B2 => 
                           n9035, C1 => n12358, C2 => n8909, ZN => n12743);
   U952 : OAI222_X1 port map( A1 => n8805, A2 => n12359, B1 => n12186, B2 => 
                           n9113, C1 => n12743, C2 => n8802, ZN => n11861);
   U953 : AOI22_X1 port map( A1 => n8902, A2 => n11861, B1 => n9110, B2 => 
                           n8800, ZN => n11862);
   U954 : NAND4_X1 port map( A1 => n8956, A2 => n8632, A3 => n8631, A4 => 
                           n11862, ZN => OUTALU(3));
   U955 : INV_X1 port map( A => n11863, ZN => n11868);
   U956 : NOR2_X1 port map( A1 => n12613, A2 => n12545, ZN => n11867);
   U957 : NAND2_X1 port map( A1 => DATA1(14), A2 => n11917, ZN => n11865);
   U958 : OAI211_X1 port map( C1 => n12341, C2 => n12687, A => n11865, B => 
                           n11864, ZN => n11866);
   U959 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(15), A => n11867, B => 
                           n11866, ZN => n11878);
   U960 : OAI222_X1 port map( A1 => n12237, A2 => n11868, B1 => n11906, B2 => 
                           n11879, C1 => n13220, C2 => n11878, ZN => n11902);
   U961 : AOI22_X1 port map( A1 => n13123, A2 => n11882, B1 => n13121, B2 => 
                           n11902, ZN => n3885);
   U962 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n4212);
   U963 : NOR2_X1 port map( A1 => n11870, A2 => n11869, ZN => n4205);
   U964 : INV_X1 port map( A => n1847, ZN => n11890);
   U965 : OAI22_X1 port map( A1 => n13138, A2 => n1842, B1 => n1869, B2 => 
                           n1848, ZN => n11871);
   U966 : AOI21_X1 port map( B1 => n13123, B2 => n11890, A => n11871, ZN => 
                           n11872);
   U967 : OAI21_X1 port map( B1 => n13134, B2 => n13100, A => n11872, ZN => 
                           n6502);
   U968 : OAI211_X1 port map( C1 => n12163, C2 => n12613, A => n11874, B => 
                           n11873, ZN => n11875);
   U969 : AOI211_X1 port map( C1 => n12541, C2 => DATA1(17), A => n11876, B => 
                           n11875, ZN => n11907);
   U970 : INV_X1 port map( A => n11877, ZN => n11905);
   U971 : OAI222_X1 port map( A1 => n12237, A2 => n11878, B1 => n11906, B2 => 
                           n11907, C1 => n13220, C2 => n11905, ZN => n6561);
   U972 : OAI222_X1 port map( A1 => n12237, A2 => n11879, B1 => n11906, B2 => 
                           n11878, C1 => n13220, C2 => n11907, ZN => n11908);
   U973 : AOI22_X1 port map( A1 => n13221, A2 => n11882, B1 => n13123, B2 => 
                           n11908, ZN => n11881);
   U974 : AOI22_X1 port map( A1 => n1872, A2 => n11902, B1 => n13121, B2 => 
                           n6561, ZN => n11880);
   U975 : OAI211_X1 port map( C1 => n13108, C2 => n1848, A => n11881, B => 
                           n11880, ZN => n6533);
   U976 : AOI22_X1 port map( A1 => n1872, A2 => n11882, B1 => n13121, B2 => 
                           n11908, ZN => n11884);
   U977 : AOI22_X1 port map( A1 => n13123, A2 => n11902, B1 => n13222, B2 => 
                           n11890, ZN => n11883);
   U978 : OAI211_X1 port map( C1 => n1848, C2 => n13135, A => n11884, B => 
                           n11883, ZN => n6523);
   U979 : INV_X1 port map( A => n11885, ZN => n11889);
   U980 : AOI22_X1 port map( A1 => n13223, A2 => n11887, B1 => n1865, B2 => 
                           n11886, ZN => n11888);
   U981 : OAI21_X1 port map( B1 => n11889, B2 => n13220, A => n11888, ZN => 
                           n6516);
   U982 : AOI22_X1 port map( A1 => n13221, A2 => n11890, B1 => n13222, B2 => 
                           n6516, ZN => n6505);
   U983 : INV_X1 port map( A => n13134, ZN => n11901);
   U984 : AOI22_X1 port map( A1 => n13221, A2 => n6516, B1 => n13222, B2 => 
                           n11901, ZN => n6506);
   U985 : NOR2_X1 port map( A1 => n12239, A2 => n12341, ZN => n12236);
   U986 : OAI211_X1 port map( C1 => n12232, C2 => n12700, A => n11892, B => 
                           n11891, ZN => n11893);
   U987 : AOI211_X1 port map( C1 => n12216, C2 => DATA1(25), A => n12236, B => 
                           n11893, ZN => n1840);
   U988 : INV_X1 port map( A => n11894, ZN => n11900);
   U989 : OAI22_X1 port map( A1 => n11900, A2 => n11906, B1 => n1840, B2 => 
                           n12237, ZN => n6510);
   U990 : NOR2_X1 port map( A1 => n11895, A2 => n12700, ZN => n11899);
   U991 : NOR2_X1 port map( A1 => n12572, A2 => n12545, ZN => n11897);
   U992 : OAI22_X1 port map( A1 => n12710, A2 => n12341, B1 => n12239, B2 => 
                           n12163, ZN => n11896);
   U993 : NOR4_X1 port map( A1 => n11899, A2 => n11898, A3 => n11897, A4 => 
                           n11896, ZN => n11335);
   U994 : OAI222_X1 port map( A1 => n12237, A2 => n11335, B1 => n11906, B2 => 
                           n1840, C1 => n13220, C2 => n11900, ZN => n6671);
   U995 : AOI22_X1 port map( A1 => n13123, A2 => n11901, B1 => n13121, B2 => 
                           n6516, ZN => n6517);
   U996 : INV_X1 port map( A => n11902, ZN => n11909);
   U997 : OAI22_X1 port map( A1 => n13138, A2 => n11903, B1 => n11909, B2 => 
                           n13135, ZN => n6525);
   U998 : OAI222_X1 port map( A1 => n12237, A2 => n11907, B1 => n11906, B2 => 
                           n11905, C1 => n13220, C2 => n11904, ZN => n11922);
   U999 : INV_X1 port map( A => n11922, ZN => n13127);
   U1000 : INV_X1 port map( A => n11908, ZN => n13129);
   U1001 : OAI22_X1 port map( A1 => n13127, A2 => n1869, B1 => n13129, B2 => 
                           n13133, ZN => n6524);
   U1002 : OAI22_X1 port map( A1 => n13138, A2 => n11909, B1 => n13129, B2 => 
                           n13100, ZN => n6530);
   U1003 : OAI22_X1 port map( A1 => n13127, A2 => n11315, B1 => n13130, B2 => 
                           n1869, ZN => n6529);
   U1004 : NOR2_X1 port map( A1 => n12710, A2 => n12163, ZN => n12234);
   U1005 : NOR2_X1 port map( A1 => n11910, A2 => n12234, ZN => n11913);
   U1006 : NAND2_X1 port map( A1 => DATA1(29), A2 => n12541, ZN => n12204);
   U1007 : NAND4_X1 port map( A1 => n11913, A2 => n11912, A3 => n11911, A4 => 
                           n12204, ZN => n6677);
   U1008 : OAI22_X1 port map( A1 => n13128, A2 => n11315, B1 => n13130, B2 => 
                           n13133, ZN => n11915);
   U1009 : INV_X1 port map( A => n11921, ZN => n13114);
   U1010 : OAI22_X1 port map( A1 => n13127, A2 => n13100, B1 => n1869, B2 => 
                           n13114, ZN => n11914);
   U1011 : AOI211_X1 port map( C1 => n13222, C2 => n6561, A => n11915, B => 
                           n11914, ZN => n6618);
   U1012 : AOI21_X1 port map( B1 => n12541, B2 => DATA1(30), A => n11916, ZN =>
                           n11920);
   U1013 : NAND2_X1 port map( A1 => DATA1(26), A2 => n11917, ZN => n11919);
   U1014 : NAND2_X1 port map( A1 => DATA1(29), A2 => n12332, ZN => n12217);
   U1015 : NAND4_X1 port map( A1 => n11920, A2 => n11919, A3 => n12217, A4 => 
                           n11918, ZN => n6675);
   U1016 : AOI22_X1 port map( A1 => n13123, A2 => n11921, B1 => n13121, B2 => 
                           n13117, ZN => n11925);
   U1017 : AOI22_X1 port map( A1 => n1872, A2 => n11923, B1 => n13222, B2 => 
                           n11922, ZN => n11924);
   U1018 : OAI211_X1 port map( C1 => n13130, C2 => n13135, A => n11925, B => 
                           n11924, ZN => n1851);
   U1019 : INV_X1 port map( A => n1855, ZN => n11926);
   U1020 : AOI22_X1 port map( A1 => n11927, A2 => n1851, B1 => n1868, B2 => 
                           n11926, ZN => n6617);
   U1021 : AOI222_X1 port map( A1 => n11928, A2 => n11781, B1 => n11931, B2 => 
                           n13223, C1 => n11930, C2 => n1865, ZN => n13106);
   U1022 : INV_X1 port map( A => n11929, ZN => n11932);
   U1023 : AOI222_X1 port map( A1 => n13223, A2 => n11932, B1 => n1865, B2 => 
                           n11931, C1 => n11781, C2 => n11930, ZN => n13113);
   U1024 : OAI22_X1 port map( A1 => n13133, A2 => n13113, B1 => n13135, B2 => 
                           n13112, ZN => n11933);
   U1025 : INV_X1 port map( A => n11933, ZN => n11935);
   U1026 : INV_X1 port map( A => n11949, ZN => n11942);
   U1027 : AOI22_X1 port map( A1 => n13222, A2 => n13117, B1 => n13121, B2 => 
                           n11942, ZN => n11934);
   U1028 : OAI211_X1 port map( C1 => n13106, C2 => n11315, A => n11935, B => 
                           n11934, ZN => n7097);
   U1029 : OAI22_X1 port map( A1 => n13106, A2 => n13133, B1 => n13113, B2 => 
                           n13100, ZN => n11937);
   U1030 : OAI22_X1 port map( A1 => n13108, A2 => n13112, B1 => n1869, B2 => 
                           n11947, ZN => n11936);
   U1031 : AOI211_X1 port map( C1 => n13123, C2 => n11942, A => n11937, B => 
                           n11936, ZN => n7114);
   U1032 : NAND2_X1 port map( A1 => n12541, A2 => DATA1(31), ZN => n6742);
   U1033 : INV_X1 port map( A => DATA1(29), ZN => n12202);
   U1034 : NOR2_X1 port map( A1 => n12202, A2 => n12545, ZN => n12235);
   U1035 : AOI211_X1 port map( C1 => n12215, C2 => DATA1(28), A => n11938, B =>
                           n12235, ZN => n11939);
   U1036 : NAND2_X1 port map( A1 => DATA1(30), A2 => n12332, ZN => n12203);
   U1037 : NAND3_X1 port map( A1 => n11939, A2 => n12203, A3 => n6742, ZN => 
                           n6676);
   U1038 : OAI22_X1 port map( A1 => n13108, A2 => n13113, B1 => n1869, B2 => 
                           n11948, ZN => n11941);
   U1039 : OAI22_X1 port map( A1 => n13106, A2 => n13100, B1 => n11947, B2 => 
                           n11315, ZN => n11940);
   U1040 : AOI211_X1 port map( C1 => n1872, C2 => n11942, A => n11941, B => 
                           n11940, ZN => n7134);
   U1041 : XOR2_X1 port map( A => n1837, B => n4293, Z => n6749);
   U1042 : OAI21_X1 port map( B1 => DATA1(27), B2 => DATA2_I_27_port, A => 
                           n11943, ZN => n1800);
   U1043 : AOI21_X1 port map( B1 => n1802, B2 => n6106, A => n1800, ZN => n6869
                           );
   U1044 : OAI21_X1 port map( B1 => DATA1(29), B2 => n4395, A => n11944, ZN => 
                           n6850);
   U1045 : OAI21_X1 port map( B1 => n11944, B2 => n11946, A => n6740, ZN => 
                           n6733);
   U1046 : AOI21_X1 port map( B1 => n1802, B2 => n11945, A => n1800, ZN => 
                           n6870);
   U1047 : XOR2_X1 port map( A => DATA2_I_28_port, B => DATA1(28), Z => n6860);
   U1048 : OAI21_X1 port map( B1 => n4421, B2 => n6870, A => n6860, ZN => n6858
                           );
   U1049 : NAND2_X1 port map( A1 => n12756, A2 => n11946, ZN => n6739);
   U1050 : OAI221_X1 port map( B1 => DATA1(31), B2 => n1835, C1 => n1837, C2 =>
                           n12530, A => n12466, ZN => n6744);
   U1051 : OAI22_X1 port map( A1 => n13108, A2 => n13106, B1 => n11947, B2 => 
                           n13133, ZN => n6763);
   U1052 : OAI22_X1 port map( A1 => n11949, A2 => n13100, B1 => n11948, B2 => 
                           n11315, ZN => n6762);
   U1053 : AOI21_X1 port map( B1 => n9176, B2 => n8890, A => n8621, ZN => 
                           n12076);
   U1054 : OAI22_X1 port map( A1 => n8889, A2 => n12076, B1 => n9199, B2 => 
                           n8960, ZN => n11950);
   U1055 : AOI211_X1 port map( C1 => n8538, C2 => n8852, A => n9200, B => 
                           n11950, ZN => n11998);
   U1056 : AOI21_X1 port map( B1 => n8538, B2 => n9016, A => n8954, ZN => 
                           n11957);
   U1057 : OAI22_X1 port map( A1 => n13142, A2 => n11957, B1 => n13140, B2 => 
                           n11338, ZN => n11951);
   U1058 : INV_X1 port map( A => n11951, ZN => n11953);
   U1059 : OAI211_X1 port map( C1 => n8676, C2 => n9177, A => n8629, B => n8622
                           , ZN => n11994);
   U1060 : OAI211_X1 port map( C1 => n8676, C2 => n9178, A => n8628, B => n8623
                           , ZN => n11966);
   U1061 : AOI22_X1 port map( A1 => n8806, A2 => n11994, B1 => n9216, B2 => 
                           n11966, ZN => n11952);
   U1062 : OAI211_X1 port map( C1 => n11998, C2 => n9018, A => n11953, B => 
                           n11952, ZN => n12007);
   U1063 : OAI22_X1 port map( A1 => n13179, A2 => n11338, B1 => n13140, B2 => 
                           n11339, ZN => n11954);
   U1064 : INV_X1 port map( A => n11954, ZN => n11956);
   U1065 : AOI22_X1 port map( A1 => n8809, A2 => n11994, B1 => n8806, B2 => 
                           n11966, ZN => n11955);
   U1066 : OAI211_X1 port map( C1 => n11957, C2 => n9018, A => n11956, B => 
                           n11955, ZN => n11969);
   U1067 : INV_X1 port map( A => n11957, ZN => n11999);
   U1068 : AOI22_X1 port map( A1 => n8806, A2 => n11999, B1 => n9216, B2 => 
                           n11994, ZN => n11960);
   U1069 : INV_X1 port map( A => n12076, ZN => n12001);
   U1070 : AOI22_X1 port map( A1 => n9186, A2 => n12001, B1 => n9014, B2 => 
                           n13176, ZN => n11958);
   U1071 : OAI211_X1 port map( C1 => n8676, C2 => n9199, A => n8620, B => 
                           n11958, ZN => n12083);
   U1072 : AOI22_X1 port map( A1 => n8906, A2 => n12083, B1 => n9215, B2 => 
                           n11966, ZN => n11959);
   U1073 : OAI211_X1 port map( C1 => n9104, C2 => n11998, A => n11960, B => 
                           n11959, ZN => n12008);
   U1074 : AOI222_X1 port map( A1 => n12007, A2 => n8907, B1 => n11969, B2 => 
                           n9098, C1 => n12008, C2 => n9218, ZN => n12012);
   U1075 : INV_X1 port map( A => n12012, ZN => n12074);
   U1076 : OAI22_X1 port map( A1 => n9022, A2 => n11338, B1 => n8972, B2 => 
                           n11339, ZN => n11963);
   U1077 : AOI211_X1 port map( C1 => n8850, C2 => n8852, A => n8619, B => n8618
                           , ZN => n11979);
   U1078 : INV_X1 port map( A => n11994, ZN => n11961);
   U1079 : OAI22_X1 port map( A1 => n8895, A2 => n11979, B1 => n11961, B2 => 
                           n13164, ZN => n11962);
   U1080 : AOI211_X1 port map( C1 => n13144, C2 => n11966, A => n11963, B => 
                           n11962, ZN => n11975);
   U1081 : INV_X1 port map( A => n11975, ZN => n11968);
   U1082 : AOI222_X1 port map( A1 => n8907, A2 => n11969, B1 => n12007, B2 => 
                           n13147, C1 => n13156, C2 => n11968, ZN => n12073);
   U1083 : OAI22_X1 port map( A1 => n9181, A2 => n11338, B1 => n11339, B2 => 
                           n13139, ZN => n11965);
   U1084 : AOI211_X1 port map( C1 => n8850, C2 => n9016, A => n8617, B => n8616
                           , ZN => n11982);
   U1085 : OAI22_X1 port map( A1 => n9019, A2 => n11982, B1 => n9021, B2 => 
                           n11979, ZN => n11964);
   U1086 : AOI211_X1 port map( C1 => n13141, C2 => n11966, A => n11965, B => 
                           n11964, ZN => n11976);
   U1087 : INV_X1 port map( A => n11976, ZN => n11967);
   U1088 : AOI222_X1 port map( A1 => n11969, A2 => n13147, B1 => n13171, B2 => 
                           n11968, C1 => n11967, C2 => n13156, ZN => n12011);
   U1089 : OAI22_X1 port map( A1 => n9106, A2 => n12073, B1 => n8561, B2 => 
                           n12011, ZN => n11978);
   U1090 : OAI22_X1 port map( A1 => n9104, A2 => n11339, B1 => n9018, B2 => 
                           n11338, ZN => n11971);
   U1091 : OAI22_X1 port map( A1 => n9022, A2 => n11979, B1 => n9021, B2 => 
                           n11982, ZN => n11970);
   U1092 : AOI211_X1 port map( C1 => n9215, C2 => n8613, A => n11971, B => 
                           n11970, ZN => n11986);
   U1093 : INV_X1 port map( A => n11982, ZN => n11974);
   U1094 : OAI22_X1 port map( A1 => n8895, A2 => n8612, B1 => n13145, B2 => 
                           n13186, ZN => n11973);
   U1095 : OAI22_X1 port map( A1 => n9104, A2 => n11979, B1 => n9018, B2 => 
                           n11339, ZN => n11972);
   U1096 : AOI211_X1 port map( C1 => n13153, C2 => n11974, A => n11973, B => 
                           n11972, ZN => n11987);
   U1097 : OAI222_X1 port map( A1 => n9029, A2 => n11986, B1 => n11976, B2 => 
                           n9030, C1 => n8974, C2 => n11987, ZN => n12025);
   U1098 : INV_X1 port map( A => n12025, ZN => n12035);
   U1099 : OAI222_X1 port map( A1 => n9029, A2 => n11976, B1 => n9030, B2 => 
                           n11975, C1 => n8974, C2 => n11986, ZN => n12015);
   U1100 : INV_X1 port map( A => n12015, ZN => n12022);
   U1101 : OAI22_X1 port map( A1 => n13168, A2 => n12035, B1 => n9107, B2 => 
                           n12022, ZN => n11977);
   U1102 : AOI211_X1 port map( C1 => n13184, C2 => n12074, A => n11978, B => 
                           n11977, ZN => n12098);
   U1103 : INV_X1 port map( A => n12098, ZN => n12027);
   U1104 : OAI22_X1 port map( A1 => n13139, A2 => n13186, B1 => n9020, B2 => 
                           n8612, ZN => n11981);
   U1105 : OAI22_X1 port map( A1 => n9182, A2 => n11979, B1 => n9181, B2 => 
                           n11982, ZN => n11980);
   U1106 : AOI211_X1 port map( C1 => n13151, C2 => n13194, A => n11981, B => 
                           n11980, ZN => n12021);
   U1107 : INV_X1 port map( A => n12021, ZN => n11989);
   U1108 : OAI22_X1 port map( A1 => n9165, A2 => n8612, B1 => n9021, B2 => 
                           n8610, ZN => n11984);
   U1109 : OAI22_X1 port map( A1 => n9181, A2 => n9198, B1 => n11982, B2 => 
                           n9023, ZN => n11983);
   U1110 : AOI211_X1 port map( C1 => n9215, C2 => n8609, A => n11984, B => 
                           n11983, ZN => n12033);
   U1111 : OAI22_X1 port map( A1 => n9030, A2 => n11987, B1 => n8974, B2 => 
                           n12033, ZN => n11985);
   U1112 : AOI21_X1 port map( B1 => n13171, B2 => n11989, A => n11985, ZN => 
                           n12053);
   U1113 : OAI22_X1 port map( A1 => n9106, A2 => n12022, B1 => n12053, B2 => 
                           n13168, ZN => n11991);
   U1114 : OAI22_X1 port map( A1 => n9029, A2 => n11987, B1 => n9030, B2 => 
                           n11986, ZN => n11988);
   U1115 : AOI21_X1 port map( B1 => n13156, B2 => n11989, A => n11988, ZN => 
                           n12054);
   U1116 : OAI22_X1 port map( A1 => n8897, A2 => n12011, B1 => n9032, B2 => 
                           n12054, ZN => n11990);
   U1117 : AOI211_X1 port map( C1 => n13155, C2 => n12025, A => n11991, B => 
                           n11990, ZN => n12038);
   U1118 : OAI22_X1 port map( A1 => n8897, A2 => n12073, B1 => n12054, B2 => 
                           n13168, ZN => n11993);
   U1119 : OAI22_X1 port map( A1 => n8561, A2 => n12022, B1 => n9031, B2 => 
                           n12011, ZN => n11992);
   U1120 : AOI211_X1 port map( C1 => n13193, C2 => n12025, A => n11993, B => 
                           n11992, ZN => n12099);
   U1121 : OAI22_X1 port map( A1 => n9101, A2 => n12038, B1 => n9167, B2 => 
                           n12099, ZN => n12017);
   U1122 : OAI22_X1 port map( A1 => n9107, A2 => n12073, B1 => n9217, B2 => 
                           n12011, ZN => n12010);
   U1123 : AOI22_X1 port map( A1 => n9017, A2 => n11994, B1 => n9216, B2 => 
                           n11999, ZN => n11997);
   U1124 : AOI222_X1 port map( A1 => n8891, A2 => n8560, B1 => n9013, B2 => 
                           n8627, C1 => n8615, C2 => n9015, ZN => n12000);
   U1125 : AOI22_X1 port map( A1 => n9187, A2 => n13176, B1 => n9185, B2 => 
                           n12001, ZN => n11995);
   U1126 : OAI211_X1 port map( C1 => n8889, C2 => n12000, A => n8614, B => 
                           n11995, ZN => n12084);
   U1127 : AOI22_X1 port map( A1 => n8809, A2 => n12083, B1 => n13141, B2 => 
                           n12084, ZN => n11996);
   U1128 : OAI211_X1 port map( C1 => n11998, C2 => n13139, A => n11997, B => 
                           n11996, ZN => n12091);
   U1129 : INV_X1 port map( A => n12083, ZN => n12006);
   U1130 : INV_X1 port map( A => n11998, ZN => n12082);
   U1131 : AOI22_X1 port map( A1 => n9216, A2 => n12082, B1 => n9215, B2 => 
                           n11999, ZN => n12005);
   U1132 : AOI222_X1 port map( A1 => n8891, A2 => n8627, B1 => n9013, B2 => 
                           n8615, C1 => n9015, C2 => n8611, ZN => n12077);
   U1133 : AOI22_X1 port map( A1 => n9185, A2 => n13176, B1 => n8854, B2 => 
                           n8537, ZN => n12003);
   U1134 : INV_X1 port map( A => n12000, ZN => n12081);
   U1135 : AOI22_X1 port map( A1 => n9187, A2 => n12081, B1 => n8852, B2 => 
                           n12001, ZN => n12002);
   U1136 : OAI211_X1 port map( C1 => n8889, C2 => n12077, A => n12003, B => 
                           n12002, ZN => n12085);
   U1137 : AOI22_X1 port map( A1 => n8809, A2 => n12084, B1 => n8906, B2 => 
                           n12085, ZN => n12004);
   U1138 : OAI211_X1 port map( C1 => n9022, C2 => n12006, A => n12005, B => 
                           n12004, ZN => n12089);
   U1139 : AOI222_X1 port map( A1 => n12091, A2 => n8907, B1 => n12008, B2 => 
                           n9098, C1 => n12089, C2 => n9218, ZN => n12093);
   U1140 : AOI222_X1 port map( A1 => n12008, A2 => n8907, B1 => n12007, B2 => 
                           n9098, C1 => n12091, C2 => n9218, ZN => n12097);
   U1141 : OAI22_X1 port map( A1 => n8897, A2 => n12093, B1 => n9031, B2 => 
                           n12097, ZN => n12009);
   U1142 : AOI211_X1 port map( C1 => n9025, C2 => n12074, A => n12010, B => 
                           n12009, ZN => n12100);
   U1143 : OAI22_X1 port map( A1 => n8561, A2 => n12073, B1 => n9032, B2 => 
                           n12011, ZN => n12014);
   U1144 : OAI22_X1 port map( A1 => n8897, A2 => n12097, B1 => n12012, B2 => 
                           n13148, ZN => n12013);
   U1145 : AOI211_X1 port map( C1 => n13169, C2 => n12015, A => n12014, B => 
                           n12013, ZN => n12101);
   U1146 : OAI22_X1 port map( A1 => n8801, A2 => n12100, B1 => n12101, B2 => 
                           n9036, ZN => n12016);
   U1147 : AOI211_X1 port map( C1 => n13202, C2 => n12027, A => n12017, B => 
                           n12016, ZN => n12018);
   U1148 : INV_X1 port map( A => n12018, ZN => n12106);
   U1149 : AOI22_X1 port map( A1 => n9017, A2 => n8608, B1 => n8906, B2 => 
                           n8613, ZN => n12019);
   U1150 : OAI211_X1 port map( C1 => n9104, C2 => n8612, A => n8607, B => 
                           n12019, ZN => n12020);
   U1151 : INV_X1 port map( A => n12020, ZN => n12044);
   U1152 : OAI222_X1 port map( A1 => n8974, A2 => n12044, B1 => n12033, B2 => 
                           n9029, C1 => n12021, C2 => n9030, ZN => n12059);
   U1153 : INV_X1 port map( A => n12059, ZN => n12034);
   U1154 : OAI22_X1 port map( A1 => n8897, A2 => n12022, B1 => n12034, B2 => 
                           n13168, ZN => n12024);
   U1155 : OAI22_X1 port map( A1 => n8561, A2 => n12054, B1 => n9032, B2 => 
                           n12053, ZN => n12023);
   U1156 : AOI211_X1 port map( C1 => n13167, C2 => n12025, A => n12024, B => 
                           n12023, ZN => n12026);
   U1157 : INV_X1 port map( A => n12026, ZN => n12070);
   U1158 : INV_X1 port map( A => n12038, ZN => n12069);
   U1159 : AOI22_X1 port map( A1 => n13212, A2 => n12070, B1 => n12069, B2 => 
                           n8804, ZN => n12030);
   U1160 : INV_X1 port map( A => n12101, ZN => n12028);
   U1161 : AOI22_X1 port map( A1 => n13166, A2 => n12028, B1 => n13157, B2 => 
                           n12027, ZN => n12029);
   U1162 : OAI211_X1 port map( C1 => n8678, C2 => n12099, A => n12030, B => 
                           n12029, ZN => n12109);
   U1163 : INV_X1 port map( A => n12053, ZN => n12060);
   U1164 : OAI22_X1 port map( A1 => n13142, A2 => n13201, B1 => n8972, B2 => 
                           n9196, ZN => n12032);
   U1165 : OAI22_X1 port map( A1 => n9022, A2 => n9194, B1 => n9182, B2 => 
                           n8612, ZN => n12031);
   U1166 : AOI211_X1 port map( C1 => n13195, C2 => n13152, A => n12032, B => 
                           n12031, ZN => n12049);
   U1167 : OAI222_X1 port map( A1 => n8974, A2 => n12049, B1 => n12044, B2 => 
                           n9029, C1 => n12033, C2 => n9030, ZN => n12058);
   U1168 : INV_X1 port map( A => n12058, ZN => n12136);
   U1169 : OAI22_X1 port map( A1 => n9217, A2 => n12136, B1 => n12034, B2 => 
                           n13150, ZN => n12037);
   U1170 : OAI22_X1 port map( A1 => n12035, A2 => n13189, B1 => n12054, B2 => 
                           n13148, ZN => n12036);
   U1171 : AOI211_X1 port map( C1 => n9025, C2 => n12060, A => n12037, B => 
                           n12036, ZN => n12140);
   U1172 : OAI22_X1 port map( A1 => n8677, A2 => n12038, B1 => n12140, B2 => 
                           n13165, ZN => n12040);
   U1173 : OAI22_X1 port map( A1 => n8801, A2 => n12098, B1 => n12099, B2 => 
                           n9036, ZN => n12039);
   U1174 : AOI211_X1 port map( C1 => n13172, C2 => n12070, A => n12040, B => 
                           n12039, ZN => n12041);
   U1175 : INV_X1 port map( A => n12041, ZN => n12108);
   U1176 : AOI222_X1 port map( A1 => n8909, A2 => n12106, B1 => n9035, B2 => 
                           n12109, C1 => n9034, C2 => n12108, ZN => n12149);
   U1177 : INV_X1 port map( A => n12149, ZN => n12114);
   U1178 : OAI22_X1 port map( A1 => n8610, A2 => n9023, B1 => n13140, B2 => 
                           n13154, ZN => n12043);
   U1179 : OAI22_X1 port map( A1 => n9022, A2 => n9196, B1 => n9181, B2 => 
                           n9194, ZN => n12042);
   U1180 : AOI211_X1 port map( C1 => n13146, C2 => n13152, A => n12043, B => 
                           n12042, ZN => n12050);
   U1181 : OAI222_X1 port map( A1 => n9029, A2 => n12049, B1 => n9030, B2 => 
                           n12044, C1 => n8974, C2 => n12050, ZN => n12374);
   U1182 : OAI22_X1 port map( A1 => n9104, A2 => n9196, B1 => n13179, B2 => 
                           n13154, ZN => n12046);
   U1183 : OAI22_X1 port map( A1 => n9019, A2 => n8849, B1 => n9023, B2 => 
                           n9194, ZN => n12045);
   U1184 : AOI211_X1 port map( C1 => n13170, C2 => n13152, A => n12046, B => 
                           n12045, ZN => n12132);
   U1185 : OAI22_X1 port map( A1 => n9023, A2 => n9196, B1 => n13139, B2 => 
                           n13154, ZN => n12048);
   U1186 : OAI22_X1 port map( A1 => n9181, A2 => n9195, B1 => n9019, B2 => 
                           n8604, ZN => n12047);
   U1187 : AOI211_X1 port map( C1 => n13146, C2 => n13197, A => n12048, B => 
                           n12047, ZN => n12443);
   U1188 : OAI222_X1 port map( A1 => n9029, A2 => n12132, B1 => n9030, B2 => 
                           n12050, C1 => n8974, C2 => n12443, ZN => n12410);
   U1189 : AOI22_X1 port map( A1 => n9025, A2 => n12374, B1 => n9026, B2 => 
                           n12410, ZN => n12052);
   U1190 : OAI222_X1 port map( A1 => n9029, A2 => n12050, B1 => n9030, B2 => 
                           n12049, C1 => n8974, C2 => n12132, ZN => n12389);
   U1191 : AOI22_X1 port map( A1 => n8807, A2 => n12389, B1 => n9183, B2 => 
                           n12059, ZN => n12051);
   U1192 : OAI211_X1 port map( C1 => n9106, C2 => n12136, A => n12052, B => 
                           n12051, ZN => n12288);
   U1193 : AOI22_X1 port map( A1 => n9025, A2 => n12059, B1 => n9026, B2 => 
                           n12374, ZN => n12057);
   U1194 : OAI22_X1 port map( A1 => n13143, A2 => n12054, B1 => n9106, B2 => 
                           n12053, ZN => n12055);
   U1195 : INV_X1 port map( A => n12055, ZN => n12056);
   U1196 : OAI211_X1 port map( C1 => n12136, C2 => n13150, A => n12057, B => 
                           n12056, ZN => n12067);
   U1197 : AOI22_X1 port map( A1 => n8973, A2 => n12288, B1 => n13202, B2 => 
                           n12067, ZN => n12064);
   U1198 : INV_X1 port map( A => n12374, ZN => n12135);
   U1199 : AOI22_X1 port map( A1 => n9025, A2 => n12058, B1 => n9026, B2 => 
                           n12389, ZN => n12062);
   U1200 : AOI22_X1 port map( A1 => n9183, A2 => n12060, B1 => n13167, B2 => 
                           n12059, ZN => n12061);
   U1201 : OAI211_X1 port map( C1 => n12135, C2 => n13150, A => n12062, B => 
                           n12061, ZN => n12139);
   U1202 : AOI22_X1 port map( A1 => n8804, A2 => n12139, B1 => n9010, B2 => 
                           n12070, ZN => n12063);
   U1203 : OAI211_X1 port map( C1 => n12140, C2 => n13181, A => n12064, B => 
                           n12063, ZN => n12144);
   U1204 : INV_X1 port map( A => n12140, ZN => n12068);
   U1205 : AOI22_X1 port map( A1 => n8804, A2 => n12068, B1 => n8973, B2 => 
                           n12067, ZN => n12066);
   U1206 : AOI22_X1 port map( A1 => n13202, A2 => n12070, B1 => n13157, B2 => 
                           n12069, ZN => n12065);
   U1207 : OAI211_X1 port map( C1 => n8801, C2 => n12099, A => n12066, B => 
                           n12065, ZN => n12110);
   U1208 : INV_X1 port map( A => n12067, ZN => n12287);
   U1209 : AOI22_X1 port map( A1 => n8973, A2 => n12139, B1 => n9173, B2 => 
                           n12068, ZN => n12072);
   U1210 : AOI22_X1 port map( A1 => n8899, A2 => n12070, B1 => n9164, B2 => 
                           n12069, ZN => n12071);
   U1211 : OAI211_X1 port map( C1 => n9167, C2 => n12287, A => n12072, B => 
                           n12071, ZN => n12143);
   U1212 : AOI222_X1 port map( A1 => n12144, A2 => n9034, B1 => n12110, B2 => 
                           n8909, C1 => n12143, C2 => n9035, ZN => n12127);
   U1213 : AOI222_X1 port map( A1 => n12143, A2 => n9034, B1 => n12108, B2 => 
                           n8909, C1 => n12110, C2 => n9035, ZN => n12128);
   U1214 : OAI22_X1 port map( A1 => n12127, A2 => n8970, B1 => n12128, B2 => 
                           n9169, ZN => n12113);
   U1215 : INV_X1 port map( A => n12073, ZN => n12075);
   U1216 : AOI22_X1 port map( A1 => n13169, A2 => n12075, B1 => n12074, B2 => 
                           n8807, ZN => n12096);
   U1217 : OAI22_X1 port map( A1 => n9180, A2 => n11304, B1 => n9028, B2 => 
                           n12076, ZN => n12080);
   U1218 : AOI222_X1 port map( A1 => n8891, A2 => n8615, B1 => n9013, B2 => 
                           n8611, C1 => n9015, C2 => n8605, ZN => n12078);
   U1219 : OAI22_X1 port map( A1 => n8889, A2 => n12078, B1 => n8960, B2 => 
                           n12077, ZN => n12079);
   U1220 : AOI211_X1 port map( C1 => n9185, C2 => n12081, A => n12080, B => 
                           n12079, ZN => n12088);
   U1221 : AOI22_X1 port map( A1 => n9216, A2 => n12083, B1 => n9215, B2 => 
                           n12082, ZN => n12087);
   U1222 : AOI22_X1 port map( A1 => n8809, A2 => n12085, B1 => n8806, B2 => 
                           n12084, ZN => n12086);
   U1223 : OAI211_X1 port map( C1 => n9182, C2 => n12088, A => n12087, B => 
                           n12086, ZN => n12090);
   U1224 : AOI222_X1 port map( A1 => n12091, A2 => n9008, B1 => n12090, B2 => 
                           n9011, C1 => n12089, C2 => n8907, ZN => n12092);
   U1225 : OAI22_X1 port map( A1 => n9106, A2 => n12093, B1 => n8897, B2 => 
                           n12092, ZN => n12094);
   U1226 : INV_X1 port map( A => n12094, ZN => n12095);
   U1227 : OAI211_X1 port map( C1 => n8561, C2 => n12097, A => n12096, B => 
                           n12095, ZN => n12104);
   U1228 : OAI22_X1 port map( A1 => n9101, A2 => n12099, B1 => n9167, B2 => 
                           n12098, ZN => n12103);
   U1229 : OAI22_X1 port map( A1 => n8678, A2 => n12101, B1 => n9166, B2 => 
                           n12100, ZN => n12102);
   U1230 : AOI211_X1 port map( C1 => n13166, C2 => n12104, A => n12103, B => 
                           n12102, ZN => n12105);
   U1231 : INV_X1 port map( A => n12105, ZN => n12107);
   U1232 : AOI222_X1 port map( A1 => n12109, A2 => n9175, B1 => n12107, B2 => 
                           n8910, C1 => n12106, C2 => n9111, ZN => n12111);
   U1233 : AOI222_X1 port map( A1 => n12110, A2 => n9034, B1 => n12109, B2 => 
                           n8909, C1 => n12108, C2 => n9035, ZN => n12146);
   U1234 : OAI22_X1 port map( A1 => n8802, A2 => n12111, B1 => n9037, B2 => 
                           n12146, ZN => n12112);
   U1235 : AOI211_X1 port map( C1 => n9112, C2 => n12114, A => n12113, B => 
                           n12112, ZN => n12152);
   U1236 : OAI21_X1 port map( B1 => n8848, B2 => n8901, A => n8951, ZN => 
                           n12224);
   U1237 : AOI21_X1 port map( B1 => n8955, B2 => n12224, A => n8847, ZN => 
                           n12157);
   U1238 : AOI21_X1 port map( B1 => n8955, B2 => n8844, A => n8847, ZN => 
                           n12156);
   U1239 : OAI22_X1 port map( A1 => n9039, A2 => n12157, B1 => n8961, B2 => 
                           n12156, ZN => n12115);
   U1240 : INV_X1 port map( A => n12115, ZN => n12207);
   U1241 : OAI21_X1 port map( B1 => n12207, B2 => n9192, A => n8843, ZN => 
                           n12116);
   U1242 : INV_X1 port map( A => n12116, ZN => n12161);
   U1243 : NOR2_X1 port map( A1 => n12161, A2 => n8952, ZN => n12126);
   U1244 : AOI22_X1 port map( A1 => n9179, A2 => n8554, B1 => n8949, B2 => 
                           n9209, ZN => n12124);
   U1245 : INV_X1 port map( A => n12157, ZN => n12118);
   U1246 : INV_X1 port map( A => n12156, ZN => n12117);
   U1247 : OAI22_X1 port map( A1 => n9114, A2 => n12118, B1 => n8962, B2 => 
                           n12117, ZN => n12120);
   U1248 : NAND2_X1 port map( A1 => n9114, A2 => n8962, ZN => n12119);
   U1249 : AOI22_X1 port map( A1 => n9193, A2 => n12120, B1 => n8846, B2 => 
                           n12119, ZN => n12121);
   U1250 : INV_X1 port map( A => n12121, ZN => n12122);
   U1251 : AOI22_X1 port map( A1 => n8952, A2 => n12122, B1 => n9210, B2 => 
                           n8679, ZN => n12123);
   U1252 : OAI211_X1 port map( C1 => n9100, C2 => n8953, A => n12124, B => 
                           n12123, ZN => n12125);
   U1253 : AOI21_X1 port map( B1 => n12126, B2 => n8950, A => n12125, ZN => 
                           n12151);
   U1254 : INV_X1 port map( A => n12127, ZN => n12241);
   U1255 : INV_X1 port map( A => n12128, ZN => n12223);
   U1256 : AOI22_X1 port map( A1 => n8808, A2 => n12241, B1 => n8904, B2 => 
                           n12223, ZN => n12148);
   U1257 : AOI211_X1 port map( C1 => n8540, C2 => n8853, A => n8603, B => n8602
                           , ZN => n12526);
   U1258 : AOI22_X1 port map( A1 => n8809, A2 => n8606, B1 => n13141, B2 => 
                           n13152, ZN => n12131);
   U1259 : OAI22_X1 port map( A1 => n9022, A2 => n8849, B1 => n8972, B2 => 
                           n8604, ZN => n12129);
   U1260 : INV_X1 port map( A => n12129, ZN => n12130);
   U1261 : OAI211_X1 port map( C1 => n9019, C2 => n12526, A => n12131, B => 
                           n12130, ZN => n12460);
   U1262 : INV_X1 port map( A => n12460, ZN => n12133);
   U1263 : OAI222_X1 port map( A1 => n8974, A2 => n12133, B1 => n12443, B2 => 
                           n9029, C1 => n12132, C2 => n9030, ZN => n12420);
   U1264 : AOI22_X1 port map( A1 => n13155, A2 => n12389, B1 => n12420, B2 => 
                           n9026, ZN => n12134);
   U1265 : INV_X1 port map( A => n12134, ZN => n12138);
   U1266 : OAI22_X1 port map( A1 => n8897, A2 => n12136, B1 => n12135, B2 => 
                           n13148, ZN => n12137);
   U1267 : AOI211_X1 port map( C1 => n8807, C2 => n12410, A => n12138, B => 
                           n12137, ZN => n12323);
   U1268 : OAI22_X1 port map( A1 => n9101, A2 => n12323, B1 => n12287, B2 => 
                           n13181, ZN => n12142);
   U1269 : INV_X1 port map( A => n12139, ZN => n12303);
   U1270 : OAI22_X1 port map( A1 => n8677, A2 => n12303, B1 => n8801, B2 => 
                           n12140, ZN => n12141);
   U1271 : AOI211_X1 port map( C1 => n13172, C2 => n12288, A => n12142, B => 
                           n12141, ZN => n12271);
   U1272 : INV_X1 port map( A => n12143, ZN => n12145);
   U1273 : INV_X1 port map( A => n12144, ZN => n12261);
   U1274 : OAI222_X1 port map( A1 => n9219, A2 => n12271, B1 => n9163, B2 => 
                           n12145, C1 => n8908, C2 => n12261, ZN => n12252);
   U1275 : INV_X1 port map( A => n12146, ZN => n12208);
   U1276 : AOI22_X1 port map( A1 => n9099, A2 => n12252, B1 => n9112, B2 => 
                           n12208, ZN => n12147);
   U1277 : OAI211_X1 port map( C1 => n8802, C2 => n12149, A => n12148, B => 
                           n12147, ZN => n12159);
   U1278 : NAND3_X1 port map( A1 => n9212, A2 => n8626, A3 => n12159, ZN => 
                           n12150);
   U1279 : OAI211_X1 port map( C1 => n9109, C2 => n12152, A => n12151, B => 
                           n12150, ZN => OUTALU(31));
   U1280 : INV_X1 port map( A => DATA2(30), ZN => n12758);
   U1281 : AOI22_X1 port map( A1 => DATA1(30), A2 => n12758, B1 => DATA2(30), 
                           B2 => n12586, ZN => n12712);
   U1282 : INV_X1 port map( A => n1833, ZN => n12220);
   U1283 : OAI22_X1 port map( A1 => n12586, A2 => n12341, B1 => n12163, B2 => 
                           n1837, ZN => n12153);
   U1284 : AOI22_X1 port map( A1 => n13224, A2 => n8681, B1 => n12220, B2 => 
                           n12153, ZN => n12155);
   U1285 : OAI211_X1 port map( C1 => n12518, C2 => n12519, A => DATA1(30), B =>
                           DATA2(30), ZN => n12154);
   U1286 : OAI211_X1 port map( C1 => n12712, C2 => n1835, A => n12155, B => 
                           n12154, ZN => n6793);
   U1287 : AOI22_X1 port map( A1 => n12157, A2 => n8903, B1 => n12156, B2 => 
                           n9115, ZN => n12162);
   U1288 : NOR2_X1 port map( A1 => n8843, A2 => n13211, ZN => n12158);
   U1289 : AOI211_X1 port map( C1 => n8969, C2 => n12159, A => n8601, B => 
                           n12158, ZN => n12160);
   U1290 : OAI221_X1 port map( B1 => n9193, B2 => n12162, C1 => n13209, C2 => 
                           n12161, A => n12160, ZN => OUTALU(30));
   U1291 : NOR2_X1 port map( A1 => n9205, A2 => n12341, ZN => n12164);
   U1292 : NOR2_X1 port map( A1 => n12163, A2 => n11332, ZN => n12542);
   U1293 : AOI211_X1 port map( C1 => n12216, C2 => n9221, A => n12164, B => 
                           n12542, ZN => n3875);
   U1294 : AOI211_X1 port map( C1 => n12167, C2 => n12171, A => n12166, B => 
                           n12165, ZN => n12176);
   U1295 : AOI22_X1 port map( A1 => DATA2(2), A2 => n9223, B1 => n9205, B2 => 
                           n13077, ZN => n12590);
   U1296 : INV_X1 port map( A => n12590, ZN => n12640);
   U1297 : OAI211_X1 port map( C1 => n12518, C2 => n13177, A => DATA2(2), B => 
                           n12477, ZN => n12174);
   U1298 : NOR2_X1 port map( A1 => n12168, A2 => n12328, ZN => n12170);
   U1299 : AOI211_X1 port map( C1 => n12171, C2 => n12170, A => n12327, B => 
                           n12169, ZN => n12172);
   U1300 : INV_X1 port map( A => n12172, ZN => n12173);
   U1301 : OAI211_X1 port map( C1 => n12640, C2 => n1835, A => n12174, B => 
                           n12173, ZN => n12175);
   U1302 : AOI211_X1 port map( C1 => n8861, C2 => n13224, A => n12176, B => 
                           n12175, ZN => n6837);
   U1303 : AOI211_X1 port map( C1 => n12179, C2 => DATA1(5), A => n12178, B => 
                           n12177, ZN => n12181);
   U1304 : NAND2_X1 port map( A1 => DATA1(4), A2 => n12216, ZN => n12180);
   U1305 : OAI211_X1 port map( C1 => n9205, C2 => n12341, A => n12181, B => 
                           n12180, ZN => n12548);
   U1306 : AOI222_X1 port map( A1 => n12183, A2 => n11781, B1 => n12548, B2 => 
                           n12182, C1 => n12342, C2 => n1865, ZN => n12538);
   U1307 : OAI22_X1 port map( A1 => n13108, A2 => n12538, B1 => n13102, B2 => 
                           n13133, ZN => n12185);
   U1308 : OAI22_X1 port map( A1 => n1869, A2 => n13118, B1 => n13101, B2 => 
                           n11315, ZN => n12184);
   U1309 : AOI211_X1 port map( C1 => n13221, C2 => n12553, A => n12185, B => 
                           n12184, ZN => n7284);
   U1310 : OAI22_X1 port map( A1 => n12359, A2 => n9037, B1 => n12186, B2 => 
                           n9040, ZN => n12200);
   U1311 : INV_X1 port map( A => n12187, ZN => n12190);
   U1312 : OAI22_X1 port map( A1 => n9165, A2 => n9191, B1 => n8630, B2 => 
                           n13142, ZN => n12189);
   U1313 : OAI22_X1 port map( A1 => n9182, A2 => n8598, B1 => n8895, B2 => 
                           n8641, ZN => n12188);
   U1314 : AOI211_X1 port map( C1 => n13146, C2 => n13187, A => n12189, B => 
                           n12188, ZN => n12723);
   U1315 : OAI222_X1 port map( A1 => n8975, A2 => n12190, B1 => n9103, B2 => 
                           n12347, C1 => n8896, C2 => n12723, ZN => n12725);
   U1316 : AOI22_X1 port map( A1 => n9183, A2 => n12725, B1 => n12348, B2 => 
                           n13199, ZN => n12193);
   U1317 : AOI22_X1 port map( A1 => n12191, A2 => n13169, B1 => n12727, B2 => 
                           n13155, ZN => n12192);
   U1318 : OAI211_X1 port map( C1 => n12349, C2 => n9032, A => n12193, B => 
                           n12192, ZN => n12731);
   U1319 : AOI22_X1 port map( A1 => n9164, A2 => n12731, B1 => n12354, B2 => 
                           n13178, ZN => n12196);
   U1320 : AOI22_X1 port map( A1 => n8899, A2 => n12733, B1 => n8804, B2 => 
                           n12194, ZN => n12195);
   U1321 : OAI211_X1 port map( C1 => n12197, C2 => n13165, A => n12196, B => 
                           n12195, ZN => n12739);
   U1322 : AOI222_X1 port map( A1 => n12198, A2 => n9034, B1 => n12358, B2 => 
                           n9035, C1 => n12739, C2 => n8909, ZN => n12742);
   U1323 : OAI22_X1 port map( A1 => n8805, A2 => n12743, B1 => n12742, B2 => 
                           n8802, ZN => n12199);
   U1324 : OAI21_X1 port map( B1 => n12200, B2 => n12199, A => n8902, ZN => 
                           n12201);
   U1325 : OAI211_X1 port map( C1 => n9109, C2 => n8600, A => n8599, B => 
                           n12201, ZN => OUTALU(2));
   U1326 : INV_X1 port map( A => DATA2(29), ZN => n12759);
   U1327 : NAND2_X1 port map( A1 => DATA1(29), A2 => n12759, ZN => n12709);
   U1328 : NAND2_X1 port map( A1 => DATA2(29), A2 => n12202, ZN => n12711);
   U1329 : NAND2_X1 port map( A1 => n12709, A2 => n12711, ZN => n1838);
   U1330 : AOI22_X1 port map( A1 => n12535, A2 => n1838, B1 => n6095, B2 => 
                           n8682, ZN => n6853);
   U1331 : OAI21_X1 port map( B1 => n12530, B2 => n12202, A => n12466, ZN => 
                           n12206);
   U1332 : OAI211_X1 port map( C1 => n1837, C2 => n12545, A => n12204, B => 
                           n12203, ZN => n12205);
   U1333 : AOI22_X1 port map( A1 => DATA2(29), A2 => n12206, B1 => n12220, B2 
                           => n12205, ZN => n6852);
   U1334 : OAI22_X1 port map( A1 => n8961, A2 => n8844, B1 => n9039, B2 => 
                           n12224, ZN => n12213);
   U1335 : AOI21_X1 port map( B1 => n8955, B2 => n8847, A => n12207, ZN => 
                           n12212);
   U1336 : AOI22_X1 port map( A1 => n9112, A2 => n12223, B1 => n8904, B2 => 
                           n12241, ZN => n12210);
   U1337 : AOI22_X1 port map( A1 => n8808, A2 => n12252, B1 => n9168, B2 => 
                           n12208, ZN => n12209);
   U1338 : AOI21_X1 port map( B1 => n12210, B2 => n12209, A => n9109, ZN => 
                           n12211);
   U1339 : AOI211_X1 port map( C1 => n8847, C2 => n12213, A => n12212, B => 
                           n12211, ZN => n12214);
   U1340 : NAND3_X1 port map( A1 => n8596, A2 => n8595, A3 => n12214, ZN => 
                           OUTALU(29));
   U1341 : NAND3_X1 port map( A1 => n12477, A2 => DATA1(28), A3 => DATA2(28), 
                           ZN => n12222);
   U1342 : AOI22_X1 port map( A1 => DATA1(30), A2 => n12216, B1 => n12215, B2 
                           => DATA1(31), ZN => n12218);
   U1343 : OAI211_X1 port map( C1 => n12341, C2 => n12710, A => n12218, B => 
                           n12217, ZN => n12219);
   U1344 : INV_X1 port map( A => DATA2(28), ZN => n12760);
   U1345 : OAI22_X1 port map( A1 => n12760, A2 => n12710, B1 => DATA1(28), B2 
                           => DATA2(28), ZN => n12580);
   U1346 : INV_X1 port map( A => n12580, ZN => n12705);
   U1347 : AOI22_X1 port map( A1 => n12220, A2 => n12219, B1 => n12535, B2 => 
                           n12705, ZN => n12221);
   U1348 : NAND2_X1 port map( A1 => n12222, A2 => n12221, ZN => n6865);
   U1349 : NOR2_X1 port map( A1 => n4421, A2 => n6860, ZN => n6862);
   U1350 : AOI222_X1 port map( A1 => n12241, A2 => n9112, B1 => n12252, B2 => 
                           n8904, C1 => n12223, C2 => n9168, ZN => n12231);
   U1351 : AOI21_X1 port map( B1 => n8683, B2 => n9211, A => n8594, ZN => 
                           n12230);
   U1352 : OAI21_X1 port map( B1 => n13163, B2 => n8848, A => n12224, ZN => 
                           n12225);
   U1353 : INV_X1 port map( A => n12225, ZN => n12228);
   U1354 : AOI22_X1 port map( A1 => n13210, A2 => n8845, B1 => n13163, B2 => 
                           n8844, ZN => n12226);
   U1355 : INV_X1 port map( A => n12226, ZN => n12227);
   U1356 : AOI22_X1 port map( A1 => n8903, A2 => n12228, B1 => n9038, B2 => 
                           n12227, ZN => n12229);
   U1357 : OAI211_X1 port map( C1 => n9109, C2 => n12231, A => n12230, B => 
                           n12229, ZN => OUTALU(28));
   U1358 : INV_X1 port map( A => DATA2(27), ZN => n12761);
   U1359 : OAI21_X1 port map( B1 => n12530, B2 => n12761, A => n12466, ZN => 
                           n4078);
   U1360 : OAI22_X1 port map( A1 => n11895, A2 => n1837, B1 => n12586, B2 => 
                           n12232, ZN => n12233);
   U1361 : NOR4_X1 port map( A1 => n12236, A2 => n12235, A3 => n12234, A4 => 
                           n12233, ZN => n6881);
   U1362 : NOR3_X1 port map( A1 => n6881, A2 => n1833, A3 => n12237, ZN => 
                           n6874);
   U1363 : INV_X1 port map( A => n1803, ZN => n12238);
   U1364 : NOR2_X1 port map( A1 => n6870, A2 => n12238, ZN => n6876);
   U1365 : NOR2_X1 port map( A1 => DATA2(27), A2 => n12239, ZN => n12627);
   U1366 : NOR2_X1 port map( A1 => DATA1(27), A2 => n12761, ZN => n12706);
   U1367 : OR2_X1 port map( A1 => n12627, A2 => n12706, ZN => n12240);
   U1368 : AOI22_X1 port map( A1 => n12535, A2 => n12240, B1 => n6095, B2 => 
                           n8685, ZN => n6871);
   U1369 : AOI22_X1 port map( A1 => n9112, A2 => n12252, B1 => n9168, B2 => 
                           n12241, ZN => n12247);
   U1370 : AOI22_X1 port map( A1 => n8947, A2 => n9171, B1 => n8842, B2 => 
                           n9002, ZN => n12245);
   U1371 : NOR2_X1 port map( A1 => n8848, A2 => n9114, ZN => n12242);
   U1372 : AOI21_X1 port map( B1 => n9207, B2 => n12242, A => n8841, ZN => 
                           n12244);
   U1373 : OAI22_X1 port map( A1 => n12242, A2 => n8947, B1 => n8965, B2 => 
                           n8799, ZN => n12243);
   U1374 : AND4_X1 port map( A1 => n12245, A2 => n8840, A3 => n12244, A4 => 
                           n12243, ZN => n12246);
   U1375 : OAI21_X1 port map( B1 => n9033, B2 => n12247, A => n12246, ZN => 
                           OUTALU(27));
   U1376 : INV_X1 port map( A => DATA2(26), ZN => n12762);
   U1377 : AOI22_X1 port map( A1 => DATA1(26), A2 => n12762, B1 => DATA2(26), 
                           B2 => n12572, ZN => n12702);
   U1378 : NAND3_X1 port map( A1 => DATA2(26), A2 => DATA1(26), A3 => n12477, 
                           ZN => n12250);
   U1379 : NAND3_X1 port map( A1 => n12257, A2 => n12269, A3 => n12248, ZN => 
                           n12249);
   U1380 : OAI211_X1 port map( C1 => n12702, C2 => n1835, A => n12250, B => 
                           n12249, ZN => n6889);
   U1381 : OAI22_X1 port map( A1 => n8968, A2 => n8672, B1 => n8668, B2 => 
                           n8967, ZN => n12251);
   U1382 : NAND2_X1 port map( A1 => n13204, A2 => n12251, ZN => n12255);
   U1383 : AOI211_X1 port map( C1 => n8686, C2 => n9211, A => n8593, B => n8839
                           , ZN => n12254);
   U1384 : NAND3_X1 port map( A1 => n8969, A2 => n9168, A3 => n12252, ZN => 
                           n12253);
   U1385 : NAND3_X1 port map( A1 => n12255, A2 => n12254, A3 => n12253, ZN => 
                           OUTALU(26));
   U1386 : INV_X1 port map( A => DATA2(25), ZN => n12763);
   U1387 : NAND2_X1 port map( A1 => n12763, A2 => DATA1(25), ZN => n12633);
   U1388 : NAND2_X1 port map( A1 => DATA2(25), A2 => n12256, ZN => n12701);
   U1389 : NAND2_X1 port map( A1 => n12633, A2 => n12701, ZN => n12560);
   U1390 : AOI22_X1 port map( A1 => n12535, A2 => n12560, B1 => n6095, B2 => 
                           n8690, ZN => n3867);
   U1391 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n12477, 
                           ZN => n3866);
   U1392 : AOI211_X1 port map( C1 => n12268, C2 => n12259, A => n12257, B => 
                           n1804, ZN => n6896);
   U1393 : AOI21_X1 port map( B1 => n12259, B2 => n12265, A => n12258, ZN => 
                           n12260);
   U1394 : NAND2_X1 port map( A1 => n1803, A2 => n12260, ZN => n6899);
   U1395 : OAI22_X1 port map( A1 => n9163, A2 => n12261, B1 => n8908, B2 => 
                           n12271, ZN => n12262);
   U1396 : AOI211_X1 port map( C1 => n8969, C2 => n12262, A => n8591, B => 
                           n13215, ZN => n12264);
   U1397 : INV_X1 port map( A => n12302, ZN => n12289);
   U1398 : OR3_X1 port map( A1 => n8889, A2 => n12289, A3 => n9009, ZN => 
                           n12263);
   U1399 : NAND4_X1 port map( A1 => n8838, A2 => n8946, A3 => n12264, A4 => 
                           n12263, ZN => OUTALU(25));
   U1400 : INV_X1 port map( A => DATA2(24), ZN => n12764);
   U1401 : OAI22_X1 port map( A1 => n12700, A2 => DATA2(24), B1 => n12764, B2 
                           => DATA1(24), ZN => n12556);
   U1402 : AOI22_X1 port map( A1 => n8692, A2 => n13224, B1 => n12535, B2 => 
                           n12556, ZN => n3865);
   U1403 : INV_X1 port map( A => n12268, ZN => n12266);
   U1404 : NAND3_X1 port map( A1 => n1803, A2 => n12266, A3 => n12265, ZN => 
                           n4075);
   U1405 : AOI22_X1 port map( A1 => DATA2(24), A2 => n12519, B1 => n12269, B2 
                           => DATA2_I_24_port, ZN => n12267);
   U1406 : AOI21_X1 port map( B1 => n12267, B2 => n12466, A => n12700, ZN => 
                           n6905);
   U1407 : NAND2_X1 port map( A1 => n12269, A2 => n12268, ZN => n6908);
   U1408 : OAI22_X1 port map( A1 => n8889, A2 => n12300, B1 => n12289, B2 => 
                           n8960, ZN => n12270);
   U1409 : AOI211_X1 port map( C1 => n8902, C2 => n12270, A => n8836, B => 
                           n13216, ZN => n12273);
   U1410 : OR3_X1 port map( A1 => n9163, A2 => n12271, A3 => n9109, ZN => 
                           n12272);
   U1411 : NAND4_X1 port map( A1 => n8837, A2 => n8945, A3 => n12273, A4 => 
                           n12272, ZN => OUTALU(24));
   U1412 : INV_X1 port map( A => DATA2(23), ZN => n12765);
   U1413 : NAND2_X1 port map( A1 => DATA1(23), A2 => n12765, ZN => n12274);
   U1414 : NOR2_X1 port map( A1 => n12765, A2 => DATA1(23), ZN => n12569);
   U1415 : INV_X1 port map( A => n12569, ZN => n12695);
   U1416 : AOI21_X1 port map( B1 => n12274, B2 => n12695, A => n1835, ZN => 
                           n4074);
   U1417 : AOI21_X1 port map( B1 => DATA2(23), B2 => n12519, A => n12518, ZN =>
                           n4073);
   U1418 : INV_X1 port map( A => n12283, ZN => n12286);
   U1419 : INV_X1 port map( A => n12282, ZN => n12278);
   U1420 : INV_X1 port map( A => n12279, ZN => n12277);
   U1421 : OAI21_X1 port map( B1 => n12307, B2 => n1805, A => n12275, ZN => 
                           n12280);
   U1422 : OAI21_X1 port map( B1 => n12403, B2 => n12280, A => n12281, ZN => 
                           n12276);
   U1423 : AOI21_X1 port map( B1 => n12277, B2 => n1808, A => n12276, ZN => 
                           n12296);
   U1424 : NOR3_X1 port map( A1 => n12278, A2 => n12296, A3 => n13225, ZN => 
                           n12285);
   U1425 : AOI22_X1 port map( A1 => n12388, A2 => n12280, B1 => n1808, B2 => 
                           n12279, ZN => n12298);
   U1426 : INV_X1 port map( A => n12281, ZN => n12297);
   U1427 : OAI22_X1 port map( A1 => n12298, A2 => n12297, B1 => n13225, B2 => 
                           n12282, ZN => n12284);
   U1428 : AOI22_X1 port map( A1 => n12286, A2 => n12285, B1 => n12284, B2 => 
                           n12283, ZN => n3863);
   U1429 : NAND2_X1 port map( A1 => n13224, A2 => n8694, ZN => n6932);
   U1430 : OAI22_X1 port map( A1 => n8801, A2 => n12287, B1 => n9166, B2 => 
                           n12303, ZN => n12294);
   U1431 : INV_X1 port map( A => n12288, ZN => n12311);
   U1432 : OAI22_X1 port map( A1 => n8677, A2 => n12311, B1 => n9167, B2 => 
                           n12323, ZN => n12293);
   U1433 : OAI222_X1 port map( A1 => n13191, A2 => n8889, B1 => n12300, B2 => 
                           n8960, C1 => n12289, C2 => n8676, ZN => n12290);
   U1434 : AOI21_X1 port map( B1 => n12290, B2 => n8902, A => n8835, ZN => 
                           n12291);
   U1435 : NAND2_X1 port map( A1 => n8589, A2 => n12291, ZN => n12292);
   U1436 : AOI221_X1 port map( B1 => n12294, B2 => n8969, C1 => n12293, C2 => 
                           n8969, A => n12292, ZN => n12295);
   U1437 : OAI211_X1 port map( C1 => n8834, C2 => n9208, A => n8944, B => 
                           n12295, ZN => OUTALU(23));
   U1438 : NAND2_X1 port map( A1 => DATA2(22), A2 => n12554, ZN => n12622);
   U1439 : OAI21_X1 port map( B1 => DATA2(22), B2 => n12554, A => n12622, ZN =>
                           n12691);
   U1440 : AOI22_X1 port map( A1 => n8696, A2 => n13224, B1 => n12535, B2 => 
                           n12691, ZN => n3861);
   U1441 : AOI21_X1 port map( B1 => n12298, B2 => n12297, A => n12296, ZN => 
                           n6935);
   U1442 : AOI22_X1 port map( A1 => n9186, A2 => n8544, B1 => n11337, B2 => 
                           n9014, ZN => n12299);
   U1443 : OAI21_X1 port map( B1 => n12300, B2 => n13208, A => n12299, ZN => 
                           n12301);
   U1444 : AOI21_X1 port map( B1 => n8852, B2 => n12302, A => n12301, ZN => 
                           n12306);
   U1445 : OAI222_X1 port map( A1 => n8677, A2 => n12323, B1 => n8801, B2 => 
                           n12303, C1 => n9166, C2 => n12311, ZN => n12304);
   U1446 : AOI211_X1 port map( C1 => n8969, C2 => n12304, A => n8587, B => 
                           n8892, ZN => n12305);
   U1447 : OAI211_X1 port map( C1 => n9100, C2 => n12306, A => n8588, B => 
                           n12305, ZN => OUTALU(22));
   U1448 : INV_X1 port map( A => DATA2(21), ZN => n12767);
   U1449 : AOI22_X1 port map( A1 => DATA1(21), A2 => DATA2(21), B1 => n12767, 
                           B2 => n12692, ZN => n12570);
   U1450 : AOI22_X1 port map( A1 => n12535, A2 => n12570, B1 => n6095, B2 => 
                           n8698, ZN => n3859);
   U1451 : AOI22_X1 port map( A1 => n12308, A2 => n1808, B1 => n12388, B2 => 
                           n12307, ZN => n12310);
   U1452 : AOI21_X1 port map( B1 => n12519, B2 => DATA2(21), A => n12518, ZN =>
                           n12309);
   U1453 : OAI22_X1 port map( A1 => n12310, A2 => n1805, B1 => n12309, B2 => 
                           n12692, ZN => n6949);
   U1454 : OAI22_X1 port map( A1 => n8801, A2 => n12311, B1 => n9166, B2 => 
                           n12323, ZN => n12312);
   U1455 : AOI211_X1 port map( C1 => n8969, C2 => n12312, A => n8584, B => 
                           n13217, ZN => n12314);
   U1456 : NAND3_X1 port map( A1 => n12392, A2 => n13162, A3 => n13204, ZN => 
                           n12313);
   U1457 : OAI211_X1 port map( C1 => n8963, C2 => n8586, A => n12314, B => 
                           n12313, ZN => OUTALU(21));
   U1458 : AOI22_X1 port map( A1 => n12388, A2 => n12316, B1 => n1808, B2 => 
                           n12317, ZN => n3858);
   U1459 : NOR2_X1 port map( A1 => DATA2(20), A2 => n12319, ZN => n12688);
   U1460 : NAND2_X1 port map( A1 => n12319, A2 => DATA2(20), ZN => n12620);
   U1461 : INV_X1 port map( A => n12620, ZN => n12634);
   U1462 : NOR2_X1 port map( A1 => n12688, A2 => n12634, ZN => n12564);
   U1463 : INV_X1 port map( A => n12564, ZN => n12315);
   U1464 : AOI22_X1 port map( A1 => n12535, A2 => n12315, B1 => n13224, B2 => 
                           n8700, ZN => n3856);
   U1465 : OAI22_X1 port map( A1 => n12317, A2 => n12406, B1 => n12403, B2 => 
                           n12316, ZN => n12318);
   U1466 : INV_X1 port map( A => n12318, ZN => n12321);
   U1467 : AOI21_X1 port map( B1 => n12519, B2 => DATA2(20), A => n12518, ZN =>
                           n12320);
   U1468 : OAI22_X1 port map( A1 => n12321, A2 => n1806, B1 => n12320, B2 => 
                           n12319, ZN => n6957);
   U1469 : AOI22_X1 port map( A1 => n13144, A2 => n12392, B1 => n12393, B2 => 
                           n13162, ZN => n12326);
   U1470 : OAI21_X1 port map( B1 => n8964, B2 => n8583, A => n8582, ZN => 
                           n12322);
   U1471 : NOR2_X1 port map( A1 => n8833, A2 => n12322, ZN => n12325);
   U1472 : OR3_X1 port map( A1 => n8801, A2 => n12323, A3 => n9109, ZN => 
                           n12324);
   U1473 : OAI211_X1 port map( C1 => n12326, C2 => n13203, A => n12325, B => 
                           n12324, ZN => OUTALU(20));
   U1474 : AOI211_X1 port map( C1 => n12531, C2 => n12333, A => n12328, B => 
                           n12327, ZN => n12330);
   U1475 : NOR2_X1 port map( A1 => n13088, A2 => n9222, ZN => n12637);
   U1476 : INV_X1 port map( A => n12637, ZN => n12593);
   U1477 : NOR2_X1 port map( A1 => DATA2(1), A2 => n11332, ZN => n12591);
   U1478 : INV_X1 port map( A => n12591, ZN => n12639);
   U1479 : AOI21_X1 port map( B1 => n12593, B2 => n12639, A => n1835, ZN => 
                           n12329);
   U1480 : AOI211_X1 port map( C1 => n8528, C2 => n13224, A => n12330, B => 
                           n12329, ZN => n3854);
   U1481 : AOI21_X1 port map( B1 => n12541, B2 => n12331, A => n12518, ZN => 
                           n12529);
   U1482 : OAI21_X1 port map( B1 => n13088, B2 => n12530, A => n12529, ZN => 
                           n4070);
   U1483 : NAND3_X1 port map( A1 => n9221, A2 => n12332, A3 => n12331, ZN => 
                           n4069);
   U1484 : OAI221_X1 port map( B1 => n12532, B2 => n12335, C1 => n12334, C2 => 
                           n12333, A => n7166, ZN => n3822);
   U1485 : OAI22_X1 port map( A1 => n13102, A2 => n11315, B1 => n12538, B2 => 
                           n13100, ZN => n12344);
   U1486 : NOR4_X1 port map( A1 => n12339, A2 => n12338, A3 => n12337, A4 => 
                           n12336, ZN => n12340);
   U1487 : OAI21_X1 port map( B1 => n11332, B2 => n12341, A => n12340, ZN => 
                           n12546);
   U1488 : AOI222_X1 port map( A1 => n12342, A2 => n11528, B1 => n12546, B2 => 
                           n13223, C1 => n12548, C2 => n1865, ZN => n12549);
   U1489 : OAI22_X1 port map( A1 => n13108, A2 => n12549, B1 => n1869, B2 => 
                           n13101, ZN => n12343);
   U1490 : AOI211_X1 port map( C1 => n1872, C2 => n12553, A => n12344, B => 
                           n12343, ZN => n7286);
   U1491 : OAI22_X1 port map( A1 => n8895, A2 => n8637, B1 => n13145, B2 => 
                           n13158, ZN => n12346);
   U1492 : OAI22_X1 port map( A1 => n9182, A2 => n8580, B1 => n9181, B2 => 
                           n8598, ZN => n12345);
   U1493 : AOI211_X1 port map( C1 => n13153, C2 => n13198, A => n12346, B => 
                           n12345, ZN => n12722);
   U1494 : OAI222_X1 port map( A1 => n8975, A2 => n12347, B1 => n9103, B2 => 
                           n12723, C1 => n8896, C2 => n12722, ZN => n12726);
   U1495 : AOI22_X1 port map( A1 => n9183, A2 => n12726, B1 => n9025, B2 => 
                           n12348, ZN => n12352);
   U1496 : INV_X1 port map( A => n12349, ZN => n12350);
   U1497 : AOI22_X1 port map( A1 => n9102, A2 => n12350, B1 => n8905, B2 => 
                           n12725, ZN => n12351);
   U1498 : OAI211_X1 port map( C1 => n12353, C2 => n9032, A => n12352, B => 
                           n12351, ZN => n12734);
   U1499 : AOI22_X1 port map( A1 => n9164, A2 => n12734, B1 => n12731, B2 => 
                           n13157, ZN => n12356);
   U1500 : AOI22_X1 port map( A1 => n9173, A2 => n12733, B1 => n8804, B2 => 
                           n12354, ZN => n12355);
   U1501 : OAI211_X1 port map( C1 => n12357, C2 => n13165, A => n12356, B => 
                           n12355, ZN => n12738);
   U1502 : AOI222_X1 port map( A1 => n12738, A2 => n8910, B1 => n12739, B2 => 
                           n9111, C1 => n12358, C2 => n9175, ZN => n12744);
   U1503 : OAI22_X1 port map( A1 => n9113, A2 => n12743, B1 => n8802, B2 => 
                           n12744, ZN => n12361);
   U1504 : OAI22_X1 port map( A1 => n12359, A2 => n13206, B1 => n8805, B2 => 
                           n12742, ZN => n12360);
   U1505 : AOI211_X1 port map( C1 => n9099, C2 => n12362, A => n12361, B => 
                           n12360, ZN => n12753);
   U1506 : INV_X1 port map( A => n12753, ZN => n12363);
   U1507 : AOI22_X1 port map( A1 => n9006, A2 => n8832, B1 => n8902, B2 => 
                           n12363, ZN => n12364);
   U1508 : NAND4_X1 port map( A1 => n8553, A2 => n8581, A3 => n8831, A4 => 
                           n12364, ZN => OUTALU(1));
   U1509 : INV_X1 port map( A => DATA2(19), ZN => n12769);
   U1510 : OAI21_X1 port map( B1 => n12530, B2 => n12769, A => n12466, ZN => 
                           n12365);
   U1511 : AOI22_X1 port map( A1 => DATA1(19), A2 => n12365, B1 => n6095, B2 =>
                           n8702, ZN => n3851);
   U1512 : NAND2_X1 port map( A1 => DATA1(19), A2 => n12769, ZN => n12685);
   U1513 : INV_X1 port map( A => n12685, ZN => n12577);
   U1514 : NOR2_X1 port map( A1 => DATA1(19), A2 => n12769, ZN => n12635);
   U1515 : OAI21_X1 port map( B1 => n12577, B2 => n12635, A => n12535, ZN => 
                           n4068);
   U1516 : INV_X1 port map( A => n12369, ZN => n12372);
   U1517 : AOI22_X1 port map( A1 => n12366, A2 => n1808, B1 => n12388, B2 => 
                           n12367, ZN => n12371);
   U1518 : OAI22_X1 port map( A1 => n12403, A2 => n12367, B1 => n12406, B2 => 
                           n12366, ZN => n12368);
   U1519 : INV_X1 port map( A => n12368, ZN => n12370);
   U1520 : AOI22_X1 port map( A1 => n12372, A2 => n12371, B1 => n12370, B2 => 
                           n12369, ZN => n7007);
   U1521 : AOI222_X1 port map( A1 => n12373, A2 => n13162, B1 => n12392, B2 => 
                           n13170, C1 => n12393, C2 => n13144, ZN => n12381);
   U1522 : INV_X1 port map( A => n12420, ZN => n12376);
   U1523 : AOI22_X1 port map( A1 => n8905, A2 => n12389, B1 => n9024, B2 => 
                           n12374, ZN => n12375);
   U1524 : OAI21_X1 port map( B1 => n12376, B2 => n13150, A => n12375, ZN => 
                           n12377);
   U1525 : AOI21_X1 port map( B1 => n9025, B2 => n12410, A => n12377, ZN => 
                           n12378);
   U1526 : OAI21_X1 port map( B1 => n9033, B2 => n12378, A => n8579, ZN => 
                           n12379);
   U1527 : NOR2_X1 port map( A1 => n8578, A2 => n12379, ZN => n12380);
   U1528 : OAI211_X1 port map( C1 => n12381, C2 => n13203, A => n8830, B => 
                           n12380, ZN => OUTALU(19));
   U1529 : INV_X1 port map( A => DATA2(18), ZN => n12770);
   U1530 : OAI21_X1 port map( B1 => n12530, B2 => n12770, A => n12466, ZN => 
                           n4067);
   U1531 : AOI211_X1 port map( C1 => n12383, C2 => n12386, A => n12382, B => 
                           n12406, ZN => n3850);
   U1532 : OAI22_X1 port map( A1 => n12687, A2 => DATA2(18), B1 => n12770, B2 
                           => DATA1(18), ZN => n12615);
   U1533 : AOI22_X1 port map( A1 => n8704, A2 => n13224, B1 => n12535, B2 => 
                           n12615, ZN => n3849);
   U1534 : AOI21_X1 port map( B1 => n12386, B2 => n12385, A => n12384, ZN => 
                           n12387);
   U1535 : NAND2_X1 port map( A1 => n12388, A2 => n12387, ZN => n3848);
   U1536 : AOI222_X1 port map( A1 => n12410, A2 => n8905, B1 => n12420, B2 => 
                           n9025, C1 => n12389, C2 => n9024, ZN => n12401);
   U1537 : NAND2_X1 port map( A1 => n9003, A2 => n8829, ZN => n12390);
   U1538 : NAND3_X1 port map( A1 => n8575, A2 => n8576, A3 => n12390, ZN => 
                           n12391);
   U1539 : NOR2_X1 port map( A1 => n8577, A2 => n12391, ZN => n12400);
   U1540 : AOI22_X1 port map( A1 => n12393, A2 => n8806, B1 => n12392, B2 => 
                           n9105, ZN => n12394);
   U1541 : INV_X1 port map( A => n12394, ZN => n12398);
   U1542 : OAI22_X1 port map( A1 => n12396, A2 => n13164, B1 => n12395, B2 => 
                           n13142, ZN => n12397);
   U1543 : OAI21_X1 port map( B1 => n12398, B2 => n12397, A => n13161, ZN => 
                           n12399);
   U1544 : OAI211_X1 port map( C1 => n9109, C2 => n12401, A => n12400, B => 
                           n12399, ZN => OUTALU(18));
   U1545 : INV_X1 port map( A => DATA2(17), ZN => n12771);
   U1546 : NAND2_X1 port map( A1 => n12771, A2 => DATA1(17), ZN => n12587);
   U1547 : NAND2_X1 port map( A1 => DATA2(17), A2 => n12402, ZN => n12681);
   U1548 : NAND2_X1 port map( A1 => n12587, A2 => n12681, ZN => n12559);
   U1549 : AOI22_X1 port map( A1 => n12535, A2 => n12559, B1 => n13224, B2 => 
                           n8706, ZN => n3847);
   U1550 : AOI211_X1 port map( C1 => n12405, C2 => n12408, A => n12404, B => 
                           n12403, ZN => n3846);
   U1551 : AOI211_X1 port map( C1 => n12409, C2 => n12408, A => n12407, B => 
                           n12406, ZN => n3845);
   U1552 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n12477, 
                           ZN => n3844);
   U1553 : AOI22_X1 port map( A1 => n12410, A2 => n9024, B1 => n12420, B2 => 
                           n8905, ZN => n12411);
   U1554 : INV_X1 port map( A => n12411, ZN => n12412);
   U1555 : AOI211_X1 port map( C1 => n8969, C2 => n12412, A => n8573, B => 
                           n8572, ZN => n12414);
   U1556 : NAND3_X1 port map( A1 => n9218, A2 => n8902, A3 => n12417, ZN => 
                           n12413);
   U1557 : NAND4_X1 port map( A1 => n8574, A2 => n8828, A3 => n12414, A4 => 
                           n12413, ZN => OUTALU(17));
   U1558 : INV_X1 port map( A => DATA2(16), ZN => n12772);
   U1559 : OAI21_X1 port map( B1 => n12530, B2 => n12772, A => n12466, ZN => 
                           n4066);
   U1560 : NAND2_X1 port map( A1 => DATA1(16), A2 => n12772, ZN => n12679);
   U1561 : OAI21_X1 port map( B1 => DATA1(16), B2 => n12772, A => n12679, ZN =>
                           n12555);
   U1562 : AOI22_X1 port map( A1 => n8708, A2 => n13224, B1 => n12535, B2 => 
                           n12555, ZN => n3843);
   U1563 : NOR2_X1 port map( A1 => n9170, A2 => n8971, ZN => n12415);
   U1564 : AOI21_X1 port map( B1 => n9004, B2 => n8827, A => n12415, ZN => 
                           n12423);
   U1565 : AOI22_X1 port map( A1 => n8907, A2 => n12417, B1 => n9218, B2 => 
                           n12416, ZN => n12418);
   U1566 : OAI21_X1 port map( B1 => n9100, B2 => n12418, A => n8571, ZN => 
                           n12419);
   U1567 : NOR2_X1 port map( A1 => n8943, A2 => n12419, ZN => n12422);
   U1568 : NAND3_X1 port map( A1 => n9024, A2 => n8969, A3 => n12420, ZN => 
                           n12421);
   U1569 : NAND3_X1 port map( A1 => n12423, A2 => n12422, A3 => n12421, ZN => 
                           OUTALU(16));
   U1570 : NAND2_X1 port map( A1 => DATA1(15), A2 => n12773, ZN => n12674);
   U1571 : NAND2_X1 port map( A1 => DATA2(15), A2 => n12424, ZN => n12676);
   U1572 : AND2_X1 port map( A1 => n12674, A2 => n12676, ZN => n12574);
   U1573 : NAND3_X1 port map( A1 => DATA1(15), A2 => DATA2(15), A3 => n12477, 
                           ZN => n12438);
   U1574 : INV_X1 port map( A => n12504, ZN => n12502);
   U1575 : INV_X1 port map( A => n12516, ZN => n12425);
   U1576 : AOI21_X1 port map( B1 => n12514, B2 => n12425, A => n12515, ZN => 
                           n12426);
   U1577 : INV_X1 port map( A => n12426, ZN => n12512);
   U1578 : NAND2_X1 port map( A1 => n12512, A2 => n12427, ZN => n12501);
   U1579 : NAND2_X1 port map( A1 => n12502, A2 => n12501, ZN => n12428);
   U1580 : NAND2_X1 port map( A1 => n12429, A2 => n12428, ZN => n12479);
   U1581 : AOI21_X1 port map( B1 => n12431, B2 => n12479, A => n12430, ZN => 
                           n12449);
   U1582 : NAND2_X1 port map( A1 => n12449, A2 => n12448, ZN => n12455);
   U1583 : INV_X1 port map( A => n12455, ZN => n12433);
   U1584 : OAI21_X1 port map( B1 => n12433, B2 => n12451, A => n12432, ZN => 
                           n12436);
   U1585 : AOI21_X1 port map( B1 => n12442, B2 => n12436, A => n12434, ZN => 
                           n12435);
   U1586 : OAI21_X1 port map( B1 => n12442, B2 => n12436, A => n12435, ZN => 
                           n12437);
   U1587 : OAI211_X1 port map( C1 => n12574, C2 => n1835, A => n12438, B => 
                           n12437, ZN => n3842);
   U1588 : INV_X1 port map( A => n12439, ZN => n12441);
   U1589 : INV_X1 port map( A => n12442, ZN => n12440);
   U1590 : INV_X1 port map( A => n12510, ZN => n12482);
   U1591 : OAI221_X1 port map( B1 => n12442, B2 => n12441, C1 => n12440, C2 => 
                           n12439, A => n12482, ZN => n3821);
   U1592 : INV_X1 port map( A => n12443, ZN => n12444);
   U1593 : AOI22_X1 port map( A1 => n13171, A2 => n12460, B1 => n13147, B2 => 
                           n12444, ZN => n12447);
   U1594 : AOI211_X1 port map( C1 => n8710, C2 => n9210, A => n8570, B => 
                           n13218, ZN => n12446);
   U1595 : OR3_X1 port map( A1 => n8897, A2 => n12488, A3 => n9100, ZN => 
                           n12445);
   U1596 : OAI211_X1 port map( C1 => n12447, C2 => n13205, A => n12446, B => 
                           n12445, ZN => OUTALU(15));
   U1597 : INV_X1 port map( A => n12448, ZN => n12452);
   U1598 : AOI22_X1 port map( A1 => n12450, A2 => n12482, B1 => n7147, B2 => 
                           n12449, ZN => n12467);
   U1599 : NOR3_X1 port map( A1 => n12452, A2 => n12467, A3 => n12451, ZN => 
                           n4065);
   U1600 : NAND2_X1 port map( A1 => n11309, A2 => n8990, ZN => n12453);
   U1601 : OAI21_X1 port map( B1 => n11309, B2 => n8990, A => n12453, ZN => 
                           n13007);
   U1602 : NOR3_X1 port map( A1 => n11301, A2 => n11340, A3 => n13007, ZN => 
                           n3020);
   U1603 : AOI221_X1 port map( B1 => n11301, B2 => n11340, C1 => n13007, C2 => 
                           n11340, A => n3020, ZN => n4200);
   U1604 : AOI22_X1 port map( A1 => n7147, A2 => n12455, B1 => n12482, B2 => 
                           n12454, ZN => n12458);
   U1605 : OAI22_X1 port map( A1 => n12774, A2 => DATA1(14), B1 => n12675, B2 
                           => DATA2(14), ZN => n12608);
   U1606 : AOI22_X1 port map( A1 => n8824, A2 => n13224, B1 => n12535, B2 => 
                           n12608, ZN => n12457);
   U1607 : OAI211_X1 port map( C1 => n12518, C2 => n12519, A => DATA1(14), B =>
                           DATA2(14), ZN => n12456);
   U1608 : OAI211_X1 port map( C1 => n12459, C2 => n12458, A => n12457, B => 
                           n12456, ZN => n7086);
   U1609 : NAND2_X1 port map( A1 => n12460, A2 => n13147, ZN => n12463);
   U1610 : OAI22_X1 port map( A1 => n12489, A2 => n13143, B1 => n12488, B2 => 
                           n13148, ZN => n12461);
   U1611 : AOI211_X1 port map( C1 => n13161, C2 => n12461, A => n8826, B => 
                           n8942, ZN => n12462);
   U1612 : OAI21_X1 port map( B1 => n9033, B2 => n12463, A => n12462, ZN => 
                           OUTALU(14));
   U1613 : INV_X1 port map( A => n12479, ZN => n12478);
   U1614 : NOR3_X1 port map( A1 => n12478, A2 => n12485, A3 => n13225, ZN => 
                           n12464);
   U1615 : OAI211_X1 port map( C1 => n12484, C2 => n12465, A => n12464, B => 
                           n12468, ZN => n3838);
   U1616 : OAI21_X1 port map( B1 => n12530, B2 => n12775, A => n12466, ZN => 
                           n4064);
   U1617 : AOI21_X1 port map( B1 => n12469, B2 => n12468, A => n12467, ZN => 
                           n4063);
   U1618 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12775, ZN => n12667);
   U1619 : NAND2_X1 port map( A1 => DATA2(13), A2 => n12470, ZN => n12669);
   U1620 : NAND2_X1 port map( A1 => n12667, A2 => n12669, ZN => n12558);
   U1621 : AOI22_X1 port map( A1 => n12535, A2 => n12558, B1 => n13224, B2 => 
                           n8727, ZN => n3837);
   U1622 : OAI222_X1 port map( A1 => n13143, A2 => n12490, B1 => n13148, B2 => 
                           n12489, C1 => n13180, C2 => n12488, ZN => n12471);
   U1623 : AOI211_X1 port map( C1 => n13161, C2 => n12471, A => n8821, B => 
                           n13219, ZN => n12476);
   U1624 : OAI22_X1 port map( A1 => n8972, A2 => n12526, B1 => n8849, B2 => 
                           n13142, ZN => n12473);
   U1625 : OAI22_X1 port map( A1 => n9022, A2 => n8604, B1 => n13154, B2 => 
                           n13164, ZN => n12472);
   U1626 : OAI21_X1 port map( B1 => n12473, B2 => n12472, A => n13207, ZN => 
                           n12475);
   U1627 : NAND2_X1 port map( A1 => n9005, A2 => n8822, ZN => n12474);
   U1628 : NAND4_X1 port map( A1 => n8823, A2 => n12476, A3 => n12475, A4 => 
                           n12474, ZN => OUTALU(13));
   U1629 : OAI22_X1 port map( A1 => n12776, A2 => n12668, B1 => DATA1(12), B2 
                           => DATA2(12), ZN => n12604);
   U1630 : NAND3_X1 port map( A1 => DATA1(12), A2 => DATA2(12), A3 => n12477, 
                           ZN => n12481);
   U1631 : INV_X1 port map( A => n12485, ZN => n12483);
   U1632 : OAI221_X1 port map( B1 => n12483, B2 => n12479, C1 => n12485, C2 => 
                           n12478, A => n7147, ZN => n12480);
   U1633 : OAI211_X1 port map( C1 => n12604, C2 => n1835, A => n12481, B => 
                           n12480, ZN => n3836);
   U1634 : INV_X1 port map( A => n12484, ZN => n12486);
   U1635 : OAI221_X1 port map( B1 => n12486, B2 => n12485, C1 => n12484, C2 => 
                           n12483, A => n12482, ZN => n3835);
   U1636 : OAI222_X1 port map( A1 => n9022, A2 => n12526, B1 => n9181, B2 => 
                           n8604, C1 => n9023, C2 => n8849, ZN => n12487);
   U1637 : AOI22_X1 port map( A1 => n9210, A2 => n8867, B1 => n8969, B2 => 
                           n12487, ZN => n12495);
   U1638 : OAI22_X1 port map( A1 => n12489, A2 => n13180, B1 => n12488, B2 => 
                           n13150, ZN => n12493);
   U1639 : OAI22_X1 port map( A1 => n12491, A2 => n13143, B1 => n12490, B2 => 
                           n13148, ZN => n12492);
   U1640 : OAI21_X1 port map( B1 => n12493, B2 => n12492, A => n13161, ZN => 
                           n12494);
   U1641 : NAND4_X1 port map( A1 => n8551, A2 => n12495, A3 => n12494, A4 => 
                           n13213, ZN => OUTALU(12));
   U1642 : NOR3_X1 port map( A1 => n12496, A2 => n12497, A3 => n12777, ZN => 
                           n12500);
   U1643 : NOR2_X1 port map( A1 => DATA2(11), A2 => n12497, ZN => n12605);
   U1644 : NOR2_X1 port map( A1 => DATA1(11), A2 => n12777, ZN => n12664);
   U1645 : OAI21_X1 port map( B1 => n12605, B2 => n12664, A => n12535, ZN => 
                           n12498);
   U1646 : INV_X1 port map( A => n12498, ZN => n12499);
   U1647 : AOI211_X1 port map( C1 => n8744, C2 => n13224, A => n12500, B => 
                           n12499, ZN => n4062);
   U1648 : XOR2_X1 port map( A => n12502, B => n12501, Z => n4199);
   U1649 : INV_X1 port map( A => n12505, ZN => n12503);
   U1650 : AOI221_X1 port map( B1 => n12505, B2 => n12504, C1 => n12503, C2 => 
                           n12502, A => n12510, ZN => n3820);
   U1651 : OAI22_X1 port map( A1 => n9181, A2 => n12526, B1 => n9023, B2 => 
                           n8604, ZN => n12506);
   U1652 : AOI22_X1 port map( A1 => n8969, A2 => n12506, B1 => n9108, B2 => 
                           n8941, ZN => n12509);
   U1653 : NOR3_X1 port map( A1 => n8801, A2 => n12523, A3 => n9100, ZN => 
                           n12507);
   U1654 : NOR2_X1 port map( A1 => n12507, A2 => n8550, ZN => n12508);
   U1655 : NAND3_X1 port map( A1 => n8567, A2 => n12509, A3 => n12508, ZN => 
                           OUTALU(11));
   U1656 : NOR2_X1 port map( A1 => n12511, A2 => n12510, ZN => n12517);
   U1657 : AOI21_X1 port map( B1 => n12512, B2 => n7147, A => n12517, ZN => 
                           n12513);
   U1658 : AOI21_X1 port map( B1 => n12514, B2 => n12515, A => n12513, ZN => 
                           n3834);
   U1659 : NAND3_X1 port map( A1 => n7147, A2 => n12516, A3 => n12515, ZN => 
                           n4061);
   U1660 : INV_X1 port map( A => n12517, ZN => n12521);
   U1661 : AOI22_X1 port map( A1 => DATA2(10), A2 => n12571, B1 => DATA1(10), 
                           B2 => n12778, ZN => n12660);
   U1662 : AOI21_X1 port map( B1 => n12519, B2 => DATA2(10), A => n12518, ZN =>
                           n12520);
   U1663 : OAI222_X1 port map( A1 => n12522, A2 => n12521, B1 => n1835, B2 => 
                           n12660, C1 => n12571, C2 => n12520, ZN => n7150);
   U1664 : NAND2_X1 port map( A1 => n13224, A2 => n8871, ZN => n7153);
   U1665 : OAI22_X1 port map( A1 => n8801, A2 => n12524, B1 => n12523, B2 => 
                           n9036, ZN => n12525);
   U1666 : AOI211_X1 port map( C1 => n8902, C2 => n12525, A => n8566, B => 
                           n8819, ZN => n12528);
   U1667 : OR3_X1 port map( A1 => n9023, A2 => n12526, A3 => n9033, ZN => 
                           n12527);
   U1668 : NAND4_X1 port map( A1 => n8820, A2 => n8940, A3 => n12528, A4 => 
                           n12527, ZN => OUTALU(10));
   U1669 : OAI21_X1 port map( B1 => n13082, B2 => n12530, A => n12529, ZN => 
                           n12536);
   U1670 : NAND2_X1 port map( A1 => n13082, A2 => n9221, ZN => n12638);
   U1671 : NAND2_X1 port map( A1 => DATA2(0), A2 => n13173, ZN => n12592);
   U1672 : NAND2_X1 port map( A1 => n12638, A2 => n12592, ZN => n12576);
   U1673 : NOR2_X1 port map( A1 => n12532, A2 => n12531, ZN => n12537);
   U1674 : INV_X1 port map( A => n12537, ZN => n12534);
   U1675 : AOI222_X1 port map( A1 => n12536, A2 => n9221, B1 => n12576, B2 => 
                           n12535, C1 => n12534, C2 => n12533, ZN => n4060);
   U1676 : AOI22_X1 port map( A1 => n13224, A2 => n8933, B1 => n7166, B2 => 
                           n12537, ZN => n3831);
   U1677 : OAI22_X1 port map( A1 => n1869, A2 => n13102, B1 => n12538, B2 => 
                           n13133, ZN => n12552);
   U1678 : AOI211_X1 port map( C1 => n12541, C2 => n9221, A => n12540, B => 
                           n12539, ZN => n12544);
   U1679 : INV_X1 port map( A => n12542, ZN => n12543);
   U1680 : OAI211_X1 port map( C1 => n9205, C2 => n12545, A => n12544, B => 
                           n12543, ZN => n12547);
   U1681 : AOI222_X1 port map( A1 => n12548, A2 => n11528, B1 => n12547, B2 => 
                           n13223, C1 => n12546, C2 => n1865, ZN => n12550);
   U1682 : OAI22_X1 port map( A1 => n13108, A2 => n12550, B1 => n12549, B2 => 
                           n13100, ZN => n12551);
   U1683 : AOI211_X1 port map( C1 => n13123, C2 => n12553, A => n12552, B => 
                           n12551, ZN => n7285);
   U1684 : OAI22_X1 port map( A1 => DATA2(22), A2 => n12554, B1 => DATA2(23), 
                           B2 => n1846, ZN => n12697);
   U1685 : OR4_X1 port map( A1 => n12608, A2 => n12555, A3 => n12615, A4 => 
                           n12697, ZN => n12584);
   U1686 : AOI21_X1 port map( B1 => DATA1(10), B2 => n12778, A => n12605, ZN =>
                           n12666);
   U1687 : INV_X1 port map( A => n12556, ZN => n12696);
   U1688 : AOI21_X1 port map( B1 => DATA1(26), B2 => n12762, A => n12627, ZN =>
                           n12708);
   U1689 : NAND4_X1 port map( A1 => n12666, A2 => n12604, A3 => n12696, A4 => 
                           n12708, ZN => n12583);
   U1690 : NOR3_X1 port map( A1 => n12637, A2 => n12591, A3 => n12557, ZN => 
                           n12563);
   U1691 : NOR4_X1 port map( A1 => n12561, A2 => n12560, A3 => n12559, A4 => 
                           n12558, ZN => n12562);
   U1692 : NAND4_X1 port map( A1 => n12565, A2 => n12564, A3 => n12563, A4 => 
                           n12562, ZN => n12582);
   U1693 : AOI21_X1 port map( B1 => n12588, B2 => DATA2(7), A => n12599, ZN => 
                           n12566);
   U1694 : INV_X1 port map( A => n12566, ZN => n12657);
   U1695 : NAND4_X1 port map( A1 => n12640, A2 => n12655, A3 => n12567, A4 => 
                           n12622, ZN => n12568);
   U1696 : NOR4_X1 port map( A1 => n12570, A2 => n12569, A3 => n12657, A4 => 
                           n12568, ZN => n12579);
   U1697 : AOI21_X1 port map( B1 => DATA2(10), B2 => n12571, A => n12664, ZN =>
                           n12607);
   U1698 : AOI21_X1 port map( B1 => DATA2(26), B2 => n12572, A => n12706, ZN =>
                           n12629);
   U1699 : NAND4_X1 port map( A1 => n12607, A2 => n12629, A3 => n12574, A4 => 
                           n12573, ZN => n12575);
   U1700 : NOR4_X1 port map( A1 => n12577, A2 => n12635, A3 => n12576, A4 => 
                           n12575, ZN => n12578);
   U1701 : NAND4_X1 port map( A1 => n12580, A2 => n12712, A3 => n12579, A4 => 
                           n12578, ZN => n12581);
   U1702 : NOR4_X1 port map( A1 => n12584, A2 => n12583, A3 => n12582, A4 => 
                           n12581, ZN => n7326);
   U1703 : AOI21_X1 port map( B1 => DATA2(30), B2 => n12586, A => n12585, ZN =>
                           n7333);
   U1704 : INV_X1 port map( A => n12587, ZN => n12684);
   U1705 : AOI22_X1 port map( A1 => DATA2(7), A2 => n12588, B1 => DATA2(6), B2 
                           => n12651, ZN => n12601);
   U1706 : INV_X1 port map( A => n12589, ZN => n12646);
   U1707 : AOI211_X1 port map( C1 => n12593, C2 => n12592, A => n12591, B => 
                           n12590, ZN => n12595);
   U1708 : OAI21_X1 port map( B1 => n9223, B2 => n13077, A => n12643, ZN => 
                           n12594);
   U1709 : OAI21_X1 port map( B1 => n12595, B2 => n12594, A => n12648, ZN => 
                           n12596);
   U1710 : OAI21_X1 port map( B1 => n12646, B2 => n12596, A => n12644, ZN => 
                           n12598);
   U1711 : INV_X1 port map( A => n12597, ZN => n12647);
   U1712 : OAI211_X1 port map( C1 => n12650, C2 => n12598, A => n12655, B => 
                           n12647, ZN => n12600);
   U1713 : AOI211_X1 port map( C1 => n12601, C2 => n12600, A => n12653, B => 
                           n12599, ZN => n12603);
   U1714 : OAI21_X1 port map( B1 => DATA1(8), B2 => n12780, A => n12659, ZN => 
                           n12602);
   U1715 : OAI211_X1 port map( C1 => n12603, C2 => n12602, A => n12660, B => 
                           n12636, ZN => n12606);
   U1716 : INV_X1 port map( A => n12604, ZN => n12663);
   U1717 : AOI211_X1 port map( C1 => n12607, C2 => n12606, A => n12605, B => 
                           n12663, ZN => n12610);
   U1718 : OAI21_X1 port map( B1 => DATA1(12), B2 => n12776, A => n12669, ZN =>
                           n12609);
   U1719 : INV_X1 port map( A => n12608, ZN => n12670);
   U1720 : OAI211_X1 port map( C1 => n12610, C2 => n12609, A => n12670, B => 
                           n12667, ZN => n12611);
   U1721 : OAI211_X1 port map( C1 => DATA1(14), C2 => n12774, A => n12676, B =>
                           n12611, ZN => n12612);
   U1722 : NAND3_X1 port map( A1 => n12679, A2 => n12674, A3 => n12612, ZN => 
                           n12614);
   U1723 : NAND2_X1 port map( A1 => DATA2(16), A2 => n12613, ZN => n12677);
   U1724 : NAND3_X1 port map( A1 => n12681, A2 => n12614, A3 => n12677, ZN => 
                           n12616);
   U1725 : INV_X1 port map( A => n12615, ZN => n12682);
   U1726 : NAND2_X1 port map( A1 => n12616, A2 => n12682, ZN => n12617);
   U1727 : OAI22_X1 port map( A1 => n12684, A2 => n12617, B1 => DATA1(18), B2 
                           => n12770, ZN => n12618);
   U1728 : OAI21_X1 port map( B1 => n12635, B2 => n12618, A => n12685, ZN => 
                           n12619);
   U1729 : AOI21_X1 port map( B1 => n12620, B2 => n12619, A => n12688, ZN => 
                           n12621);
   U1730 : AOI222_X1 port map( A1 => DATA2(21), A2 => n12621, B1 => DATA2(21), 
                           B2 => n12692, C1 => n12621, C2 => n12692, ZN => 
                           n12623);
   U1731 : OAI211_X1 port map( C1 => n12691, C2 => n12623, A => n12622, B => 
                           n12695, ZN => n12624);
   U1732 : OAI211_X1 port map( C1 => DATA2(23), C2 => n1846, A => n12696, B => 
                           n12624, ZN => n12625);
   U1733 : OAI211_X1 port map( C1 => DATA1(24), C2 => n12764, A => n12625, B =>
                           n12701, ZN => n12626);
   U1734 : NAND3_X1 port map( A1 => n12702, A2 => n12633, A3 => n12626, ZN => 
                           n12628);
   U1735 : AOI211_X1 port map( C1 => n12629, C2 => n12628, A => n12627, B => 
                           n12705, ZN => n12631);
   U1736 : OAI21_X1 port map( B1 => DATA1(28), B2 => n12760, A => n12711, ZN =>
                           n12630);
   U1737 : OAI211_X1 port map( C1 => n12631, C2 => n12630, A => n12712, B => 
                           n12709, ZN => n7332);
   U1738 : AOI21_X1 port map( B1 => DATA1(30), B2 => n12758, A => n12632, ZN =>
                           n7340);
   U1739 : INV_X1 port map( A => n12633, ZN => n12704);
   U1740 : NOR2_X1 port map( A1 => n12635, A2 => n12634, ZN => n12690);
   U1741 : INV_X1 port map( A => n12636, ZN => n12662);
   U1742 : AOI21_X1 port map( B1 => n12639, B2 => n12638, A => n12637, ZN => 
                           n12641);
   U1743 : AOI22_X1 port map( A1 => n13077, A2 => n13177, B1 => n12641, B2 => 
                           n12640, ZN => n12642);
   U1744 : INV_X1 port map( A => n12642, ZN => n12645);
   U1745 : OAI211_X1 port map( C1 => n12646, C2 => n12645, A => n12644, B => 
                           n12643, ZN => n12649);
   U1746 : OAI221_X1 port map( B1 => n12650, B2 => n12649, C1 => n12650, C2 => 
                           n12648, A => n12647, ZN => n12654);
   U1747 : NOR2_X1 port map( A1 => DATA2(6), A2 => n12651, ZN => n12652);
   U1748 : AOI211_X1 port map( C1 => n12655, C2 => n12654, A => n12653, B => 
                           n12652, ZN => n12658);
   U1749 : OAI22_X1 port map( A1 => n12658, A2 => n12657, B1 => DATA2(8), B2 =>
                           n12656, ZN => n12661);
   U1750 : OAI211_X1 port map( C1 => n12662, C2 => n12661, A => n12660, B => 
                           n12659, ZN => n12665);
   U1751 : AOI211_X1 port map( C1 => n12666, C2 => n12665, A => n12664, B => 
                           n12663, ZN => n12672);
   U1752 : OAI21_X1 port map( B1 => DATA2(12), B2 => n12668, A => n12667, ZN =>
                           n12671);
   U1753 : OAI211_X1 port map( C1 => n12672, C2 => n12671, A => n12670, B => 
                           n12669, ZN => n12673);
   U1754 : OAI211_X1 port map( C1 => DATA2(14), C2 => n12675, A => n12674, B =>
                           n12673, ZN => n12678);
   U1755 : NAND3_X1 port map( A1 => n12678, A2 => n12677, A3 => n12676, ZN => 
                           n12680);
   U1756 : NAND2_X1 port map( A1 => n12680, A2 => n12679, ZN => n12683);
   U1757 : OAI211_X1 port map( C1 => n12684, C2 => n12683, A => n12682, B => 
                           n12681, ZN => n12686);
   U1758 : OAI211_X1 port map( C1 => DATA2(18), C2 => n12687, A => n12686, B =>
                           n12685, ZN => n12689);
   U1759 : AOI21_X1 port map( B1 => n12690, B2 => n12689, A => n12688, ZN => 
                           n12694);
   U1760 : NAND2_X1 port map( A1 => n12767, A2 => DATA1(21), ZN => n12693);
   U1761 : AOI221_X1 port map( B1 => n12694, B2 => n12693, C1 => DATA2(21), C2 
                           => n12692, A => n12691, ZN => n12698);
   U1762 : OAI211_X1 port map( C1 => n12698, C2 => n12697, A => n12696, B => 
                           n12695, ZN => n12699);
   U1763 : OAI21_X1 port map( B1 => DATA2(24), B2 => n12700, A => n12699, ZN =>
                           n12703);
   U1764 : OAI211_X1 port map( C1 => n12704, C2 => n12703, A => n12702, B => 
                           n12701, ZN => n12707);
   U1765 : AOI211_X1 port map( C1 => n12708, C2 => n12707, A => n12706, B => 
                           n12705, ZN => n12714);
   U1766 : OAI21_X1 port map( B1 => DATA2(28), B2 => n12710, A => n12709, ZN =>
                           n12713);
   U1767 : OAI211_X1 port map( C1 => n12714, C2 => n12713, A => n12712, B => 
                           n12711, ZN => n7339);
   U1768 : NAND2_X1 port map( A1 => n8626, A2 => n9000, ZN => n12754);
   U1769 : NAND4_X1 port map( A1 => n8563, A2 => n8597, A3 => n9190, A4 => 
                           n8939, ZN => n12715);
   U1770 : NAND2_X1 port map( A1 => n9212, A2 => n12715, ZN => n12716);
   U1771 : AOI211_X1 port map( C1 => n8999, C2 => n12716, A => n8998, B => 
                           n9214, ZN => n12751);
   U1772 : AOI22_X1 port map( A1 => n9179, A2 => n9001, B1 => n8816, B2 => 
                           n8817, ZN => n12718);
   U1773 : OAI221_X1 port map( B1 => n8949, B2 => n8815, C1 => n8949, C2 => 
                           n8562, A => n9007, ZN => n12717);
   U1774 : OAI211_X1 port map( C1 => n9000, C2 => n12718, A => n9213, B => 
                           n12717, ZN => n12750);
   U1775 : OAI22_X1 port map( A1 => n9020, A2 => n8630, B1 => n13190, B2 => 
                           n13158, ZN => n12720);
   U1776 : OAI22_X1 port map( A1 => n9182, A2 => n8564, B1 => n9181, B2 => 
                           n8580, ZN => n12719);
   U1777 : AOI211_X1 port map( C1 => n13153, C2 => n13200, A => n12720, B => 
                           n12719, ZN => n12721);
   U1778 : OAI222_X1 port map( A1 => n8975, A2 => n12723, B1 => n9103, B2 => 
                           n12722, C1 => n8896, C2 => n12721, ZN => n12724);
   U1779 : AOI22_X1 port map( A1 => n9162, A2 => n12725, B1 => n9183, B2 => 
                           n12724, ZN => n12729);
   U1780 : AOI22_X1 port map( A1 => n9102, A2 => n12727, B1 => n8905, B2 => 
                           n12726, ZN => n12728);
   U1781 : OAI211_X1 port map( C1 => n9107, C2 => n12730, A => n12729, B => 
                           n12728, ZN => n12732);
   U1782 : AOI22_X1 port map( A1 => n9164, A2 => n12732, B1 => n13178, B2 => 
                           n12731, ZN => n12736);
   U1783 : AOI22_X1 port map( A1 => n8898, A2 => n12734, B1 => n8804, B2 => 
                           n12733, ZN => n12735);
   U1784 : OAI211_X1 port map( C1 => n12737, C2 => n13165, A => n12736, B => 
                           n12735, ZN => n12740);
   U1785 : AOI222_X1 port map( A1 => n12740, A2 => n8910, B1 => n12739, B2 => 
                           n9175, C1 => n12738, C2 => n9111, ZN => n12741);
   U1786 : OAI22_X1 port map( A1 => n12742, A2 => n9037, B1 => n8802, B2 => 
                           n12741, ZN => n12746);
   U1787 : OAI22_X1 port map( A1 => n8805, A2 => n12744, B1 => n12743, B2 => 
                           n13206, ZN => n12745);
   U1788 : AOI211_X1 port map( C1 => n9099, C2 => n12747, A => n12746, B => 
                           n12745, ZN => n12748);
   U1789 : OAI211_X1 port map( C1 => n12748, C2 => n13203, A => n8818, B => 
                           n8565, ZN => n12749);
   U1790 : AOI21_X1 port map( B1 => n12751, B2 => n12750, A => n12749, ZN => 
                           n12752);
   U1791 : OAI21_X1 port map( B1 => n12754, B2 => n12753, A => n12752, ZN => 
                           OUTALU(0));
   U1792 : NAND2_X1 port map( A1 => n12756, A2 => n12755, ZN => n12787);
   U1793 : CLKBUF_X1 port map( A => n12787, Z => n12782);
   U1794 : NAND2_X1 port map( A1 => n12756, A2 => FUNC(3), ZN => n12786);
   U1795 : AOI22_X1 port map( A1 => DATA2(31), A2 => n12782, B1 => n12781, B2 
                           => n12757, ZN => N2548);
   U1796 : AOI22_X1 port map( A1 => DATA2(30), A2 => n12787, B1 => n12786, B2 
                           => n12758, ZN => N2547);
   U1797 : AOI22_X1 port map( A1 => DATA2(29), A2 => n12782, B1 => n12781, B2 
                           => n12759, ZN => N2546);
   U1798 : AOI22_X1 port map( A1 => DATA2(28), A2 => n12787, B1 => n12786, B2 
                           => n12760, ZN => N2545);
   U1799 : AOI22_X1 port map( A1 => DATA2(27), A2 => n12782, B1 => n12781, B2 
                           => n12761, ZN => N2544);
   U1800 : AOI22_X1 port map( A1 => DATA2(26), A2 => n12787, B1 => n12786, B2 
                           => n12762, ZN => N2543);
   U1801 : AOI22_X1 port map( A1 => DATA2(25), A2 => n12782, B1 => n12781, B2 
                           => n12763, ZN => N2542);
   U1802 : AOI22_X1 port map( A1 => DATA2(24), A2 => n12787, B1 => n12786, B2 
                           => n12764, ZN => N2541);
   U1803 : AOI22_X1 port map( A1 => DATA2(23), A2 => n12782, B1 => n12781, B2 
                           => n12765, ZN => N2540);
   U1804 : AOI22_X1 port map( A1 => DATA2(22), A2 => n12787, B1 => n12786, B2 
                           => n12766, ZN => N2539);
   U1805 : AOI22_X1 port map( A1 => DATA2(21), A2 => n12787, B1 => n12786, B2 
                           => n12767, ZN => N2538);
   U1806 : INV_X1 port map( A => DATA2(20), ZN => n12768);
   U1807 : AOI22_X1 port map( A1 => DATA2(20), A2 => n12787, B1 => n12786, B2 
                           => n12768, ZN => N2537);
   U1808 : AOI22_X1 port map( A1 => DATA2(19), A2 => n12782, B1 => n12781, B2 
                           => n12769, ZN => N2536);
   U1809 : AOI22_X1 port map( A1 => DATA2(18), A2 => n12782, B1 => n12781, B2 
                           => n12770, ZN => N2535);
   U1810 : AOI22_X1 port map( A1 => DATA2(17), A2 => n12782, B1 => n12781, B2 
                           => n12771, ZN => N2534);
   U1811 : AOI22_X1 port map( A1 => DATA2(16), A2 => n12782, B1 => n12781, B2 
                           => n12772, ZN => N2533);
   U1812 : AOI22_X1 port map( A1 => DATA2(15), A2 => n12782, B1 => n12781, B2 
                           => n12773, ZN => N2532);
   U1813 : AOI22_X1 port map( A1 => DATA2(14), A2 => n12782, B1 => n12781, B2 
                           => n12774, ZN => N2531);
   U1814 : AOI22_X1 port map( A1 => DATA2(13), A2 => n12782, B1 => n12781, B2 
                           => n12775, ZN => N2530);
   U1815 : AOI22_X1 port map( A1 => DATA2(12), A2 => n12782, B1 => n12781, B2 
                           => n12776, ZN => N2529);
   U1816 : AOI22_X1 port map( A1 => DATA2(11), A2 => n12782, B1 => n12781, B2 
                           => n12777, ZN => N2528);
   U1817 : AOI22_X1 port map( A1 => DATA2(10), A2 => n12782, B1 => n12781, B2 
                           => n12778, ZN => N2527);
   U1818 : AOI22_X1 port map( A1 => DATA2(9), A2 => n12782, B1 => n12781, B2 =>
                           n12779, ZN => N2526);
   U1819 : AOI22_X1 port map( A1 => DATA2(8), A2 => n12782, B1 => n12781, B2 =>
                           n12780, ZN => N2525);
   U1820 : AOI22_X1 port map( A1 => DATA2(7), A2 => n12787, B1 => n12786, B2 =>
                           n12783, ZN => N2524);
   U1821 : AOI22_X1 port map( A1 => DATA2(6), A2 => n12787, B1 => n12786, B2 =>
                           n12784, ZN => N2523);
   U1822 : AOI22_X1 port map( A1 => DATA2(5), A2 => n12787, B1 => n12786, B2 =>
                           n12785, ZN => N2522);
   U1823 : AOI22_X1 port map( A1 => DATA2(4), A2 => n12787, B1 => n12786, B2 =>
                           n13076, ZN => N2521);
   U1824 : AOI22_X1 port map( A1 => DATA2(3), A2 => n12787, B1 => n12786, B2 =>
                           n13078, ZN => N2520);
   U1825 : AOI22_X1 port map( A1 => DATA2(2), A2 => n12787, B1 => n12786, B2 =>
                           n13077, ZN => N2519);
   U1826 : AOI22_X1 port map( A1 => DATA2(1), A2 => n12787, B1 => n12786, B2 =>
                           n13088, ZN => N2518);
   U1827 : AOI22_X1 port map( A1 => DATA2(0), A2 => n12787, B1 => n12786, B2 =>
                           n13082, ZN => N2517);
   U1828 : NOR2_X1 port map( A1 => n12788, A2 => n1826, ZN => n4192);
   U1829 : NAND2_X1 port map( A1 => n12827, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, ZN 
                           => n12792);
   U1830 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , ZN => n12823);
   U1831 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n12823, ZN => n12822);
   U1832 : INV_X1 port map( A => n12789, ZN => n12790);
   U1833 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n12825, B1 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B2 => 
                           n12819, ZN => n12791);
   U1834 : OAI221_X1 port map( B1 => n1826, B2 => n12792, C1 => n1826, C2 => 
                           n12822, A => n12791, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1835 : INV_X1 port map( A => n12792, ZN => n12824);
   U1836 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n12825, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n12824, ZN => n12794);
   U1837 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_63_port, A2
                           => n12819, ZN => n12793);
   U1838 : OAI211_X1 port map( C1 => n1825, C2 => n12822, A => n12794, B => 
                           n12793, ZN => boothmul_pipelined_i_mux_out_1_4_port)
                           ;
   U1839 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n12824, B1 => n12825, B2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n12796);
   U1840 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, ZN => 
                           n12795);
   U1841 : OAI211_X1 port map( C1 => n12822, C2 => n1824, A => n12796, B => 
                           n12795, ZN => boothmul_pipelined_i_mux_out_1_5_port)
                           ;
   U1842 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n12798);
   U1843 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, ZN => 
                           n12797);
   U1844 : OAI211_X1 port map( C1 => n1823, C2 => n12822, A => n12798, B => 
                           n12797, ZN => boothmul_pipelined_i_mux_out_1_6_port)
                           ;
   U1845 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n12800);
   U1846 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, ZN => 
                           n12799);
   U1847 : OAI211_X1 port map( C1 => n1822, C2 => n12822, A => n12800, B => 
                           n12799, ZN => boothmul_pipelined_i_mux_out_1_7_port)
                           ;
   U1848 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n12802);
   U1849 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, ZN => 
                           n12801);
   U1850 : OAI211_X1 port map( C1 => n1820, C2 => n12822, A => n12802, B => 
                           n12801, ZN => boothmul_pipelined_i_mux_out_1_8_port)
                           ;
   U1851 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n12804);
   U1852 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_34_port, ZN => 
                           n12803);
   U1853 : OAI211_X1 port map( C1 => n1819, C2 => n12822, A => n12804, B => 
                           n12803, ZN => boothmul_pipelined_i_mux_out_1_9_port)
                           ;
   U1854 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n12806);
   U1855 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_33_port, ZN => 
                           n12805);
   U1856 : OAI211_X1 port map( C1 => n1818, C2 => n12822, A => n12806, B => 
                           n12805, ZN => boothmul_pipelined_i_mux_out_1_10_port
                           );
   U1857 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n12808);
   U1858 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_32_port, ZN => 
                           n12807);
   U1859 : OAI211_X1 port map( C1 => n1817, C2 => n12822, A => n12808, B => 
                           n12807, ZN => boothmul_pipelined_i_mux_out_1_11_port
                           );
   U1860 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n12810);
   U1861 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_31_port, ZN => 
                           n12809);
   U1862 : OAI211_X1 port map( C1 => n1816, C2 => n12822, A => n12810, B => 
                           n12809, ZN => boothmul_pipelined_i_mux_out_1_12_port
                           );
   U1863 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n12812);
   U1864 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_30_port, ZN => 
                           n12811);
   U1865 : OAI211_X1 port map( C1 => n1815, C2 => n12822, A => n12812, B => 
                           n12811, ZN => boothmul_pipelined_i_mux_out_1_13_port
                           );
   U1866 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n12814);
   U1867 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_29_port, ZN => 
                           n12813);
   U1868 : OAI211_X1 port map( C1 => n1814, C2 => n12822, A => n12814, B => 
                           n12813, ZN => boothmul_pipelined_i_mux_out_1_14_port
                           );
   U1869 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n12816);
   U1870 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_28_port, ZN => 
                           n12815);
   U1871 : OAI211_X1 port map( C1 => n1813, C2 => n12822, A => n12816, B => 
                           n12815, ZN => boothmul_pipelined_i_mux_out_1_15_port
                           );
   U1872 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n12818);
   U1873 : NAND2_X1 port map( A1 => n12819, A2 => 
                           boothmul_pipelined_i_muxes_in_4_27_port, ZN => 
                           n12817);
   U1874 : OAI211_X1 port map( C1 => n1812, C2 => n12822, A => n12818, B => 
                           n12817, ZN => boothmul_pipelined_i_mux_out_1_16_port
                           );
   U1875 : AOI22_X1 port map( A1 => n12825, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n12821);
   U1876 : NAND2_X1 port map( A1 => n12819, A2 => data1_mul_15_port, ZN => 
                           n12820);
   U1877 : OAI211_X1 port map( C1 => n1811, C2 => n12822, A => n12821, B => 
                           n12820, ZN => boothmul_pipelined_i_mux_out_1_17_port
                           );
   U1878 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n12823, ZN => 
                           n12828);
   U1879 : AOI22_X1 port map( A1 => n12825, A2 => n1809, B1 => n12824, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n12826);
   U1880 : OAI21_X1 port map( B1 => n12828, B2 => n12827, A => n12826, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1881 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           ZN => n13084);
   U1882 : OR2_X1 port map( A1 => n13084, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n4055);
   U1883 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n9093, B1 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B2 => n8887
                           , ZN => n12829);
   U1884 : OAI221_X1 port map( B1 => n1826, B2 => n9116, C1 => n1826, C2 => 
                           n8932, A => n12829, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1885 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n8803, B1 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B2 => n8887
                           , ZN => n12831);
   U1886 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n9093, ZN => n12830);
   U1887 : OAI211_X1 port map( C1 => n8932, C2 => n1825, A => n12831, B => 
                           n12830, ZN => boothmul_pipelined_i_mux_out_2_6_port)
                           ;
   U1888 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_62_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n9093, ZN => n12833);
   U1889 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n8803, ZN => n12832);
   U1890 : OAI211_X1 port map( C1 => n8932, C2 => n1824, A => n12833, B => 
                           n12832, ZN => boothmul_pipelined_i_mux_out_2_7_port)
                           ;
   U1891 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_61_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n9093, ZN => n12835);
   U1892 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n8803, ZN => n12834);
   U1893 : OAI211_X1 port map( C1 => n8932, C2 => n1823, A => n12835, B => 
                           n12834, ZN => boothmul_pipelined_i_mux_out_2_8_port)
                           ;
   U1894 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_60_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n9093, ZN => n12837);
   U1895 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n8803, ZN => n12836);
   U1896 : OAI211_X1 port map( C1 => n8932, C2 => n1822, A => n12837, B => 
                           n12836, ZN => boothmul_pipelined_i_mux_out_2_9_port)
                           ;
   U1897 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_59_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n9093, ZN => n12839);
   U1898 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n8803, ZN => n12838);
   U1899 : OAI211_X1 port map( C1 => n8932, C2 => n1820, A => n12839, B => 
                           n12838, ZN => boothmul_pipelined_i_mux_out_2_10_port
                           );
   U1900 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_34_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n9093, ZN => n12841);
   U1901 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n8803, ZN => n12840);
   U1902 : OAI211_X1 port map( C1 => n8932, C2 => n1819, A => n12841, B => 
                           n12840, ZN => boothmul_pipelined_i_mux_out_2_11_port
                           );
   U1903 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_33_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n9093, ZN => n12843);
   U1904 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n8803, ZN => n12842);
   U1905 : OAI211_X1 port map( C1 => n8932, C2 => n1818, A => n12843, B => 
                           n12842, ZN => boothmul_pipelined_i_mux_out_2_12_port
                           );
   U1906 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_32_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n9093, ZN => n12845);
   U1907 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n8803, ZN => n12844);
   U1908 : OAI211_X1 port map( C1 => n8932, C2 => n1817, A => n12845, B => 
                           n12844, ZN => boothmul_pipelined_i_mux_out_2_13_port
                           );
   U1909 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_31_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n9093, ZN => n12847);
   U1910 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n8803, ZN => n12846);
   U1911 : OAI211_X1 port map( C1 => n8932, C2 => n1816, A => n12847, B => 
                           n12846, ZN => boothmul_pipelined_i_mux_out_2_14_port
                           );
   U1912 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_30_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n9093, ZN => n12849);
   U1913 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n8803, ZN => n12848);
   U1914 : OAI211_X1 port map( C1 => n8932, C2 => n1815, A => n12849, B => 
                           n12848, ZN => boothmul_pipelined_i_mux_out_2_15_port
                           );
   U1915 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_29_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n9093, ZN => n12851);
   U1916 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n8803, ZN => n12850);
   U1917 : OAI211_X1 port map( C1 => n8932, C2 => n1814, A => n12851, B => 
                           n12850, ZN => boothmul_pipelined_i_mux_out_2_16_port
                           );
   U1918 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_28_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n9093, ZN => n12853);
   U1919 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n8803, ZN => n12852);
   U1920 : OAI211_X1 port map( C1 => n8932, C2 => n1813, A => n12853, B => 
                           n12852, ZN => boothmul_pipelined_i_mux_out_2_17_port
                           );
   U1921 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_27_port, A2
                           => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n9093, ZN => n12855);
   U1922 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n8803, ZN => n12854);
   U1923 : OAI211_X1 port map( C1 => n8932, C2 => n1812, A => n12855, B => 
                           n12854, ZN => boothmul_pipelined_i_mux_out_2_18_port
                           );
   U1924 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n8887, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n9093, ZN => n12857);
   U1925 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n8803, ZN => n12856);
   U1926 : OAI211_X1 port map( C1 => n8932, C2 => n1811, A => n12857, B => 
                           n12856, ZN => boothmul_pipelined_i_mux_out_2_19_port
                           );
   U1927 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_102_port, ZN 
                           => n12889);
   U1928 : INV_X1 port map( A => n1809, ZN => n12888);
   U1929 : OAI222_X1 port map( A1 => n12889, A2 => n9116, B1 => n1810, B2 => 
                           n8888, C1 => n8976, C2 => n12888, ZN => n3800);
   U1930 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n4295, ZN => n12858);
   U1931 : NAND2_X1 port map( A1 => n12858, A2 => n7769, ZN => n7485);
   U1932 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n8977, B1 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B2 => n8930
                           , ZN => n12859);
   U1933 : OAI221_X1 port map( B1 => n1826, B2 => n8931, C1 => n1826, C2 => 
                           n8814, A => n12859, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1934 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_116_port, ZN 
                           => n13046);
   U1935 : OAI22_X1 port map( A1 => n8931, A2 => n13046, B1 => n8814, B2 => 
                           n1825, ZN => n12860);
   U1936 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           B2 => n8977, A => n12860, ZN => n12861);
   U1937 : OAI21_X1 port map( B1 => n9189, B2 => n1824, A => n12861, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1938 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_115_port, ZN 
                           => n13047);
   U1939 : OAI22_X1 port map( A1 => n8814, A2 => n1824, B1 => n9189, B2 => 
                           n1823, ZN => n12862);
   U1940 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           B2 => n8977, A => n12862, ZN => n12863);
   U1941 : OAI21_X1 port map( B1 => n8931, B2 => n13047, A => n12863, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1942 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_114_port, ZN 
                           => n13048);
   U1943 : OAI22_X1 port map( A1 => n8931, A2 => n13048, B1 => n9189, B2 => 
                           n1822, ZN => n12864);
   U1944 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           B2 => n8977, A => n12864, ZN => n12865);
   U1945 : OAI21_X1 port map( B1 => n8814, B2 => n1823, A => n12865, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1946 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_113_port, ZN 
                           => n13049);
   U1947 : OAI22_X1 port map( A1 => n8931, A2 => n13049, B1 => n9189, B2 => 
                           n1820, ZN => n12866);
   U1948 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           B2 => n8977, A => n12866, ZN => n12867);
   U1949 : OAI21_X1 port map( B1 => n8814, B2 => n1822, A => n12867, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1950 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_112_port, ZN 
                           => n13050);
   U1951 : OAI22_X1 port map( A1 => n8931, A2 => n13050, B1 => n9189, B2 => 
                           n1819, ZN => n12868);
   U1952 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           B2 => n8977, A => n12868, ZN => n12869);
   U1953 : OAI21_X1 port map( B1 => n8814, B2 => n1820, A => n12869, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1954 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_111_port, ZN 
                           => n13051);
   U1955 : OAI22_X1 port map( A1 => n8931, A2 => n13051, B1 => n9189, B2 => 
                           n1818, ZN => n12870);
   U1956 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           B2 => n8977, A => n12870, ZN => n12871);
   U1957 : OAI21_X1 port map( B1 => n8814, B2 => n1819, A => n12871, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U1958 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_110_port, ZN 
                           => n13052);
   U1959 : OAI22_X1 port map( A1 => n8931, A2 => n13052, B1 => n9189, B2 => 
                           n1817, ZN => n12872);
   U1960 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           B2 => n8977, A => n12872, ZN => n12873);
   U1961 : OAI21_X1 port map( B1 => n8814, B2 => n1818, A => n12873, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U1962 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_109_port, ZN 
                           => n13053);
   U1963 : OAI22_X1 port map( A1 => n8931, A2 => n13053, B1 => n9189, B2 => 
                           n1816, ZN => n12874);
   U1964 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           B2 => n8977, A => n12874, ZN => n12875);
   U1965 : OAI21_X1 port map( B1 => n8814, B2 => n1817, A => n12875, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U1966 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_108_port, ZN 
                           => n13054);
   U1967 : OAI22_X1 port map( A1 => n8931, A2 => n13054, B1 => n9189, B2 => 
                           n1815, ZN => n12876);
   U1968 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           B2 => n8977, A => n12876, ZN => n12877);
   U1969 : OAI21_X1 port map( B1 => n8814, B2 => n1816, A => n12877, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U1970 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_107_port, ZN 
                           => n13055);
   U1971 : OAI22_X1 port map( A1 => n8931, A2 => n13055, B1 => n9189, B2 => 
                           n1814, ZN => n12878);
   U1972 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           B2 => n8977, A => n12878, ZN => n12879);
   U1973 : OAI21_X1 port map( B1 => n8814, B2 => n1815, A => n12879, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U1974 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_106_port, ZN 
                           => n13056);
   U1975 : OAI22_X1 port map( A1 => n8931, A2 => n13056, B1 => n9189, B2 => 
                           n1813, ZN => n12880);
   U1976 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           B2 => n8977, A => n12880, ZN => n12881);
   U1977 : OAI21_X1 port map( B1 => n8814, B2 => n1814, A => n12881, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U1978 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_105_port, ZN 
                           => n13057);
   U1979 : OAI22_X1 port map( A1 => n8931, A2 => n13057, B1 => n9189, B2 => 
                           n1812, ZN => n12882);
   U1980 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           B2 => n8977, A => n12882, ZN => n12883);
   U1981 : OAI21_X1 port map( B1 => n8814, B2 => n1813, A => n12883, ZN => 
                           n4190);
   U1982 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_104_port, ZN 
                           => n13059);
   U1983 : OAI22_X1 port map( A1 => n8931, A2 => n13059, B1 => n9189, B2 => 
                           n1811, ZN => n12884);
   U1984 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           B2 => n8977, A => n12884, ZN => n12885);
   U1985 : OAI21_X1 port map( B1 => n8814, B2 => n1812, A => n12885, ZN => 
                           n4189);
   U1986 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_103_port, ZN 
                           => n13061);
   U1987 : OAI22_X1 port map( A1 => n8931, A2 => n13061, B1 => n9189, B2 => 
                           n1810, ZN => n12886);
   U1988 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           B2 => n8977, A => n12886, ZN => n12887);
   U1989 : OAI21_X1 port map( B1 => n8814, B2 => n1811, A => n12887, ZN => 
                           n4188);
   U1990 : OAI222_X1 port map( A1 => n12889, A2 => n8931, B1 => n1810, B2 => 
                           n8929, C1 => n9188, C2 => n12888, ZN => n4187);
   U1991 : NAND3_X1 port map( A1 => n11328, A2 => n8978, A3 => n11306, ZN => 
                           n12927);
   U1992 : OR2_X1 port map( A1 => n8978, A2 => n11306, ZN => n12890);
   U1993 : INV_X1 port map( A => n12925, ZN => n12894);
   U1994 : NAND2_X1 port map( A1 => n11328, A2 => n12892, ZN => n12928);
   U1995 : INV_X1 port map( A => n12928, ZN => n12921);
   U1996 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n12924, B1 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B2 => 
                           n12921, ZN => n12893);
   U1997 : OAI221_X1 port map( B1 => n1826, B2 => n12927, C1 => n1826, C2 => 
                           n12894, A => n12893, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U1998 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n12924, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n12925, ZN => n12896);
   U1999 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_63_port, A2
                           => n12921, ZN => n12895);
   U2000 : OAI211_X1 port map( C1 => n12927, C2 => n1825, A => n12896, B => 
                           n12895, ZN => boothmul_pipelined_i_mux_out_4_10_port
                           );
   U2001 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n12924, ZN => n12898);
   U2002 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_62_port, A2
                           => n12921, ZN => n12897);
   U2003 : OAI211_X1 port map( C1 => n12927, C2 => n1824, A => n12898, B => 
                           n12897, ZN => boothmul_pipelined_i_mux_out_4_11_port
                           );
   U2004 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n12924, ZN => n12900);
   U2005 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_61_port, A2
                           => n12921, ZN => n12899);
   U2006 : OAI211_X1 port map( C1 => n12927, C2 => n1823, A => n12900, B => 
                           n12899, ZN => boothmul_pipelined_i_mux_out_4_12_port
                           );
   U2007 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n12924, ZN => n12902);
   U2008 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_60_port, A2
                           => n12921, ZN => n12901);
   U2009 : OAI211_X1 port map( C1 => n12927, C2 => n1822, A => n12902, B => 
                           n12901, ZN => boothmul_pipelined_i_mux_out_4_13_port
                           );
   U2010 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n12924, ZN => n12904);
   U2011 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_59_port, A2
                           => n12921, ZN => n12903);
   U2012 : OAI211_X1 port map( C1 => n12927, C2 => n1820, A => n12904, B => 
                           n12903, ZN => boothmul_pipelined_i_mux_out_4_14_port
                           );
   U2013 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n12924, ZN => n12906);
   U2014 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_34_port, A2
                           => n12921, ZN => n12905);
   U2015 : OAI211_X1 port map( C1 => n12927, C2 => n1819, A => n12906, B => 
                           n12905, ZN => boothmul_pipelined_i_mux_out_4_15_port
                           );
   U2016 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n12924, ZN => n12908);
   U2017 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_33_port, A2
                           => n12921, ZN => n12907);
   U2018 : OAI211_X1 port map( C1 => n12927, C2 => n1818, A => n12908, B => 
                           n12907, ZN => boothmul_pipelined_i_mux_out_4_16_port
                           );
   U2019 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n12924, ZN => n12910);
   U2020 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_32_port, A2
                           => n12921, ZN => n12909);
   U2021 : OAI211_X1 port map( C1 => n12927, C2 => n1817, A => n12910, B => 
                           n12909, ZN => boothmul_pipelined_i_mux_out_4_17_port
                           );
   U2022 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n12924, ZN => n12912);
   U2023 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_31_port, A2
                           => n12921, ZN => n12911);
   U2024 : OAI211_X1 port map( C1 => n12927, C2 => n1816, A => n12912, B => 
                           n12911, ZN => boothmul_pipelined_i_mux_out_4_18_port
                           );
   U2025 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n12924, ZN => n12914);
   U2026 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_30_port, A2
                           => n12921, ZN => n12913);
   U2027 : OAI211_X1 port map( C1 => n12927, C2 => n1815, A => n12914, B => 
                           n12913, ZN => boothmul_pipelined_i_mux_out_4_19_port
                           );
   U2028 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n12924, ZN => n12916);
   U2029 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_29_port, A2
                           => n12921, ZN => n12915);
   U2030 : OAI211_X1 port map( C1 => n12927, C2 => n1814, A => n12916, B => 
                           n12915, ZN => boothmul_pipelined_i_mux_out_4_20_port
                           );
   U2031 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n12924, ZN => n12918);
   U2032 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_28_port, A2
                           => n12921, ZN => n12917);
   U2033 : OAI211_X1 port map( C1 => n12927, C2 => n1813, A => n12918, B => 
                           n12917, ZN => boothmul_pipelined_i_mux_out_4_21_port
                           );
   U2034 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n12924, ZN => n12920);
   U2035 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_27_port, A2
                           => n12921, ZN => n12919);
   U2036 : OAI211_X1 port map( C1 => n12927, C2 => n1812, A => n12920, B => 
                           n12919, ZN => n4186);
   U2037 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n12925, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n12924, ZN => n12923);
   U2038 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n12921, ZN => 
                           n12922);
   U2039 : OAI211_X1 port map( C1 => n12927, C2 => n1811, A => n12923, B => 
                           n12922, ZN => n4185);
   U2040 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n12925, B1 => n12924, B2 => n1809, ZN => 
                           n12926);
   U2041 : OAI221_X1 port map( B1 => n1810, B2 => n12928, C1 => n1810, C2 => 
                           n12927, A => n12926, ZN => n4184);
   U2042 : NAND3_X1 port map( A1 => n11326, A2 => n8980, A3 => n11307, ZN => 
                           n12966);
   U2043 : NOR2_X1 port map( A1 => n8980, A2 => n11307, ZN => n12929);
   U2044 : NAND2_X1 port map( A1 => n12929, A2 => n13174, ZN => n12932);
   U2045 : AOI22_X1 port map( A1 => n12959, A2 => n9085, B1 => n12963, B2 => 
                           n9119, ZN => n12931);
   U2046 : OAI221_X1 port map( B1 => n11310, B2 => n12966, C1 => n11310, C2 => 
                           n12932, A => n12931, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2047 : INV_X1 port map( A => n12966, ZN => n12960);
   U2048 : INV_X1 port map( A => n12932, ZN => n12964);
   U2049 : AOI22_X1 port map( A1 => n9085, A2 => n12960, B1 => n12964, B2 => 
                           n9119, ZN => n12934);
   U2050 : AOI22_X1 port map( A1 => n12959, A2 => n9082, B1 => n12963, B2 => 
                           n9122, ZN => n12933);
   U2051 : NAND2_X1 port map( A1 => n12934, A2 => n12933, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2052 : AOI22_X1 port map( A1 => n12960, A2 => n9082, B1 => n12964, B2 => 
                           n9122, ZN => n12936);
   U2053 : AOI22_X1 port map( A1 => n12959, A2 => n9079, B1 => n12963, B2 => 
                           n9125, ZN => n12935);
   U2054 : NAND2_X1 port map( A1 => n12936, A2 => n12935, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2055 : AOI22_X1 port map( A1 => n12960, A2 => n9079, B1 => n12964, B2 => 
                           n9125, ZN => n12938);
   U2056 : AOI22_X1 port map( A1 => n12959, A2 => n9076, B1 => n12963, B2 => 
                           n9128, ZN => n12937);
   U2057 : NAND2_X1 port map( A1 => n12938, A2 => n12937, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2058 : AOI22_X1 port map( A1 => n12960, A2 => n9076, B1 => n12964, B2 => 
                           n9128, ZN => n12940);
   U2059 : AOI22_X1 port map( A1 => n12959, A2 => n9073, B1 => n12963, B2 => 
                           n9131, ZN => n12939);
   U2060 : NAND2_X1 port map( A1 => n12940, A2 => n12939, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2061 : AOI22_X1 port map( A1 => n12960, A2 => n9073, B1 => n12964, B2 => 
                           n9131, ZN => n12942);
   U2062 : AOI22_X1 port map( A1 => n12959, A2 => n9070, B1 => n12963, B2 => 
                           n9134, ZN => n12941);
   U2063 : NAND2_X1 port map( A1 => n12942, A2 => n12941, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2064 : AOI22_X1 port map( A1 => n12960, A2 => n9070, B1 => n12964, B2 => 
                           n9134, ZN => n12944);
   U2065 : AOI22_X1 port map( A1 => n12959, A2 => n9067, B1 => n12963, B2 => 
                           n9137, ZN => n12943);
   U2066 : NAND2_X1 port map( A1 => n12944, A2 => n12943, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2067 : AOI22_X1 port map( A1 => n12960, A2 => n9067, B1 => n12964, B2 => 
                           n9137, ZN => n12946);
   U2068 : AOI22_X1 port map( A1 => n12959, A2 => n9064, B1 => n12963, B2 => 
                           n9140, ZN => n12945);
   U2069 : NAND2_X1 port map( A1 => n12946, A2 => n12945, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2070 : AOI22_X1 port map( A1 => n12960, A2 => n9064, B1 => n12964, B2 => 
                           n9140, ZN => n12948);
   U2071 : AOI22_X1 port map( A1 => n12959, A2 => n9061, B1 => n12963, B2 => 
                           n9143, ZN => n12947);
   U2072 : NAND2_X1 port map( A1 => n12948, A2 => n12947, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2073 : AOI22_X1 port map( A1 => n12960, A2 => n9061, B1 => n12964, B2 => 
                           n9143, ZN => n12950);
   U2074 : AOI22_X1 port map( A1 => n12959, A2 => n9058, B1 => n12963, B2 => 
                           n9146, ZN => n12949);
   U2075 : NAND2_X1 port map( A1 => n12950, A2 => n12949, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2076 : AOI22_X1 port map( A1 => n12960, A2 => n9058, B1 => n12964, B2 => 
                           n9146, ZN => n12952);
   U2077 : AOI22_X1 port map( A1 => n12959, A2 => n9055, B1 => n12963, B2 => 
                           n9149, ZN => n12951);
   U2078 : NAND2_X1 port map( A1 => n12952, A2 => n12951, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2079 : AOI22_X1 port map( A1 => n12960, A2 => n9055, B1 => n12964, B2 => 
                           n9149, ZN => n12954);
   U2080 : AOI22_X1 port map( A1 => n12959, A2 => n9052, B1 => n12963, B2 => 
                           n9152, ZN => n12953);
   U2081 : NAND2_X1 port map( A1 => n12954, A2 => n12953, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2082 : AOI22_X1 port map( A1 => n12960, A2 => n9052, B1 => n12964, B2 => 
                           n9152, ZN => n12956);
   U2083 : AOI22_X1 port map( A1 => n12959, A2 => n9049, B1 => n12963, B2 => 
                           n9155, ZN => n12955);
   U2084 : NAND2_X1 port map( A1 => n12956, A2 => n12955, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2085 : AOI22_X1 port map( A1 => n12960, A2 => n9049, B1 => n12964, B2 => 
                           n9155, ZN => n12958);
   U2086 : AOI22_X1 port map( A1 => n12959, A2 => n9046, B1 => n12963, B2 => 
                           n9158, ZN => n12957);
   U2087 : NAND2_X1 port map( A1 => n12958, A2 => n12957, ZN => n4183);
   U2088 : INV_X1 port map( A => n12959, ZN => n12967);
   U2089 : AOI22_X1 port map( A1 => n12960, A2 => n9046, B1 => n12964, B2 => 
                           n9158, ZN => n12962);
   U2090 : NAND2_X1 port map( A1 => n12963, A2 => n9161, ZN => n12961);
   U2091 : OAI211_X1 port map( C1 => n11302, C2 => n12967, A => n12962, B => 
                           n12961, ZN => n4182);
   U2092 : AOI22_X1 port map( A1 => n12964, A2 => n9161, B1 => n12963, B2 => 
                           n9097, ZN => n12965);
   U2093 : OAI221_X1 port map( B1 => n11302, B2 => n12967, C1 => n11302, C2 => 
                           n12966, A => n12965, ZN => n4181);
   U2094 : NAND3_X1 port map( A1 => n11329, A2 => n8984, A3 => n11308, ZN => 
                           n13005);
   U2095 : NOR2_X1 port map( A1 => n8984, A2 => n11308, ZN => n12968);
   U2096 : NAND2_X1 port map( A1 => n12968, A2 => n13175, ZN => n12971);
   U2097 : AOI22_X1 port map( A1 => n12998, A2 => n9084, B1 => n13002, B2 => 
                           n9118, ZN => n12970);
   U2098 : OAI221_X1 port map( B1 => n11300, B2 => n13005, C1 => n11300, C2 => 
                           n12971, A => n12970, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2099 : INV_X1 port map( A => n13005, ZN => n12999);
   U2100 : INV_X1 port map( A => n12971, ZN => n13003);
   U2101 : AOI22_X1 port map( A1 => n9084, A2 => n12999, B1 => n13003, B2 => 
                           n9118, ZN => n12973);
   U2102 : AOI22_X1 port map( A1 => n12998, A2 => n9081, B1 => n13002, B2 => 
                           n9121, ZN => n12972);
   U2103 : NAND2_X1 port map( A1 => n12973, A2 => n12972, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2104 : AOI22_X1 port map( A1 => n12999, A2 => n9081, B1 => n13003, B2 => 
                           n9121, ZN => n12975);
   U2105 : AOI22_X1 port map( A1 => n12998, A2 => n9078, B1 => n13002, B2 => 
                           n9124, ZN => n12974);
   U2106 : NAND2_X1 port map( A1 => n12975, A2 => n12974, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2107 : AOI22_X1 port map( A1 => n12999, A2 => n9078, B1 => n13003, B2 => 
                           n9124, ZN => n12977);
   U2108 : AOI22_X1 port map( A1 => n12998, A2 => n9075, B1 => n13002, B2 => 
                           n9127, ZN => n12976);
   U2109 : NAND2_X1 port map( A1 => n12977, A2 => n12976, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2110 : AOI22_X1 port map( A1 => n12999, A2 => n9075, B1 => n13003, B2 => 
                           n9127, ZN => n12979);
   U2111 : AOI22_X1 port map( A1 => n12998, A2 => n9072, B1 => n13002, B2 => 
                           n9130, ZN => n12978);
   U2112 : NAND2_X1 port map( A1 => n12979, A2 => n12978, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2113 : AOI22_X1 port map( A1 => n12999, A2 => n9072, B1 => n13003, B2 => 
                           n9130, ZN => n12981);
   U2114 : AOI22_X1 port map( A1 => n12998, A2 => n9069, B1 => n13002, B2 => 
                           n9133, ZN => n12980);
   U2115 : NAND2_X1 port map( A1 => n12981, A2 => n12980, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2116 : AOI22_X1 port map( A1 => n12999, A2 => n9069, B1 => n13003, B2 => 
                           n9133, ZN => n12983);
   U2117 : AOI22_X1 port map( A1 => n12998, A2 => n9066, B1 => n13002, B2 => 
                           n9136, ZN => n12982);
   U2118 : NAND2_X1 port map( A1 => n12983, A2 => n12982, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2119 : AOI22_X1 port map( A1 => n12999, A2 => n9066, B1 => n13003, B2 => 
                           n9136, ZN => n12985);
   U2120 : AOI22_X1 port map( A1 => n12998, A2 => n9063, B1 => n13002, B2 => 
                           n9139, ZN => n12984);
   U2121 : NAND2_X1 port map( A1 => n12985, A2 => n12984, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2122 : AOI22_X1 port map( A1 => n12999, A2 => n9063, B1 => n13003, B2 => 
                           n9139, ZN => n12987);
   U2123 : AOI22_X1 port map( A1 => n12998, A2 => n9060, B1 => n13002, B2 => 
                           n9142, ZN => n12986);
   U2124 : NAND2_X1 port map( A1 => n12987, A2 => n12986, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2125 : AOI22_X1 port map( A1 => n12999, A2 => n9060, B1 => n13003, B2 => 
                           n9142, ZN => n12989);
   U2126 : AOI22_X1 port map( A1 => n12998, A2 => n9057, B1 => n13002, B2 => 
                           n9145, ZN => n12988);
   U2127 : NAND2_X1 port map( A1 => n12989, A2 => n12988, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2128 : AOI22_X1 port map( A1 => n12999, A2 => n9057, B1 => n13003, B2 => 
                           n9145, ZN => n12991);
   U2129 : AOI22_X1 port map( A1 => n12998, A2 => n9054, B1 => n13002, B2 => 
                           n9148, ZN => n12990);
   U2130 : NAND2_X1 port map( A1 => n12991, A2 => n12990, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2131 : AOI22_X1 port map( A1 => n12999, A2 => n9054, B1 => n13003, B2 => 
                           n9148, ZN => n12993);
   U2132 : AOI22_X1 port map( A1 => n12998, A2 => n9051, B1 => n13002, B2 => 
                           n9151, ZN => n12992);
   U2133 : NAND2_X1 port map( A1 => n12993, A2 => n12992, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2134 : AOI22_X1 port map( A1 => n12999, A2 => n9051, B1 => n13003, B2 => 
                           n9151, ZN => n12995);
   U2135 : AOI22_X1 port map( A1 => n12998, A2 => n9048, B1 => n13002, B2 => 
                           n9154, ZN => n12994);
   U2136 : NAND2_X1 port map( A1 => n12995, A2 => n12994, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2137 : AOI22_X1 port map( A1 => n12999, A2 => n9048, B1 => n13003, B2 => 
                           n9154, ZN => n12997);
   U2138 : AOI22_X1 port map( A1 => n12998, A2 => n9045, B1 => n13002, B2 => 
                           n9157, ZN => n12996);
   U2139 : NAND2_X1 port map( A1 => n12997, A2 => n12996, ZN => n4180);
   U2140 : INV_X1 port map( A => n12998, ZN => n13006);
   U2141 : AOI22_X1 port map( A1 => n12999, A2 => n9045, B1 => n13003, B2 => 
                           n9157, ZN => n13001);
   U2142 : NAND2_X1 port map( A1 => n13002, A2 => n9160, ZN => n13000);
   U2143 : OAI211_X1 port map( C1 => n11303, C2 => n13006, A => n13001, B => 
                           n13000, ZN => n4179);
   U2144 : AOI22_X1 port map( A1 => n13003, A2 => n9160, B1 => n13002, B2 => 
                           n9096, ZN => n13004);
   U2145 : OAI221_X1 port map( B1 => n11303, B2 => n13006, C1 => n11303, C2 => 
                           n13005, A => n13004, ZN => n4178);
   U2146 : NAND3_X1 port map( A1 => n11325, A2 => n11309, A3 => n8990, ZN => 
                           n13010);
   U2147 : INV_X1 port map( A => n13042, ZN => n13009);
   U2148 : AOI22_X1 port map( A1 => n13040, A2 => n9083, B1 => n13041, B2 => 
                           n9117, ZN => n13008);
   U2149 : OAI221_X1 port map( B1 => n11301, B2 => n13010, C1 => n11301, C2 => 
                           n13009, A => n13008, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2150 : INV_X1 port map( A => n13010, ZN => n13039);
   U2151 : AOI22_X1 port map( A1 => n9083, A2 => n13039, B1 => n13042, B2 => 
                           n9117, ZN => n13012);
   U2152 : AOI22_X1 port map( A1 => n13040, A2 => n9080, B1 => n13041, B2 => 
                           n9120, ZN => n13011);
   U2153 : NAND2_X1 port map( A1 => n13012, A2 => n13011, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2154 : AOI22_X1 port map( A1 => n13039, A2 => n9080, B1 => n13042, B2 => 
                           n9120, ZN => n13014);
   U2155 : AOI22_X1 port map( A1 => n13040, A2 => n9077, B1 => n13041, B2 => 
                           n9123, ZN => n13013);
   U2156 : NAND2_X1 port map( A1 => n13014, A2 => n13013, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2157 : AOI22_X1 port map( A1 => n13039, A2 => n9077, B1 => n13042, B2 => 
                           n9123, ZN => n13016);
   U2158 : AOI22_X1 port map( A1 => n13040, A2 => n9074, B1 => n13041, B2 => 
                           n9126, ZN => n13015);
   U2159 : NAND2_X1 port map( A1 => n13016, A2 => n13015, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2160 : AOI22_X1 port map( A1 => n13039, A2 => n9074, B1 => n13042, B2 => 
                           n9126, ZN => n13018);
   U2161 : AOI22_X1 port map( A1 => n13040, A2 => n9071, B1 => n13041, B2 => 
                           n9129, ZN => n13017);
   U2162 : NAND2_X1 port map( A1 => n13018, A2 => n13017, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2163 : AOI22_X1 port map( A1 => n13039, A2 => n9071, B1 => n13042, B2 => 
                           n9129, ZN => n13020);
   U2164 : AOI22_X1 port map( A1 => n13040, A2 => n9068, B1 => n13041, B2 => 
                           n9132, ZN => n13019);
   U2165 : NAND2_X1 port map( A1 => n13020, A2 => n13019, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2166 : AOI22_X1 port map( A1 => n13039, A2 => n9068, B1 => n13042, B2 => 
                           n9132, ZN => n13022);
   U2167 : AOI22_X1 port map( A1 => n13040, A2 => n9065, B1 => n13041, B2 => 
                           n9135, ZN => n13021);
   U2168 : NAND2_X1 port map( A1 => n13022, A2 => n13021, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2169 : AOI22_X1 port map( A1 => n13039, A2 => n9065, B1 => n13042, B2 => 
                           n9135, ZN => n13024);
   U2170 : AOI22_X1 port map( A1 => n13040, A2 => n9062, B1 => n13041, B2 => 
                           n9138, ZN => n13023);
   U2171 : NAND2_X1 port map( A1 => n13024, A2 => n13023, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2172 : AOI22_X1 port map( A1 => n13039, A2 => n9062, B1 => n13042, B2 => 
                           n9138, ZN => n13026);
   U2173 : AOI22_X1 port map( A1 => n13040, A2 => n9059, B1 => n13041, B2 => 
                           n9141, ZN => n13025);
   U2174 : NAND2_X1 port map( A1 => n13026, A2 => n13025, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2175 : AOI22_X1 port map( A1 => n13039, A2 => n9059, B1 => n13042, B2 => 
                           n9141, ZN => n13028);
   U2176 : AOI22_X1 port map( A1 => n13040, A2 => n9056, B1 => n13041, B2 => 
                           n9144, ZN => n13027);
   U2177 : NAND2_X1 port map( A1 => n13028, A2 => n13027, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2178 : AOI22_X1 port map( A1 => n13039, A2 => n9056, B1 => n13042, B2 => 
                           n9144, ZN => n13030);
   U2179 : AOI22_X1 port map( A1 => n13040, A2 => n9053, B1 => n13041, B2 => 
                           n9147, ZN => n13029);
   U2180 : NAND2_X1 port map( A1 => n13030, A2 => n13029, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2181 : AOI22_X1 port map( A1 => n13039, A2 => n9053, B1 => n13042, B2 => 
                           n9147, ZN => n13032);
   U2182 : AOI22_X1 port map( A1 => n13040, A2 => n9050, B1 => n13041, B2 => 
                           n9150, ZN => n13031);
   U2183 : NAND2_X1 port map( A1 => n13032, A2 => n13031, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2184 : AOI22_X1 port map( A1 => n13039, A2 => n9050, B1 => n13042, B2 => 
                           n9150, ZN => n13034);
   U2185 : AOI22_X1 port map( A1 => n13040, A2 => n9047, B1 => n13041, B2 => 
                           n9153, ZN => n13033);
   U2186 : NAND2_X1 port map( A1 => n13034, A2 => n13033, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2187 : AOI22_X1 port map( A1 => n13039, A2 => n9047, B1 => n13042, B2 => 
                           n9153, ZN => n13036);
   U2188 : AOI22_X1 port map( A1 => n13040, A2 => n9044, B1 => n13041, B2 => 
                           n9156, ZN => n13035);
   U2189 : NAND2_X1 port map( A1 => n13036, A2 => n13035, ZN => n4177);
   U2190 : AOI22_X1 port map( A1 => n13039, A2 => n9044, B1 => n13042, B2 => 
                           n9156, ZN => n13038);
   U2191 : AOI22_X1 port map( A1 => n13040, A2 => n9041, B1 => n13041, B2 => 
                           n9159, ZN => n13037);
   U2192 : NAND2_X1 port map( A1 => n13038, A2 => n13037, ZN => n4176);
   U2193 : OAI21_X1 port map( B1 => n13040, B2 => n13039, A => n9041, ZN => 
                           n13044);
   U2194 : AOI22_X1 port map( A1 => n13042, A2 => n9159, B1 => n13041, B2 => 
                           n9095, ZN => n13043);
   U2195 : NAND2_X1 port map( A1 => n13044, A2 => n13043, ZN => n4175);
   U2196 : INV_X1 port map( A => n13045, ZN => n13066);
   U2197 : OAI222_X1 port map( A1 => n1826, A2 => n13058, B1 => n13046, B2 => 
                           n13060, C1 => n13066, C2 => n1825, ZN => n3794);
   U2198 : OAI222_X1 port map( A1 => n13047, A2 => n13058, B1 => n13048, B2 => 
                           n13060, C1 => n1823, C2 => n13066, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U2199 : OAI222_X1 port map( A1 => n1822, A2 => n13066, B1 => n13049, B2 => 
                           n13060, C1 => n13048, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U2200 : OAI222_X1 port map( A1 => n1820, A2 => n13066, B1 => n13050, B2 => 
                           n13060, C1 => n13049, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U2201 : OAI222_X1 port map( A1 => n1819, A2 => n13066, B1 => n13051, B2 => 
                           n13060, C1 => n13050, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U2202 : OAI222_X1 port map( A1 => n1818, A2 => n13066, B1 => n13052, B2 => 
                           n13060, C1 => n13051, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U2203 : OAI222_X1 port map( A1 => n1817, A2 => n13066, B1 => n13053, B2 => 
                           n13060, C1 => n13052, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U2204 : OAI222_X1 port map( A1 => n1816, A2 => n13066, B1 => n13054, B2 => 
                           n13060, C1 => n13053, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U2205 : OAI222_X1 port map( A1 => n1815, A2 => n13066, B1 => n13055, B2 => 
                           n13060, C1 => n13054, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U2206 : OAI222_X1 port map( A1 => n1814, A2 => n13066, B1 => n13056, B2 => 
                           n13060, C1 => n13055, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U2207 : OAI222_X1 port map( A1 => n1813, A2 => n13066, B1 => n13057, B2 => 
                           n13060, C1 => n13056, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U2208 : OAI222_X1 port map( A1 => n1812, A2 => n13066, B1 => n13059, B2 => 
                           n13060, C1 => n13057, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U2209 : OAI222_X1 port map( A1 => n1811, A2 => n13066, B1 => n13061, B2 => 
                           n13060, C1 => n13059, C2 => n13058, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U2210 : AOI22_X1 port map( A1 => n13064, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n13063, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n13062);
   U2211 : OAI21_X1 port map( B1 => n13066, B2 => n1810, A => n13062, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2212 : AOI22_X1 port map( A1 => n13064, A2 => n1809, B1 => n13063, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n13065);
   U2213 : OAI21_X1 port map( B1 => n13066, B2 => n1810, A => n13065, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U2214 : AOI21_X1 port map( B1 => n13069, B2 => n13068, A => n13067, ZN => 
                           n4216);
   U2215 : NAND2_X1 port map( A1 => n13070, A2 => n7769, ZN => n11305);
   U2216 : NAND2_X1 port map( A1 => n13092, A2 => n13086, ZN => n11311);
   U2217 : INV_X1 port map( A => n13073, ZN => n13071);
   U2218 : NAND2_X1 port map( A1 => n13072, A2 => n13071, ZN => n11312);
   U2219 : NOR2_X1 port map( A1 => DATA2(2), A2 => DATA2(1), ZN => n13097);
   U2220 : NOR2_X1 port map( A1 => n13097, A2 => n13089, ZN => n7654);
   U2221 : NOR3_X1 port map( A1 => n7654, A2 => n13089, A3 => n13082, ZN => 
                           n11313);
   U2222 : NAND2_X1 port map( A1 => n13099, A2 => n4506, ZN => n11314);
   U2223 : NAND2_X1 port map( A1 => n13081, A2 => n13086, ZN => n11316);
   U2224 : NOR3_X1 port map( A1 => DATA2(2), A2 => n13075, A3 => n13089, ZN => 
                           n11317);
   U2225 : NAND2_X1 port map( A1 => n13074, A2 => n13073, ZN => n11318);
   U2226 : NOR2_X1 port map( A1 => n13076, A2 => n13075, ZN => n13098);
   U2227 : NAND3_X1 port map( A1 => DATA2(2), A2 => n13098, A3 => n13078, ZN =>
                           n11319);
   U2228 : NAND2_X1 port map( A1 => n13077, A2 => n13078, ZN => n13093);
   U2229 : INV_X1 port map( A => n13093, ZN => n13080);
   U2230 : NAND2_X1 port map( A1 => n13098, A2 => n13080, ZN => n11320);
   U2231 : NOR2_X1 port map( A1 => n13077, A2 => n13076, ZN => n13079);
   U2232 : INV_X1 port map( A => n13079, ZN => n13094);
   U2233 : NOR4_X1 port map( A1 => DATA2(0), A2 => n13096, A3 => n13088, A4 => 
                           n13094, ZN => n11321);
   U2234 : NAND3_X1 port map( A1 => n13081, A2 => n13079, A3 => n13078, ZN => 
                           n11322);
   U2235 : NAND3_X1 port map( A1 => n13081, A2 => n13080, A3 => n1870, ZN => 
                           n11323);
   U2236 : AOI21_X1 port map( B1 => n13097, B2 => n13082, A => n13089, ZN => 
                           n11324);
   U2237 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           ZN => n13083);
   U2238 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n13083, ZN => n11330);
   U2239 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n13084, ZN => n4111);
   U2240 : NOR2_X1 port map( A1 => n13085, A2 => n4111, ZN => n11331);
   U2241 : INV_X1 port map( A => n13086, ZN => n13087);
   U2242 : NOR2_X1 port map( A1 => n13088, A2 => n13087, ZN => n1878);
   U2243 : INV_X1 port map( A => n13089, ZN => n13090);
   U2244 : OAI21_X1 port map( B1 => DATA2(2), B2 => n13091, A => n13090, ZN => 
                           n1877);
   U2245 : INV_X1 port map( A => n13092, ZN => n13095);
   U2246 : OAI21_X1 port map( B1 => n13095, B2 => n13093, A => n1870, ZN => 
                           n1876);
   U2247 : NAND2_X1 port map( A1 => n13094, A2 => n1874, ZN => n7659);
   U2248 : OAI21_X1 port map( B1 => n13096, B2 => n13095, A => n7659, ZN => 
                           n1873);
   U2249 : NOR4_X1 port map( A1 => n13099, A2 => n13098, A3 => n13097, A4 => 
                           n7659, ZN => n1871);
   U2250 : INV_X1 port map( A => n13126, ZN => n13105);
   U2251 : OAI22_X1 port map( A1 => n13108, A2 => n13102, B1 => n13101, B2 => 
                           n13100, ZN => n13104);
   U2252 : OAI22_X1 port map( A1 => n1869, A2 => n13119, B1 => n13118, B2 => 
                           n13133, ZN => n13103);
   U2253 : AOI211_X1 port map( C1 => n13123, C2 => n13105, A => n13104, B => 
                           n13103, ZN => n1858);
   U2254 : INV_X1 port map( A => n13112, ZN => n13111);
   U2255 : OAI22_X1 port map( A1 => n1869, A2 => n13106, B1 => n13113, B2 => 
                           n11315, ZN => n13110);
   U2256 : OAI22_X1 port map( A1 => n13108, A2 => n13114, B1 => n13107, B2 => 
                           n13135, ZN => n13109);
   U2257 : AOI211_X1 port map( C1 => n1872, C2 => n13111, A => n13110, B => 
                           n13109, ZN => n1857);
   U2258 : OAI22_X1 port map( A1 => n1869, A2 => n13113, B1 => n13112, B2 => 
                           n11315, ZN => n13116);
   U2259 : OAI22_X1 port map( A1 => n13128, A2 => n13138, B1 => n13114, B2 => 
                           n13135, ZN => n13115);
   U2260 : AOI211_X1 port map( C1 => n1872, C2 => n13117, A => n13116, B => 
                           n13115, ZN => n1856);
   U2261 : OAI22_X1 port map( A1 => n13133, A2 => n13119, B1 => n13138, B2 => 
                           n13118, ZN => n13120);
   U2262 : INV_X1 port map( A => n13120, ZN => n13125);
   U2263 : AOI22_X1 port map( A1 => n13123, A2 => n13122, B1 => n13121, B2 => 
                           n1853, ZN => n13124);
   U2264 : OAI211_X1 port map( C1 => n13126, C2 => n13135, A => n13125, B => 
                           n13124, ZN => n1854);
   U2265 : OAI22_X1 port map( A1 => n13128, A2 => n1869, B1 => n13127, B2 => 
                           n13133, ZN => n13132);
   U2266 : OAI22_X1 port map( A1 => n13130, A2 => n11315, B1 => n13138, B2 => 
                           n13129, ZN => n13131);
   U2267 : AOI211_X1 port map( C1 => n13221, C2 => n6561, A => n13132, B => 
                           n13131, ZN => n1850);
   U2268 : OAI22_X1 port map( A1 => n1869, A2 => n1847, B1 => n13134, B2 => 
                           n13133, ZN => n1844);
   U2269 : INV_X1 port map( A => n6198, ZN => n13136);
   U2270 : OAI22_X1 port map( A1 => n13138, A2 => n13137, B1 => n13136, B2 => 
                           n13135, ZN => n1841);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, 
      n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, 
      n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, 
      n10097, n10098, n10099, n10100, n10101, n10102, n11132, n11133, n11136, 
      n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11149, n11150, 
      n11151, n11152, n11153, n11154, n11157, n11162, n11165, n11166, n11167, 
      n11168, n11172, n11173, n11174, n11175, n11186, n11187, n11188, n11189, 
      n11190, n11191, n11225, n11226, n11227, n11228, n11229, n11230, n11231, 
      n11232, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, 
      n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, 
      n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, 
      n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, 
      n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, 
      n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, 
      n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, 
      n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, 
      n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, 
      n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, 
      n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, 
      n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, 
      n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, 
      n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, 
      n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, 
      n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, 
      n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, 
      n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, 
      n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, 
      n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, 
      n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, 
      n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, 
      n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, 
      n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, 
      n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, 
      n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, 
      n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, 
      n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, 
      n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, 
      n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, 
      n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, 
      n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, 
      n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, 
      n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, 
      n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, 
      n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, 
      n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, 
      n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, 
      n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, 
      n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, 
      n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, 
      n13837, n13838, n13839, n13840, n13841, n13843, n13845, n13847, n13849, 
      n13851, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, 
      n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, 
      n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, 
      n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, 
      n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, 
      n13897, n13898, n13899, n13901, n13902, n13903, n13904, n13905, n13906, 
      n13907, n13908, n13909, n13910, n13911, n13913, n13914, n13915, n13917, 
      n13919, n13920, n13922, n13923, n13924, n13925, n13926, n13927, n13928, 
      n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, 
      n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, 
      n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, 
      n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, 
      n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, 
      n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, 
      n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, 
      n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, 
      n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, 
      n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, 
      n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, 
      n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, 
      n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, 
      n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, 
      n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, 
      n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, 
      n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, 
      n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, 
      n14091, n14092, n14094, n14095, n14096, n14097, n14098, n14099, n14100, 
      n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, 
      n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, 
      n14119, n14120, n14121, n14123, n14124, n14126, n14128, n14130, n14132, 
      n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, 
      n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, 
      n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, 
      n14160, n14161, n14162, n14164, n14166, n14168, n14170, n14172, n14174, 
      n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, 
      n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, 
      n14193, n14194, n14196, n14197, n14198, n14199, n14200, n14201, n14202, 
      n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14211, n14212, 
      n14213, n14214, n14215, n14216, n14217, n14219, n14221, n14222, n14223, 
      n14225, n14226, n14227, n14228, n14230, n14231, n14232, n14233, n14234, 
      n14235, n14236, n14237, n14238, n14239, n14240, n14242, n14243, n14244, 
      n14245, n14246, n14248, n14249, n14250, n14251, n14252, n14254, n14255, 
      n14256, n14257, n14258, n14259, n14260, n14262, n14263, n14264, n14265, 
      n14266, n14268, n14269, n14270, n14272, n14273, n14275, n14277, n14278, 
      n14279, n14281, n14283, n14284, n14286, n14288, n14290, n14292, n14294, 
      n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, 
      n14305, n14307, n14309, n14310, n14311, n14312, n14313, n14315, n14317, 
      n14319, n14321, n14322, n14324, n14325, n14326, n14328, n14329, n14331, 
      n14333, n14335, n14336, n14338, n14339, n14340, n14341, n14342, n14343, 
      n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14354, 
      n14356, n14357, n14359, n14360, n14362, n14364, n14366, n14367, n14368, 
      n14369, n14370, n14371, n14372, n14374, n14376, n14377, n14378, n14379, 
      n14380, n14382, n14383, n14385, n14386, n14387, n14388, n14389, n14390, 
      n14391, n14392, n14393, n14394, n14396, n14397, n14398, n14399, n14401, 
      n14402, n14403, n14405, n14407, n14409, n14411, n14413, n14415, n14416, 
      n14418, n14421, n14424, n14425, n14426, n14427, n14428, n14429, n14430, 
      n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, 
      n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, 
      n14449, n14451, n14452, n14453, n14455, n14457, n14459, n14461, n14463, 
      n14465, n14467, n14469, n14471, n14473, n14475, n14477, n14480, n14481, 
      n14482, n14483, n14485, n14486, n14487, n14489, n14491, n14492, n14494, 
      n14495, n14496, n14497, n14498, n14500, n14501, n14503, n14504, n14506, 
      n14507, n14509, n14512, n14514, n14517, n14518, n14519, n14520, n14521, 
      n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, 
      n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, 
      n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, 
      n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, 
      n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, 
      n14567, n14568, n14569, n14570, n14571, n14572, n14574, n14575, n14576, 
      n14577, n14578, n14579, n14581, n14582, n14584, n14585, n14586, n14587, 
      n14589, n14590, n14592, n14593, n14595, n14596, n14598, n14600, n14602, 
      n14605, n14607, n14609, n14611, n14613, n14615, n14617, n14620, n14632, 
      n14633, n14634, n14635, n14636, n14637, n14638, n14640, n18281, n18282, 
      n18283, n18284, n18288, n18290, n18291, n18292, n18293, n18294, n18295, 
      n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, 
      n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, 
      n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, 
      n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, 
      n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, 
      n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, 
      n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, 
      n18359, n18360, n18363, n18364, n18367, n18368, n18369, n18370, n18371, 
      n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, 
      n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, 
      n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, 
      n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, 
      n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, 
      n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, 
      n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, 
      n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, 
      n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, 
      n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, 
      n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, 
      n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, 
      n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, 
      n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, 
      n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, 
      n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, 
      n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, 
      n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, 
      n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, 
      n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, 
      n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, 
      n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, 
      n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, 
      n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, 
      n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, 
      n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, 
      n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, 
      n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, 
      n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, 
      n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, 
      n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, 
      n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, 
      n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, 
      n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, 
      n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, 
      n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, 
      n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, 
      n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, 
      n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, 
      n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, 
      n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, 
      n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, 
      n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, 
      n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, 
      n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, 
      n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, 
      n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, 
      n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, 
      n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, 
      n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, 
      n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, 
      n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, 
      n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, 
      n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, 
      n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, 
      n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, 
      n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, 
      n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, 
      n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, 
      n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, 
      n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, 
      n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, 
      n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, 
      n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, 
      n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, 
      n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, 
      n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, 
      n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, 
      n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, 
      n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, 
      n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, 
      n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, 
      n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, 
      n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, 
      n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, 
      n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, 
      n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, 
      n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, 
      n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, 
      n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, 
      n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, 
      n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, 
      n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, 
      n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, 
      n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, 
      n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, 
      n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, 
      n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, 
      n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, 
      n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, 
      n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, 
      n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, 
      n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, 
      n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, 
      n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, 
      n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, 
      n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, 
      n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, 
      n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, 
      n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, 
      n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, 
      n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, 
      n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, 
      n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, 
      n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, 
      n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, 
      n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, 
      n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, 
      n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, 
      n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, 
      n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, 
      n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, 
      n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, 
      n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, 
      n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, 
      n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, 
      n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, 
      n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, 
      n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, 
      n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, 
      n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, 
      n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, 
      n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, 
      n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, 
      n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, 
      n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, 
      n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, 
      n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, 
      n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, 
      n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, 
      n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, 
      n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, 
      n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, 
      n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, 
      n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, 
      n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, 
      n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, 
      n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, 
      n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, 
      n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, 
      n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, 
      n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, 
      n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, 
      n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, 
      n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, 
      n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, 
      n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, 
      n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, 
      n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, 
      n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, 
      n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, 
      n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, 
      n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, 
      n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, 
      n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, 
      n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, 
      n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, 
      n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, 
      n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, 
      n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, 
      n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, 
      n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, 
      n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, 
      n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, 
      n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, 
      n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, 
      n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, 
      n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, 
      n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, 
      n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, 
      n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, 
      n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, 
      n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, 
      n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, 
      n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, 
      n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, 
      n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, 
      n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, 
      n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, 
      n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, 
      n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, 
      n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, 
      n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, 
      n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, 
      n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, 
      n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, 
      n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, 
      n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, 
      n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, 
      n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, 
      n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, 
      n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, 
      n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, 
      n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, 
      n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, 
      n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, 
      n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, 
      n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, 
      n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, 
      n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, 
      n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, 
      n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, 
      n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, 
      n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, 
      n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, 
      n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, 
      n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, 
      n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, 
      n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, 
      n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, 
      n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, 
      n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, 
      n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, 
      n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, 
      n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, 
      n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, 
      n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, 
      n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, 
      n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, 
      n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, 
      n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, 
      n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, 
      n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, 
      n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, 
      n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, 
      n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, 
      n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, 
      n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, 
      n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, 
      n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, 
      n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, 
      n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, 
      n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, 
      n20470, n25143, n25144, n25145, n25146, n25147, n25148, n25150, n25151, 
      n25152, n25153, n25154, n25155, n25157, n25158, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n25183, n25184, n25185, 
      n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, 
      n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, 
      n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, 
      n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, 
      n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, 
      n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, 
      n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, 
      n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, 
      n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, 
      n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, 
      n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, 
      n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, 
      n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, 
      n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, 
      n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, 
      n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, 
      n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, 
      n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, 
      n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, 
      n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, 
      n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, 
      n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, 
      n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, 
      n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, 
      n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, 
      n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, 
      n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, 
      n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, 
      n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, 
      n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, 
      n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, 
      n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, 
      n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, 
      n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, 
      n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, 
      n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, 
      n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, 
      n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, 
      n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, 
      n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, 
      n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, 
      n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, 
      n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, 
      n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, 
      n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, 
      n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, 
      n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, 
      n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, 
      n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, 
      n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, 
      n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, 
      n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, 
      n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, 
      n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, 
      n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, 
      n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, 
      n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, 
      n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, 
      n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, 
      n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, 
      n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, 
      n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, 
      n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, 
      n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, 
      n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, 
      n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, 
      n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, 
      n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, 
      n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, 
      n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, 
      n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, 
      n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, 
      n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, 
      n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, 
      n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, 
      n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, 
      n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, 
      n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, 
      n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, 
      n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, 
      n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, 
      n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, 
      n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, 
      n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, 
      n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, 
      n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, 
      n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, 
      n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, 
      n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, 
      n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, 
      n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, 
      n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, 
      n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, 
      n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, 
      n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, 
      n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, 
      n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, 
      n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, 
      n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, 
      n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, 
      n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, 
      n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, 
      n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, 
      n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, 
      n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, 
      n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, 
      n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, 
      n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, 
      n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, 
      n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, 
      n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, 
      n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, 
      n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, 
      n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, 
      n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, 
      n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, 
      n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, 
      n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, 
      n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, 
      n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, 
      n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, 
      n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, 
      n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, 
      n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, 
      n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, 
      n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, 
      n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, 
      n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, 
      n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, 
      n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, 
      n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, 
      n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, 
      n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, 
      n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, 
      n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, 
      n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, 
      n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, 
      n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, 
      n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, 
      n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, 
      n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, 
      n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, 
      n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, 
      n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, 
      n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, 
      n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, 
      n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, 
      n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, 
      n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, 
      n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, 
      n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, 
      n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, 
      n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, 
      n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, 
      n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, 
      n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, 
      n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, 
      n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, 
      n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, 
      n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, 
      n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, 
      n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, 
      n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, 
      n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, 
      n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, 
      n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, 
      n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, 
      n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, 
      n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, 
      n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, 
      n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, 
      n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, 
      n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, 
      n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, 
      n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, 
      n26761, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, 
      n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, 
      n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, 
      n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, 
      n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, 
      n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, 
      n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, 
      n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, 
      n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, 
      n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, 
      n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, 
      n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, 
      n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, 
      n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, 
      n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, 
      n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, 
      n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, 
      n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, 
      n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, 
      n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, 
      n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, 
      n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, 
      n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, 
      n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, 
      n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, 
      n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, 
      n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, 
      n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, 
      n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, 
      n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, 
      n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, 
      n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, 
      n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, 
      n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, 
      n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, 
      n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, 
      n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, 
      n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, 
      n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, 
      n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, 
      n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, 
      n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, 
      n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, 
      n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, 
      n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, 
      n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, 
      n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, 
      n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, 
      n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, 
      n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, 
      n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, 
      n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, 
      n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, 
      n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, 
      n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, 
      n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, 
      n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, 
      n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, 
      n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, 
      n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, 
      n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, 
      n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, 
      n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, 
      n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, 
      n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, 
      n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, 
      n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, 
      n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, 
      n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, 
      n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, 
      n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, 
      n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, 
      n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, 
      n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, 
      n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, 
      n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, 
      n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, 
      n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, 
      n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, 
      n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, 
      n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, 
      n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, 
      n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, 
      n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, 
      n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, 
      n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, 
      n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, 
      n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, 
      n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, 
      n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, 
      n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, 
      n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, 
      n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, 
      n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, 
      n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, 
      n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, 
      n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, 
      n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, 
      n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, 
      n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, 
      n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, 
      n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, 
      n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, 
      n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, 
      n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, 
      n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, 
      n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, 
      n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, 
      n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, 
      n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, 
      n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, 
      n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, 
      n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, 
      n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, 
      n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, 
      n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, 
      n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, 
      n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, 
      n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, 
      n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, 
      n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, 
      n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, 
      n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, 
      n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, 
      n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, 
      n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, 
      n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, 
      n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, 
      n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, 
      n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, 
      n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, 
      n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, 
      n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, 
      n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, 
      n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, 
      n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, 
      n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, 
      n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, 
      n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, 
      n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, 
      n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, 
      n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, 
      n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, 
      n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, 
      n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, 
      n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, 
      n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, 
      n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, 
      n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, 
      n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, 
      n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, 
      n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, 
      n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, 
      n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, 
      n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, 
      n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, 
      n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, 
      n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, 
      n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, 
      n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, 
      n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, 
      n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, 
      n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, 
      n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, 
      n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, 
      n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, 
      n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, 
      n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, 
      n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, 
      n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, 
      n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, 
      n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, 
      n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, 
      n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, 
      n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, 
      n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, 
      n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, 
      n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, 
      n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, 
      n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, 
      n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, 
      n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, 
      n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, 
      n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, 
      n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, 
      n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, 
      n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, 
      n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, 
      n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, 
      n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, 
      n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, 
      n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, 
      n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, 
      n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, 
      n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, 
      n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, 
      n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, 
      n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, 
      n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, 
      n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, 
      n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, 
      n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, 
      n_3812, n_3813, n_3814, n_3815, n_3816, n_3817 : std_logic;

begin
   
   clk_r_REG6666_S6 : DFFR_X1 port map( D => ENABLE, CK => CLK, RN => RESET_BAR
                           , Q => n20470, QN => n_1635);
   clk_r_REG6703_S3 : DFFR_X1 port map( D => RD1, CK => CLK, RN => RESET_BAR, Q
                           => n20468, QN => n_1636);
   clk_r_REG6701_S3 : DFFR_X1 port map( D => RD2, CK => CLK, RN => RESET_BAR, Q
                           => n20467, QN => n_1637);
   clk_r_REG6730_S5 : DFFS_X1 port map( D => n1512, CK => CLK, SN => RESET_BAR,
                           Q => n_1638, QN => n20466);
   clk_r_REG6736_S5 : DFFS_X1 port map( D => n1513, CK => CLK, SN => RESET_BAR,
                           Q => n_1639, QN => n20465);
   clk_r_REG6830_S6 : DFFR_X1 port map( D => ADD_RD1(4), CK => CLK, RN => 
                           RESET_BAR, Q => n20464, QN => n_1640);
   clk_r_REG6884_S6 : DFFR_X1 port map( D => ADD_RD2(4), CK => CLK, RN => 
                           RESET_BAR, Q => n20463, QN => n_1641);
   clk_r_REG3578_S6 : DFFR_X1 port map( D => DATAIN(31), CK => CLK, RN => 
                           RESET_BAR, Q => n20462, QN => n_1642);
   clk_r_REG3570_S6 : DFFR_X1 port map( D => DATAIN(30), CK => CLK, RN => 
                           RESET_BAR, Q => n20461, QN => n_1643);
   clk_r_REG3626_S6 : DFFR_X1 port map( D => DATAIN(29), CK => CLK, RN => 
                           RESET_BAR, Q => n20460, QN => n_1644);
   clk_r_REG3674_S12 : DFFR_X1 port map( D => DATAIN(28), CK => CLK, RN => 
                           RESET_BAR, Q => n20459, QN => n_1645);
   clk_r_REG3560_S6 : DFFR_X1 port map( D => DATAIN(27), CK => CLK, RN => 
                           RESET_BAR, Q => n20458, QN => n_1646);
   clk_r_REG3551_S6 : DFFR_X1 port map( D => DATAIN(26), CK => CLK, RN => 
                           RESET_BAR, Q => n20457, QN => n_1647);
   clk_r_REG3766_S5 : DFFR_X1 port map( D => DATAIN(25), CK => CLK, RN => 
                           RESET_BAR, Q => n20456, QN => n_1648);
   clk_r_REG3543_S12 : DFFR_X1 port map( D => DATAIN(24), CK => CLK, RN => 
                           RESET_BAR, Q => n20455, QN => n_1649);
   clk_r_REG3699_S6 : DFFR_X1 port map( D => DATAIN(23), CK => CLK, RN => 
                           RESET_BAR, Q => n20454, QN => n_1650);
   clk_r_REG3692_S5 : DFFR_X1 port map( D => DATAIN(22), CK => CLK, RN => 
                           RESET_BAR, Q => n20453, QN => n_1651);
   clk_r_REG3751_S6 : DFFR_X1 port map( D => DATAIN(21), CK => CLK, RN => 
                           RESET_BAR, Q => n20452, QN => n_1652);
   clk_r_REG3744_S6 : DFFR_X1 port map( D => DATAIN(20), CK => CLK, RN => 
                           RESET_BAR, Q => n20451, QN => n_1653);
   clk_r_REG3737_S6 : DFFR_X1 port map( D => DATAIN(19), CK => CLK, RN => 
                           RESET_BAR, Q => n20450, QN => n_1654);
   clk_r_REG3730_S12 : DFFR_X1 port map( D => DATAIN(18), CK => CLK, RN => 
                           RESET_BAR, Q => n20449, QN => n_1655);
   clk_r_REG3614_S6 : DFFR_X1 port map( D => DATAIN(17), CK => CLK, RN => 
                           RESET_BAR, Q => n20448, QN => n_1656);
   clk_r_REG3607_S12 : DFFR_X1 port map( D => DATAIN(16), CK => CLK, RN => 
                           RESET_BAR, Q => n20447, QN => n_1657);
   clk_r_REG3828_S12 : DFFR_X1 port map( D => DATAIN(15), CK => CLK, RN => 
                           RESET_BAR, Q => n20446, QN => n_1658);
   clk_r_REG3878_S5 : DFFR_X1 port map( D => DATAIN(14), CK => CLK, RN => 
                           RESET_BAR, Q => n20445, QN => n_1659);
   clk_r_REG3947_S5 : DFFR_X1 port map( D => DATAIN(13), CK => CLK, RN => 
                           RESET_BAR, Q => n20444, QN => n_1660);
   clk_r_REG3782_S5 : DFFR_X1 port map( D => DATAIN(12), CK => CLK, RN => 
                           RESET_BAR, Q => n20443, QN => n_1661);
   clk_r_REG3853_S5 : DFFR_X1 port map( D => DATAIN(11), CK => CLK, RN => 
                           RESET_BAR, Q => n20442, QN => n_1662);
   clk_r_REG3656_S15 : DFFR_X1 port map( D => DATAIN(10), CK => CLK, RN => 
                           RESET_BAR, Q => n20441, QN => n_1663);
   clk_r_REG4059_S5 : DFFR_X1 port map( D => DATAIN(9), CK => CLK, RN => 
                           RESET_BAR, Q => n20440, QN => n_1664);
   clk_r_REG3529_S12 : DFFR_X1 port map( D => DATAIN(8), CK => CLK, RN => 
                           RESET_BAR, Q => n20439, QN => n_1665);
   clk_r_REG4126_S17 : DFFR_X1 port map( D => DATAIN(7), CK => CLK, RN => 
                           RESET_BAR, Q => n20438, QN => n_1666);
   clk_r_REG3649_S7 : DFFR_X1 port map( D => DATAIN(6), CK => CLK, RN => 
                           RESET_BAR, Q => n20437, QN => n_1667);
   clk_r_REG3991_S5 : DFFR_X1 port map( D => DATAIN(5), CK => CLK, RN => 
                           RESET_BAR, Q => n20436, QN => n_1668);
   clk_r_REG4046_S5 : DFFR_X1 port map( D => DATAIN(4), CK => CLK, RN => 
                           RESET_BAR, Q => n20435, QN => n_1669);
   clk_r_REG3977_S5 : DFFR_X1 port map( D => DATAIN(3), CK => CLK, RN => 
                           RESET_BAR, Q => n20434, QN => n_1670);
   clk_r_REG3934_S5 : DFFR_X1 port map( D => DATAIN(2), CK => CLK, RN => 
                           RESET_BAR, Q => n20433, QN => n_1671);
   clk_r_REG3713_S5 : DFFR_X1 port map( D => DATAIN(1), CK => CLK, RN => 
                           RESET_BAR, Q => n20432, QN => n_1672);
   clk_r_REG3587_S5 : DFFR_X1 port map( D => DATAIN(0), CK => CLK, RN => 
                           RESET_BAR, Q => n20431, QN => n_1673);
   clk_r_REG6848_S6 : DFFR_X1 port map( D => ADD_RD1(3), CK => CLK, RN => 
                           RESET_BAR, Q => n_1674, QN => n20430);
   clk_r_REG6878_S6 : DFFR_X1 port map( D => ADD_RD2(3), CK => CLK, RN => 
                           RESET_BAR, Q => n_1675, QN => n20429);
   clk_r_REG6256_S1 : DFF_X1 port map( D => n13469, CK => CLK, Q => n_1676, QN 
                           => n20428);
   clk_r_REG6254_S1 : DFF_X1 port map( D => n13470, CK => CLK, Q => n_1677, QN 
                           => n20427);
   clk_r_REG6252_S1 : DFF_X1 port map( D => n13471, CK => CLK, Q => n_1678, QN 
                           => n20426);
   clk_r_REG6514_S1 : DFF_X1 port map( D => n13472, CK => CLK, Q => n_1679, QN 
                           => n20425);
   clk_r_REG6449_S1 : DFF_X1 port map( D => n13473, CK => CLK, Q => n_1680, QN 
                           => n20424);
   clk_r_REG5995_S1 : DFF_X1 port map( D => n13474, CK => CLK, Q => n_1681, QN 
                           => n20423);
   clk_r_REG5993_S1 : DFF_X1 port map( D => n13475, CK => CLK, Q => n_1682, QN 
                           => n20422);
   clk_r_REG6250_S1 : DFF_X1 port map( D => n13476, CK => CLK, Q => n_1683, QN 
                           => n20421);
   clk_r_REG6248_S1 : DFF_X1 port map( D => n13477, CK => CLK, Q => n_1684, QN 
                           => n20420);
   clk_r_REG6246_S1 : DFF_X1 port map( D => n13478, CK => CLK, Q => n_1685, QN 
                           => n20419);
   clk_r_REG6244_S1 : DFF_X1 port map( D => n13479, CK => CLK, Q => n_1686, QN 
                           => n20418);
   clk_r_REG6512_S1 : DFF_X1 port map( D => n13480, CK => CLK, Q => n_1687, QN 
                           => n20417);
   clk_r_REG6447_S1 : DFF_X1 port map( D => n13481, CK => CLK, Q => n_1688, QN 
                           => n20416);
   clk_r_REG6242_S1 : DFF_X1 port map( D => n13482, CK => CLK, Q => n_1689, QN 
                           => n20415);
   clk_r_REG5192_S1 : DFF_X1 port map( D => n13483, CK => CLK, Q => n_1690, QN 
                           => n20414);
   clk_r_REG6064_S1 : DFF_X1 port map( D => n13484, CK => CLK, Q => n_1691, QN 
                           => n20413);
   clk_r_REG6510_S1 : DFF_X1 port map( D => n13485, CK => CLK, Q => n_1692, QN 
                           => n20412);
   clk_r_REG5574_S1 : DFF_X1 port map( D => n13486, CK => CLK, Q => n_1693, QN 
                           => n20411);
   clk_r_REG6445_S1 : DFF_X1 port map( D => n13487, CK => CLK, Q => n_1694, QN 
                           => n20410);
   clk_r_REG5991_S1 : DFF_X1 port map( D => n13488, CK => CLK, Q => n_1695, QN 
                           => n20409);
   clk_r_REG5509_S1 : DFF_X1 port map( D => n13489, CK => CLK, Q => n_1696, QN 
                           => n20408);
   clk_r_REG5063_S1 : DFF_X1 port map( D => n13490, CK => CLK, Q => n_1697, QN 
                           => n20407);
   clk_r_REG5381_S1 : DFF_X1 port map( D => n13491, CK => CLK, Q => n_1698, QN 
                           => n20406);
   clk_r_REG6508_S1 : DFF_X1 port map( D => n13492, CK => CLK, Q => n_1699, QN 
                           => n20405);
   clk_r_REG6443_S1 : DFF_X1 port map( D => n13493, CK => CLK, Q => n_1700, QN 
                           => n20404);
   clk_r_REG6578_S1 : DFF_X1 port map( D => n13494, CK => CLK, Q => n_1701, QN 
                           => n20403);
   clk_r_REG4317_S1 : DFF_X1 port map( D => n13495, CK => CLK, Q => n_1702, QN 
                           => n20402);
   clk_r_REG5127_S1 : DFF_X1 port map( D => n13496, CK => CLK, Q => n_1703, QN 
                           => n20401);
   clk_r_REG5256_S1 : DFF_X1 port map( D => n13497, CK => CLK, Q => n_1704, QN 
                           => n20400);
   clk_r_REG4918_S1 : DFF_X1 port map( D => n13498, CK => CLK, Q => n_1705, QN 
                           => n20399);
   clk_r_REG5061_S1 : DFF_X1 port map( D => n13499, CK => CLK, Q => n_1706, QN 
                           => n20398);
   clk_r_REG5989_S1 : DFF_X1 port map( D => n13500, CK => CLK, Q => n_1707, QN 
                           => n20397);
   clk_r_REG6129_S1 : DFF_X1 port map( D => n13501, CK => CLK, Q => n_1708, QN 
                           => n20396);
   clk_r_REG6062_S1 : DFF_X1 port map( D => n13502, CK => CLK, Q => n_1709, QN 
                           => n20395);
   clk_r_REG5190_S1 : DFF_X1 port map( D => n13503, CK => CLK, Q => n_1710, QN 
                           => n20394);
   clk_r_REG6127_S1 : DFF_X1 port map( D => n13504, CK => CLK, Q => n_1711, QN 
                           => n20393);
   clk_r_REG6060_S1 : DFF_X1 port map( D => n13505, CK => CLK, Q => n_1712, QN 
                           => n20392);
   clk_r_REG5572_S1 : DFF_X1 port map( D => n13506, CK => CLK, Q => n_1713, QN 
                           => n20391);
   clk_r_REG5507_S1 : DFF_X1 port map( D => n13507, CK => CLK, Q => n_1714, QN 
                           => n20390);
   clk_r_REG5188_S1 : DFF_X1 port map( D => n13508, CK => CLK, Q => n_1715, QN 
                           => n20389);
   clk_r_REG6058_S1 : DFF_X1 port map( D => n13509, CK => CLK, Q => n_1716, QN 
                           => n20388);
   clk_r_REG5059_S1 : DFF_X1 port map( D => n13510, CK => CLK, Q => n_1717, QN 
                           => n20387);
   clk_r_REG5379_S1 : DFF_X1 port map( D => n13511, CK => CLK, Q => n_1718, QN 
                           => n20386);
   clk_r_REG4916_S1 : DFF_X1 port map( D => n13512, CK => CLK, Q => n_1719, QN 
                           => n20385);
   clk_r_REG5254_S1 : DFF_X1 port map( D => n13513, CK => CLK, Q => n_1720, QN 
                           => n20384);
   clk_r_REG5125_S1 : DFF_X1 port map( D => n13514, CK => CLK, Q => n_1721, QN 
                           => n20383);
   clk_r_REG5570_S1 : DFF_X1 port map( D => n13515, CK => CLK, Q => n_1722, QN 
                           => n20382);
   clk_r_REG4315_S1 : DFF_X1 port map( D => n13516, CK => CLK, Q => n_1723, QN 
                           => n20381);
   clk_r_REG6576_S1 : DFF_X1 port map( D => n13517, CK => CLK, Q => n_1724, QN 
                           => n20380);
   clk_r_REG4313_S1 : DFF_X1 port map( D => n13518, CK => CLK, Q => n_1725, QN 
                           => n20379);
   clk_r_REG5505_S1 : DFF_X1 port map( D => n13519, CK => CLK, Q => n_1726, QN 
                           => n20378);
   clk_r_REG5123_S1 : DFF_X1 port map( D => n13520, CK => CLK, Q => n_1727, QN 
                           => n20377);
   clk_r_REG5252_S1 : DFF_X1 port map( D => n13521, CK => CLK, Q => n_1728, QN 
                           => n20376);
   clk_r_REG5377_S1 : DFF_X1 port map( D => n13522, CK => CLK, Q => n_1729, QN 
                           => n20375);
   clk_r_REG4914_S1 : DFF_X1 port map( D => n13523, CK => CLK, Q => n_1730, QN 
                           => n20374);
   clk_r_REG5057_S1 : DFF_X1 port map( D => n13524, CK => CLK, Q => n_1731, QN 
                           => n20373);
   clk_r_REG6574_S1 : DFF_X1 port map( D => n13525, CK => CLK, Q => n_1732, QN 
                           => n20372);
   clk_r_REG5987_S1 : DFF_X1 port map( D => n13526, CK => CLK, Q => n_1733, QN 
                           => n20371);
   clk_r_REG6441_S1 : DFF_X1 port map( D => n13527, CK => CLK, Q => n_1734, QN 
                           => n20370);
   clk_r_REG6506_S1 : DFF_X1 port map( D => n13528, CK => CLK, Q => n_1735, QN 
                           => n20369);
   clk_r_REG5375_S1 : DFF_X1 port map( D => n13529, CK => CLK, Q => n_1736, QN 
                           => n20368);
   clk_r_REG5503_S1 : DFF_X1 port map( D => n13530, CK => CLK, Q => n_1737, QN 
                           => n20367);
   clk_r_REG5568_S1 : DFF_X1 port map( D => n13531, CK => CLK, Q => n_1738, QN 
                           => n20366);
   clk_r_REG5186_S1 : DFF_X1 port map( D => n13532, CK => CLK, Q => n_1739, QN 
                           => n20365);
   clk_r_REG6125_S1 : DFF_X1 port map( D => n13533, CK => CLK, Q => n_1740, QN 
                           => n20364);
   clk_r_REG6056_S1 : DFF_X1 port map( D => n13534, CK => CLK, Q => n_1741, QN 
                           => n20363);
   clk_r_REG6123_S1 : DFF_X1 port map( D => n13535, CK => CLK, Q => n_1742, QN 
                           => n20362);
   clk_r_REG5566_S1 : DFF_X1 port map( D => n13536, CK => CLK, Q => n_1743, QN 
                           => n20361);
   clk_r_REG6572_S1 : DFF_X1 port map( D => n13537, CK => CLK, Q => n_1744, QN 
                           => n20360);
   clk_r_REG5501_S1 : DFF_X1 port map( D => n13538, CK => CLK, Q => n_1745, QN 
                           => n20359);
   clk_r_REG5121_S1 : DFF_X1 port map( D => n13539, CK => CLK, Q => n_1746, QN 
                           => n20358);
   clk_r_REG4311_S1 : DFF_X1 port map( D => n13540, CK => CLK, Q => n_1747, QN 
                           => n20357);
   clk_r_REG6054_S1 : DFF_X1 port map( D => n13541, CK => CLK, Q => n_1748, QN 
                           => n20356);
   clk_r_REG6570_S1 : DFF_X1 port map( D => n13542, CK => CLK, Q => n_1749, QN 
                           => n20355);
   clk_r_REG6121_S1 : DFF_X1 port map( D => n13543, CK => CLK, Q => n_1750, QN 
                           => n20354);
   clk_r_REG5373_S1 : DFF_X1 port map( D => n13544, CK => CLK, Q => n_1751, QN 
                           => n20353);
   clk_r_REG5184_S1 : DFF_X1 port map( D => n13545, CK => CLK, Q => n_1752, QN 
                           => n20352);
   clk_r_REG6439_S1 : DFF_X1 port map( D => n13546, CK => CLK, Q => n_1753, QN 
                           => n20351);
   clk_r_REG5055_S1 : DFF_X1 port map( D => n13547, CK => CLK, Q => n_1754, QN 
                           => n20350);
   clk_r_REG4309_S1 : DFF_X1 port map( D => n13548, CK => CLK, Q => n_1755, QN 
                           => n20349);
   clk_r_REG4912_S1 : DFF_X1 port map( D => n13549, CK => CLK, Q => n_1756, QN 
                           => n20348);
   clk_r_REG6504_S1 : DFF_X1 port map( D => n13550, CK => CLK, Q => n_1757, QN 
                           => n20347);
   clk_r_REG5250_S1 : DFF_X1 port map( D => n13551, CK => CLK, Q => n_1758, QN 
                           => n20346);
   clk_r_REG4910_S1 : DFF_X1 port map( D => n13552, CK => CLK, Q => n_1759, QN 
                           => n20345);
   clk_r_REG5985_S1 : DFF_X1 port map( D => n13553, CK => CLK, Q => n_1760, QN 
                           => n20344);
   clk_r_REG5564_S1 : DFF_X1 port map( D => n13554, CK => CLK, Q => n_1761, QN 
                           => n20343);
   clk_r_REG5248_S1 : DFF_X1 port map( D => n13555, CK => CLK, Q => n_1762, QN 
                           => n20342);
   clk_r_REG5182_S1 : DFF_X1 port map( D => n13556, CK => CLK, Q => n_1763, QN 
                           => n20341);
   clk_r_REG5499_S1 : DFF_X1 port map( D => n13557, CK => CLK, Q => n_1764, QN 
                           => n20340);
   clk_r_REG6502_S1 : DFF_X1 port map( D => n13558, CK => CLK, Q => n_1765, QN 
                           => n20339);
   clk_r_REG5119_S1 : DFF_X1 port map( D => n13559, CK => CLK, Q => n_1766, QN 
                           => n20338);
   clk_r_REG4307_S1 : DFF_X1 port map( D => n13560, CK => CLK, Q => n_1767, QN 
                           => n20337);
   clk_r_REG6119_S1 : DFF_X1 port map( D => n13561, CK => CLK, Q => n_1768, QN 
                           => n20336);
   clk_r_REG6568_S1 : DFF_X1 port map( D => n13562, CK => CLK, Q => n_1769, QN 
                           => n20335);
   clk_r_REG5246_S1 : DFF_X1 port map( D => n13563, CK => CLK, Q => n_1770, QN 
                           => n20334);
   clk_r_REG5371_S1 : DFF_X1 port map( D => n13564, CK => CLK, Q => n_1771, QN 
                           => n20333);
   clk_r_REG6437_S1 : DFF_X1 port map( D => n13565, CK => CLK, Q => n_1772, QN 
                           => n20332);
   clk_r_REG5983_S1 : DFF_X1 port map( D => n13566, CK => CLK, Q => n_1773, QN 
                           => n20331);
   clk_r_REG5117_S1 : DFF_X1 port map( D => n13567, CK => CLK, Q => n_1774, QN 
                           => n20330);
   clk_r_REG5053_S1 : DFF_X1 port map( D => n13568, CK => CLK, Q => n_1775, QN 
                           => n20329);
   clk_r_REG4908_S1 : DFF_X1 port map( D => n13569, CK => CLK, Q => n_1776, QN 
                           => n20328);
   clk_r_REG4305_S1 : DFF_X1 port map( D => n13570, CK => CLK, Q => n_1777, QN 
                           => n20327);
   clk_r_REG4303_S1 : DFF_X1 port map( D => n13571, CK => CLK, Q => n_1778, QN 
                           => n20326);
   clk_r_REG4301_S1 : DFF_X1 port map( D => n13572, CK => CLK, Q => n_1779, QN 
                           => n20325);
   clk_r_REG4299_S1 : DFF_X1 port map( D => n13573, CK => CLK, Q => n_1780, QN 
                           => n20324);
   clk_r_REG4297_S1 : DFF_X1 port map( D => n13574, CK => CLK, Q => n_1781, QN 
                           => n20323);
   clk_r_REG4295_S1 : DFF_X1 port map( D => n13575, CK => CLK, Q => n_1782, QN 
                           => n20322);
   clk_r_REG4293_S1 : DFF_X1 port map( D => n13576, CK => CLK, Q => n_1783, QN 
                           => n20321);
   clk_r_REG4291_S1 : DFF_X1 port map( D => n13577, CK => CLK, Q => n_1784, QN 
                           => n20320);
   clk_r_REG6500_S1 : DFF_X1 port map( D => n13578, CK => CLK, Q => n_1785, QN 
                           => n20319);
   clk_r_REG6498_S1 : DFF_X1 port map( D => n13579, CK => CLK, Q => n_1786, QN 
                           => n20318);
   clk_r_REG6496_S1 : DFF_X1 port map( D => n13580, CK => CLK, Q => n_1787, QN 
                           => n20317);
   clk_r_REG6494_S1 : DFF_X1 port map( D => n13581, CK => CLK, Q => n_1788, QN 
                           => n20316);
   clk_r_REG6492_S1 : DFF_X1 port map( D => n13582, CK => CLK, Q => n_1789, QN 
                           => n20315);
   clk_r_REG6490_S1 : DFF_X1 port map( D => n13583, CK => CLK, Q => n_1790, QN 
                           => n20314);
   clk_r_REG6488_S1 : DFF_X1 port map( D => n13584, CK => CLK, Q => n_1791, QN 
                           => n20313);
   clk_r_REG6566_S1 : DFF_X1 port map( D => n13585, CK => CLK, Q => n_1792, QN 
                           => n20312);
   clk_r_REG6564_S1 : DFF_X1 port map( D => n13586, CK => CLK, Q => n_1793, QN 
                           => n20311);
   clk_r_REG6562_S1 : DFF_X1 port map( D => n13587, CK => CLK, Q => n_1794, QN 
                           => n20310);
   clk_r_REG6560_S1 : DFF_X1 port map( D => n13588, CK => CLK, Q => n_1795, QN 
                           => n20309);
   clk_r_REG6558_S1 : DFF_X1 port map( D => n13589, CK => CLK, Q => n_1796, QN 
                           => n20308);
   clk_r_REG6556_S1 : DFF_X1 port map( D => n13590, CK => CLK, Q => n_1797, QN 
                           => n20307);
   clk_r_REG6554_S1 : DFF_X1 port map( D => n13591, CK => CLK, Q => n_1798, QN 
                           => n20306);
   clk_r_REG6552_S1 : DFF_X1 port map( D => n13592, CK => CLK, Q => n_1799, QN 
                           => n20305);
   clk_r_REG5981_S1 : DFF_X1 port map( D => n13593, CK => CLK, Q => n_1800, QN 
                           => n20304);
   clk_r_REG5979_S1 : DFF_X1 port map( D => n13594, CK => CLK, Q => n_1801, QN 
                           => n20303);
   clk_r_REG5977_S1 : DFF_X1 port map( D => n13595, CK => CLK, Q => n_1802, QN 
                           => n20302);
   clk_r_REG6240_S1 : DFF_X1 port map( D => n13596, CK => CLK, Q => n_1803, QN 
                           => n20301);
   clk_r_REG5975_S1 : DFF_X1 port map( D => n13597, CK => CLK, Q => n_1804, QN 
                           => n20300);
   clk_r_REG5973_S1 : DFF_X1 port map( D => n13598, CK => CLK, Q => n_1805, QN 
                           => n20299);
   clk_r_REG5971_S1 : DFF_X1 port map( D => n13599, CK => CLK, Q => n_1806, QN 
                           => n20298);
   clk_r_REG6435_S1 : DFF_X1 port map( D => n13600, CK => CLK, Q => n_1807, QN 
                           => n20297);
   clk_r_REG6433_S1 : DFF_X1 port map( D => n13601, CK => CLK, Q => n_1808, QN 
                           => n20296);
   clk_r_REG5051_S1 : DFF_X1 port map( D => n13602, CK => CLK, Q => n_1809, QN 
                           => n20295);
   clk_r_REG5049_S1 : DFF_X1 port map( D => n13603, CK => CLK, Q => n_1810, QN 
                           => n20294);
   clk_r_REG5047_S1 : DFF_X1 port map( D => n13604, CK => CLK, Q => n_1811, QN 
                           => n20293);
   clk_r_REG5045_S1 : DFF_X1 port map( D => n13605, CK => CLK, Q => n_1812, QN 
                           => n20292);
   clk_r_REG5180_S1 : DFF_X1 port map( D => n13606, CK => CLK, Q => n_1813, QN 
                           => n20291);
   clk_r_REG5043_S1 : DFF_X1 port map( D => n13607, CK => CLK, Q => n_1814, QN 
                           => n20290);
   clk_r_REG5041_S1 : DFF_X1 port map( D => n13608, CK => CLK, Q => n_1815, QN 
                           => n20289);
   clk_r_REG5039_S1 : DFF_X1 port map( D => n13609, CK => CLK, Q => n_1816, QN 
                           => n20288);
   clk_r_REG6238_S1 : DFF_X1 port map( D => n13610, CK => CLK, Q => n_1817, QN 
                           => n20287);
   clk_r_REG6431_S1 : DFF_X1 port map( D => n13611, CK => CLK, Q => n_1818, QN 
                           => n20286);
   clk_r_REG6429_S1 : DFF_X1 port map( D => n13612, CK => CLK, Q => n_1819, QN 
                           => n20285);
   clk_r_REG6427_S1 : DFF_X1 port map( D => n13613, CK => CLK, Q => n_1820, QN 
                           => n20284);
   clk_r_REG6425_S1 : DFF_X1 port map( D => n13614, CK => CLK, Q => n_1821, QN 
                           => n20283);
   clk_r_REG6236_S1 : DFF_X1 port map( D => n13615, CK => CLK, Q => n_1822, QN 
                           => n20282);
   clk_r_REG4906_S1 : DFF_X1 port map( D => n13616, CK => CLK, Q => n_1823, QN 
                           => n20281);
   clk_r_REG4904_S1 : DFF_X1 port map( D => n13617, CK => CLK, Q => n_1824, QN 
                           => n20280);
   clk_r_REG4902_S1 : DFF_X1 port map( D => n13618, CK => CLK, Q => n_1825, QN 
                           => n20279);
   clk_r_REG6234_S1 : DFF_X1 port map( D => n13619, CK => CLK, Q => n_1826, QN 
                           => n20278);
   clk_r_REG6423_S1 : DFF_X1 port map( D => n13620, CK => CLK, Q => n_1827, QN 
                           => n20277);
   clk_r_REG5969_S1 : DFF_X1 port map( D => n13621, CK => CLK, Q => n_1828, QN 
                           => n20276);
   clk_r_REG4900_S1 : DFF_X1 port map( D => n13622, CK => CLK, Q => n_1829, QN 
                           => n20275);
   clk_r_REG4898_S1 : DFF_X1 port map( D => n13623, CK => CLK, Q => n_1830, QN 
                           => n20274);
   clk_r_REG4896_S1 : DFF_X1 port map( D => n13624, CK => CLK, Q => n_1831, QN 
                           => n20273);
   clk_r_REG4894_S1 : DFF_X1 port map( D => n13625, CK => CLK, Q => n_1832, QN 
                           => n20272);
   clk_r_REG4892_S1 : DFF_X1 port map( D => n13626, CK => CLK, Q => n_1833, QN 
                           => n20271);
   clk_r_REG5244_S1 : DFF_X1 port map( D => n13627, CK => CLK, Q => n_1834, QN 
                           => n20270);
   clk_r_REG5242_S1 : DFF_X1 port map( D => n13628, CK => CLK, Q => n_1835, QN 
                           => n20269);
   clk_r_REG5562_S1 : DFF_X1 port map( D => n13629, CK => CLK, Q => n_1836, QN 
                           => n20268);
   clk_r_REG6232_S1 : DFF_X1 port map( D => n13630, CK => CLK, Q => n_1837, QN 
                           => n20267);
   clk_r_REG5240_S1 : DFF_X1 port map( D => n13631, CK => CLK, Q => n_1838, QN 
                           => n20266);
   clk_r_REG5238_S1 : DFF_X1 port map( D => n13632, CK => CLK, Q => n_1839, QN 
                           => n20265);
   clk_r_REG5236_S1 : DFF_X1 port map( D => n13633, CK => CLK, Q => n_1840, QN 
                           => n20264);
   clk_r_REG5234_S1 : DFF_X1 port map( D => n13634, CK => CLK, Q => n_1841, QN 
                           => n20263);
   clk_r_REG5232_S1 : DFF_X1 port map( D => n13635, CK => CLK, Q => n_1842, QN 
                           => n20262);
   clk_r_REG5230_S1 : DFF_X1 port map( D => n13636, CK => CLK, Q => n_1843, QN 
                           => n20261);
   clk_r_REG6052_S1 : DFF_X1 port map( D => n13637, CK => CLK, Q => n_1844, QN 
                           => n20260);
   clk_r_REG6230_S1 : DFF_X1 port map( D => n13638, CK => CLK, Q => n_1845, QN 
                           => n20259);
   clk_r_REG5115_S1 : DFF_X1 port map( D => n13639, CK => CLK, Q => n_1846, QN 
                           => n20258);
   clk_r_REG5113_S1 : DFF_X1 port map( D => n13640, CK => CLK, Q => n_1847, QN 
                           => n20257);
   clk_r_REG5111_S1 : DFF_X1 port map( D => n13641, CK => CLK, Q => n_1848, QN 
                           => n20256);
   clk_r_REG5109_S1 : DFF_X1 port map( D => n13642, CK => CLK, Q => n_1849, QN 
                           => n20255);
   clk_r_REG5107_S1 : DFF_X1 port map( D => n13643, CK => CLK, Q => n_1850, QN 
                           => n20254);
   clk_r_REG5497_S1 : DFF_X1 port map( D => n13644, CK => CLK, Q => n_1851, QN 
                           => n20253);
   clk_r_REG5105_S1 : DFF_X1 port map( D => n13645, CK => CLK, Q => n_1852, QN 
                           => n20252);
   clk_r_REG5103_S1 : DFF_X1 port map( D => n13646, CK => CLK, Q => n_1853, QN 
                           => n20251);
   clk_r_REG6117_S1 : DFF_X1 port map( D => n13647, CK => CLK, Q => n_1854, QN 
                           => n20250);
   clk_r_REG6115_S1 : DFF_X1 port map( D => n13648, CK => CLK, Q => n_1855, QN 
                           => n20249);
   clk_r_REG6113_S1 : DFF_X1 port map( D => n13649, CK => CLK, Q => n_1856, QN 
                           => n20248);
   clk_r_REG6111_S1 : DFF_X1 port map( D => n13650, CK => CLK, Q => n_1857, QN 
                           => n20247);
   clk_r_REG6109_S1 : DFF_X1 port map( D => n13651, CK => CLK, Q => n_1858, QN 
                           => n20246);
   clk_r_REG6107_S1 : DFF_X1 port map( D => n13652, CK => CLK, Q => n_1859, QN 
                           => n20245);
   clk_r_REG5101_S1 : DFF_X1 port map( D => n13653, CK => CLK, Q => n_1860, QN 
                           => n20244);
   clk_r_REG6105_S1 : DFF_X1 port map( D => n13654, CK => CLK, Q => n_1861, QN 
                           => n20243);
   clk_r_REG5369_S1 : DFF_X1 port map( D => n13655, CK => CLK, Q => n_1862, QN 
                           => n20242);
   clk_r_REG5495_S1 : DFF_X1 port map( D => n13656, CK => CLK, Q => n_1863, QN 
                           => n20241);
   clk_r_REG5367_S1 : DFF_X1 port map( D => n13657, CK => CLK, Q => n_1864, QN 
                           => n20240);
   clk_r_REG5365_S1 : DFF_X1 port map( D => n13658, CK => CLK, Q => n_1865, QN 
                           => n20239);
   clk_r_REG5493_S1 : DFF_X1 port map( D => n13659, CK => CLK, Q => n_1866, QN 
                           => n20238);
   clk_r_REG5363_S1 : DFF_X1 port map( D => n13660, CK => CLK, Q => n_1867, QN 
                           => n20237);
   clk_r_REG5361_S1 : DFF_X1 port map( D => n13661, CK => CLK, Q => n_1868, QN 
                           => n20236);
   clk_r_REG5359_S1 : DFF_X1 port map( D => n13662, CK => CLK, Q => n_1869, QN 
                           => n20235);
   clk_r_REG5357_S1 : DFF_X1 port map( D => n13663, CK => CLK, Q => n_1870, QN 
                           => n20234);
   clk_r_REG5355_S1 : DFF_X1 port map( D => n13664, CK => CLK, Q => n_1871, QN 
                           => n20233);
   clk_r_REG5560_S1 : DFF_X1 port map( D => n13665, CK => CLK, Q => n_1872, QN 
                           => n20232);
   clk_r_REG5558_S1 : DFF_X1 port map( D => n13666, CK => CLK, Q => n_1873, QN 
                           => n20231);
   clk_r_REG5556_S1 : DFF_X1 port map( D => n13667, CK => CLK, Q => n_1874, QN 
                           => n20230);
   clk_r_REG5554_S1 : DFF_X1 port map( D => n13668, CK => CLK, Q => n_1875, QN 
                           => n20229);
   clk_r_REG5552_S1 : DFF_X1 port map( D => n13669, CK => CLK, Q => n_1876, QN 
                           => n20228);
   clk_r_REG5550_S1 : DFF_X1 port map( D => n13670, CK => CLK, Q => n_1877, QN 
                           => n20227);
   clk_r_REG5548_S1 : DFF_X1 port map( D => n13671, CK => CLK, Q => n_1878, QN 
                           => n20226);
   clk_r_REG5491_S1 : DFF_X1 port map( D => n13672, CK => CLK, Q => n_1879, QN 
                           => n20225);
   clk_r_REG5489_S1 : DFF_X1 port map( D => n13673, CK => CLK, Q => n_1880, QN 
                           => n20224);
   clk_r_REG5487_S1 : DFF_X1 port map( D => n13674, CK => CLK, Q => n_1881, QN 
                           => n20223);
   clk_r_REG5485_S1 : DFF_X1 port map( D => n13675, CK => CLK, Q => n_1882, QN 
                           => n20222);
   clk_r_REG5483_S1 : DFF_X1 port map( D => n13676, CK => CLK, Q => n_1883, QN 
                           => n20221);
   clk_r_REG6192_S1 : DFF_X1 port map( D => n13677, CK => CLK, Q => n_1884, QN 
                           => n20220);
   clk_r_REG6190_S1 : DFF_X1 port map( D => n13678, CK => CLK, Q => n_1885, QN 
                           => n20219);
   clk_r_REG6188_S1 : DFF_X1 port map( D => n13679, CK => CLK, Q => n_1886, QN 
                           => n20218);
   clk_r_REG6186_S1 : DFF_X1 port map( D => n13680, CK => CLK, Q => n_1887, QN 
                           => n20217);
   clk_r_REG6184_S1 : DFF_X1 port map( D => n13681, CK => CLK, Q => n_1888, QN 
                           => n20216);
   clk_r_REG6182_S1 : DFF_X1 port map( D => n13682, CK => CLK, Q => n_1889, QN 
                           => n20215);
   clk_r_REG4768_S1 : DFF_X1 port map( D => n13683, CK => CLK, Q => n_1890, QN 
                           => n20214);
   clk_r_REG4766_S1 : DFF_X1 port map( D => n13684, CK => CLK, Q => n_1891, QN 
                           => n20213);
   clk_r_REG4764_S1 : DFF_X1 port map( D => n13685, CK => CLK, Q => n_1892, QN 
                           => n20212);
   clk_r_REG4762_S1 : DFF_X1 port map( D => n13686, CK => CLK, Q => n_1893, QN 
                           => n20211);
   clk_r_REG6642_S1 : DFF_X1 port map( D => n13687, CK => CLK, Q => n_1894, QN 
                           => n20210);
   clk_r_REG6640_S1 : DFF_X1 port map( D => n13688, CK => CLK, Q => n_1895, QN 
                           => n20209);
   clk_r_REG5178_S1 : DFF_X1 port map( D => n13689, CK => CLK, Q => n_1896, QN 
                           => n20208);
   clk_r_REG6638_S1 : DFF_X1 port map( D => n13690, CK => CLK, Q => n_1897, QN 
                           => n20207);
   clk_r_REG6636_S1 : DFF_X1 port map( D => n13691, CK => CLK, Q => n_1898, QN 
                           => n20206);
   clk_r_REG6634_S1 : DFF_X1 port map( D => n13692, CK => CLK, Q => n_1899, QN 
                           => n20205);
   clk_r_REG4760_S1 : DFF_X1 port map( D => n13693, CK => CLK, Q => n_1900, QN 
                           => n20204);
   clk_r_REG5176_S1 : DFF_X1 port map( D => n13694, CK => CLK, Q => n_1901, QN 
                           => n20203);
   clk_r_REG5174_S1 : DFF_X1 port map( D => n13695, CK => CLK, Q => n_1902, QN 
                           => n20202);
   clk_r_REG4758_S1 : DFF_X1 port map( D => n13696, CK => CLK, Q => n_1903, QN 
                           => n20201);
   clk_r_REG6632_S1 : DFF_X1 port map( D => n13697, CK => CLK, Q => n_1904, QN 
                           => n20200);
   clk_r_REG5172_S1 : DFF_X1 port map( D => n13698, CK => CLK, Q => n_1905, QN 
                           => n20199);
   clk_r_REG5170_S1 : DFF_X1 port map( D => n13699, CK => CLK, Q => n_1906, QN 
                           => n20198);
   clk_r_REG5168_S1 : DFF_X1 port map( D => n13700, CK => CLK, Q => n_1907, QN 
                           => n20197);
   clk_r_REG4756_S1 : DFF_X1 port map( D => n13701, CK => CLK, Q => n_1908, QN 
                           => n20196);
   clk_r_REG4850_S1 : DFF_X1 port map( D => n13702, CK => CLK, Q => n_1909, QN 
                           => n20195);
   clk_r_REG4848_S1 : DFF_X1 port map( D => n13703, CK => CLK, Q => n_1910, QN 
                           => n20194);
   clk_r_REG4754_S1 : DFF_X1 port map( D => n13704, CK => CLK, Q => n_1911, QN 
                           => n20193);
   clk_r_REG6630_S1 : DFF_X1 port map( D => n13705, CK => CLK, Q => n_1912, QN 
                           => n20192);
   clk_r_REG4846_S1 : DFF_X1 port map( D => n13706, CK => CLK, Q => n_1913, QN 
                           => n20191);
   clk_r_REG4566_S1 : DFF_X1 port map( D => n13707, CK => CLK, Q => n_1914, QN 
                           => n20190);
   clk_r_REG4564_S1 : DFF_X1 port map( D => n13708, CK => CLK, Q => n_1915, QN 
                           => n20189);
   clk_r_REG4996_S1 : DFF_X1 port map( D => n13709, CK => CLK, Q => n_1916, QN 
                           => n20188);
   clk_r_REG4994_S1 : DFF_X1 port map( D => n13710, CK => CLK, Q => n_1917, QN 
                           => n20187);
   clk_r_REG5166_S1 : DFF_X1 port map( D => n13711, CK => CLK, Q => n_1918, QN 
                           => n20186);
   clk_r_REG4562_S1 : DFF_X1 port map( D => n13712, CK => CLK, Q => n_1919, QN 
                           => n20185);
   clk_r_REG4992_S1 : DFF_X1 port map( D => n13713, CK => CLK, Q => n_1920, QN 
                           => n20184);
   clk_r_REG4844_S1 : DFF_X1 port map( D => n13714, CK => CLK, Q => n_1921, QN 
                           => n20183);
   clk_r_REG4842_S1 : DFF_X1 port map( D => n13715, CK => CLK, Q => n_1922, QN 
                           => n20182);
   clk_r_REG4840_S1 : DFF_X1 port map( D => n13716, CK => CLK, Q => n_1923, QN 
                           => n20181);
   clk_r_REG4838_S1 : DFF_X1 port map( D => n13717, CK => CLK, Q => n_1924, QN 
                           => n20180);
   clk_r_REG4560_S1 : DFF_X1 port map( D => n13718, CK => CLK, Q => n_1925, QN 
                           => n20179);
   clk_r_REG4558_S1 : DFF_X1 port map( D => n13719, CK => CLK, Q => n_1926, QN 
                           => n20178);
   clk_r_REG5652_S1 : DFF_X1 port map( D => n13720, CK => CLK, Q => n_1927, QN 
                           => n20177);
   clk_r_REG4990_S1 : DFF_X1 port map( D => n13721, CK => CLK, Q => n_1928, QN 
                           => n20176);
   clk_r_REG4988_S1 : DFF_X1 port map( D => n13722, CK => CLK, Q => n_1929, QN 
                           => n20175);
   clk_r_REG4836_S1 : DFF_X1 port map( D => n13723, CK => CLK, Q => n_1930, QN 
                           => n20174);
   clk_r_REG5650_S1 : DFF_X1 port map( D => n13724, CK => CLK, Q => n_1931, QN 
                           => n20173);
   clk_r_REG4556_S1 : DFF_X1 port map( D => n13725, CK => CLK, Q => n_1932, QN 
                           => n20172);
   clk_r_REG6628_S1 : DFF_X1 port map( D => n13726, CK => CLK, Q => n_1933, QN 
                           => n20171);
   clk_r_REG5648_S1 : DFF_X1 port map( D => n13727, CK => CLK, Q => n_1934, QN 
                           => n20170);
   clk_r_REG5646_S1 : DFF_X1 port map( D => n13728, CK => CLK, Q => n_1935, QN 
                           => n20169);
   clk_r_REG5644_S1 : DFF_X1 port map( D => n13729, CK => CLK, Q => n_1936, QN 
                           => n20168);
   clk_r_REG5642_S1 : DFF_X1 port map( D => n13730, CK => CLK, Q => n_1937, QN 
                           => n20167);
   clk_r_REG4986_S1 : DFF_X1 port map( D => n13731, CK => CLK, Q => n_1938, QN 
                           => n20166);
   clk_r_REG5037_S1 : DFF_X1 port map( D => n13732, CK => CLK, Q => n_1939, QN 
                           => n20165);
   clk_r_REG4984_S1 : DFF_X1 port map( D => n13733, CK => CLK, Q => n_1940, QN 
                           => n20164);
   clk_r_REG4982_S1 : DFF_X1 port map( D => n13734, CK => CLK, Q => n_1941, QN 
                           => n20163);
   clk_r_REG4554_S1 : DFF_X1 port map( D => n13735, CK => CLK, Q => n_1942, QN 
                           => n20162);
   clk_r_REG6050_S1 : DFF_X1 port map( D => n13736, CK => CLK, Q => n_1943, QN 
                           => n20161);
   clk_r_REG5640_S1 : DFF_X1 port map( D => n13737, CK => CLK, Q => n_1944, QN 
                           => n20160);
   clk_r_REG6048_S1 : DFF_X1 port map( D => n13738, CK => CLK, Q => n_1945, QN 
                           => n20159);
   clk_r_REG4552_S1 : DFF_X1 port map( D => n13739, CK => CLK, Q => n_1946, QN 
                           => n20158);
   clk_r_REG6046_S1 : DFF_X1 port map( D => n13740, CK => CLK, Q => n_1947, QN 
                           => n20157);
   clk_r_REG6103_S1 : DFF_X1 port map( D => n13741, CK => CLK, Q => n_1948, QN 
                           => n20156);
   clk_r_REG6044_S1 : DFF_X1 port map( D => n13742, CK => CLK, Q => n_1949, QN 
                           => n20155);
   clk_r_REG5638_S1 : DFF_X1 port map( D => n13743, CK => CLK, Q => n_1950, QN 
                           => n20154);
   clk_r_REG6042_S1 : DFF_X1 port map( D => n13744, CK => CLK, Q => n_1951, QN 
                           => n20153);
   clk_r_REG6040_S1 : DFF_X1 port map( D => n13745, CK => CLK, Q => n_1952, QN 
                           => n20152);
   clk_r_REG6038_S1 : DFF_X1 port map( D => n13746, CK => CLK, Q => n_1953, QN 
                           => n20151);
   clk_r_REG6180_S1 : DFF_X1 port map( D => n13747, CK => CLK, Q => n_1954, QN 
                           => n20150);
   clk_r_REG6178_S1 : DFF_X1 port map( D => n13748, CK => CLK, Q => n_1955, QN 
                           => n20149);
   clk_r_REG6176_S1 : DFF_X1 port map( D => n13749, CK => CLK, Q => n_1956, QN 
                           => n20148);
   clk_r_REG6174_S1 : DFF_X1 port map( D => n13750, CK => CLK, Q => n_1957, QN 
                           => n20147);
   clk_r_REG6172_S1 : DFF_X1 port map( D => n13751, CK => CLK, Q => n_1958, QN 
                           => n20146);
   clk_r_REG6170_S1 : DFF_X1 port map( D => n13752, CK => CLK, Q => n_1959, QN 
                           => n20145);
   clk_r_REG6168_S1 : DFF_X1 port map( D => n13753, CK => CLK, Q => n_1960, QN 
                           => n20144);
   clk_r_REG6166_S1 : DFF_X1 port map( D => n13754, CK => CLK, Q => n_1961, QN 
                           => n20143);
   clk_r_REG4830_S1 : DFF_X1 port map( D => n13755, CK => CLK, Q => n_1962, QN 
                           => n20142);
   clk_r_REG6622_S1 : DFF_X1 port map( D => n13756, CK => CLK, Q => n_1963, QN 
                           => n20141);
   clk_r_REG5632_S1 : DFF_X1 port map( D => n13757, CK => CLK, Q => n_1964, QN 
                           => n20140);
   clk_r_REG4748_S1 : DFF_X1 port map( D => n13758, CK => CLK, Q => n_1965, QN 
                           => n20139);
   clk_r_REG4746_S1 : DFF_X1 port map( D => n13759, CK => CLK, Q => n_1966, QN 
                           => n20138);
   clk_r_REG4546_S1 : DFF_X1 port map( D => n13760, CK => CLK, Q => n_1967, QN 
                           => n20137);
   clk_r_REG4828_S1 : DFF_X1 port map( D => n13761, CK => CLK, Q => n_1968, QN 
                           => n20136);
   clk_r_REG4976_S1 : DFF_X1 port map( D => n13762, CK => CLK, Q => n_1969, QN 
                           => n20135);
   clk_r_REG5630_S1 : DFF_X1 port map( D => n13763, CK => CLK, Q => n_1970, QN 
                           => n20134);
   clk_r_REG5628_S1 : DFF_X1 port map( D => n13764, CK => CLK, Q => n_1971, QN 
                           => n20133);
   clk_r_REG6620_S1 : DFF_X1 port map( D => n13765, CK => CLK, Q => n_1972, QN 
                           => n20132);
   clk_r_REG6618_S1 : DFF_X1 port map( D => n13766, CK => CLK, Q => n_1973, QN 
                           => n20131);
   clk_r_REG4974_S1 : DFF_X1 port map( D => n13767, CK => CLK, Q => n_1974, QN 
                           => n20130);
   clk_r_REG5626_S1 : DFF_X1 port map( D => n13768, CK => CLK, Q => n_1975, QN 
                           => n20129);
   clk_r_REG4972_S1 : DFF_X1 port map( D => n13769, CK => CLK, Q => n_1976, QN 
                           => n20128);
   clk_r_REG4826_S1 : DFF_X1 port map( D => n13770, CK => CLK, Q => n_1977, QN 
                           => n20127);
   clk_r_REG5624_S1 : DFF_X1 port map( D => n13771, CK => CLK, Q => n_1978, QN 
                           => n20126);
   clk_r_REG4544_S1 : DFF_X1 port map( D => n13772, CK => CLK, Q => n_1979, QN 
                           => n20125);
   clk_r_REG4744_S1 : DFF_X1 port map( D => n13773, CK => CLK, Q => n_1980, QN 
                           => n20124);
   clk_r_REG6616_S1 : DFF_X1 port map( D => n13774, CK => CLK, Q => n_1981, QN 
                           => n20123);
   clk_r_REG4542_S1 : DFF_X1 port map( D => n13775, CK => CLK, Q => n_1982, QN 
                           => n20122);
   clk_r_REG4742_S1 : DFF_X1 port map( D => n13776, CK => CLK, Q => n_1983, QN 
                           => n20121);
   clk_r_REG4540_S1 : DFF_X1 port map( D => n13777, CK => CLK, Q => n_1984, QN 
                           => n20120);
   clk_r_REG4740_S1 : DFF_X1 port map( D => n13778, CK => CLK, Q => n_1985, QN 
                           => n20119);
   clk_r_REG4970_S1 : DFF_X1 port map( D => n13779, CK => CLK, Q => n_1986, QN 
                           => n20118);
   clk_r_REG4538_S1 : DFF_X1 port map( D => n13780, CK => CLK, Q => n_1987, QN 
                           => n20117);
   clk_r_REG4536_S1 : DFF_X1 port map( D => n13781, CK => CLK, Q => n_1988, QN 
                           => n20116);
   clk_r_REG6614_S1 : DFF_X1 port map( D => n13782, CK => CLK, Q => n_1989, QN 
                           => n20115);
   clk_r_REG4824_S1 : DFF_X1 port map( D => n13783, CK => CLK, Q => n_1990, QN 
                           => n20114);
   clk_r_REG6612_S1 : DFF_X1 port map( D => n13784, CK => CLK, Q => n_1991, QN 
                           => n20113);
   clk_r_REG4968_S1 : DFF_X1 port map( D => n13785, CK => CLK, Q => n_1992, QN 
                           => n20112);
   clk_r_REG4822_S1 : DFF_X1 port map( D => n13786, CK => CLK, Q => n_1993, QN 
                           => n20111);
   clk_r_REG4738_S1 : DFF_X1 port map( D => n13787, CK => CLK, Q => n_1994, QN 
                           => n20110);
   clk_r_REG5622_S1 : DFF_X1 port map( D => n13788, CK => CLK, Q => n_1995, QN 
                           => n20109);
   clk_r_REG4820_S1 : DFF_X1 port map( D => n13789, CK => CLK, Q => n_1996, QN 
                           => n20108);
   clk_r_REG4966_S1 : DFF_X1 port map( D => n13790, CK => CLK, Q => n_1997, QN 
                           => n20107);
   clk_r_REG5909_S1 : DFF_X1 port map( D => n13791, CK => CLK, Q => n_1998, QN 
                           => n20106);
   clk_r_REG5907_S1 : DFF_X1 port map( D => n13792, CK => CLK, Q => n_1999, QN 
                           => n20105);
   clk_r_REG5905_S1 : DFF_X1 port map( D => n13793, CK => CLK, Q => n_2000, QN 
                           => n20104);
   clk_r_REG5903_S1 : DFF_X1 port map( D => n13794, CK => CLK, Q => n_2001, QN 
                           => n20103);
   clk_r_REG5901_S1 : DFF_X1 port map( D => n13795, CK => CLK, Q => n_2002, QN 
                           => n20102);
   clk_r_REG5899_S1 : DFF_X1 port map( D => n13796, CK => CLK, Q => n_2003, QN 
                           => n20101);
   clk_r_REG6220_S1 : DFF_X1 port map( D => n13797, CK => CLK, Q => n_2004, QN 
                           => n20100);
   clk_r_REG6478_S1 : DFF_X1 port map( D => n13798, CK => CLK, Q => n_2005, QN 
                           => n20099);
   clk_r_REG4283_S1 : DFF_X1 port map( D => n13799, CK => CLK, Q => n_2006, QN 
                           => n20098);
   clk_r_REG5897_S1 : DFF_X1 port map( D => n13800, CK => CLK, Q => n_2007, QN 
                           => n20097);
   clk_r_REG5542_S1 : DFF_X1 port map( D => n13801, CK => CLK, Q => n_2008, QN 
                           => n20096);
   clk_r_REG4886_S1 : DFF_X1 port map( D => n13802, CK => CLK, Q => n_2009, QN 
                           => n20095);
   clk_r_REG5961_S1 : DFF_X1 port map( D => n13803, CK => CLK, Q => n_2010, QN 
                           => n20094);
   clk_r_REG5959_S1 : DFF_X1 port map( D => n13804, CK => CLK, Q => n_2011, QN 
                           => n20093);
   clk_r_REG6546_S1 : DFF_X1 port map( D => n13805, CK => CLK, Q => n_2012, QN 
                           => n20092);
   clk_r_REG6415_S1 : DFF_X1 port map( D => n13806, CK => CLK, Q => n_2013, QN 
                           => n20091);
   clk_r_REG5095_S1 : DFF_X1 port map( D => n13807, CK => CLK, Q => n_2014, QN 
                           => n20090);
   clk_r_REG4281_S1 : DFF_X1 port map( D => n13808, CK => CLK, Q => n_2015, QN 
                           => n20089);
   clk_r_REG4884_S1 : DFF_X1 port map( D => n13809, CK => CLK, Q => n_2016, QN 
                           => n20088);
   clk_r_REG5093_S1 : DFF_X1 port map( D => n13810, CK => CLK, Q => n_2017, QN 
                           => n20087);
   clk_r_REG5224_S1 : DFF_X1 port map( D => n13811, CK => CLK, Q => n_2018, QN 
                           => n20086);
   clk_r_REG5349_S1 : DFF_X1 port map( D => n13812, CK => CLK, Q => n_2019, QN 
                           => n20085);
   clk_r_REG6097_S1 : DFF_X1 port map( D => n13813, CK => CLK, Q => n_2020, QN 
                           => n20084);
   clk_r_REG5957_S1 : DFF_X1 port map( D => n13814, CK => CLK, Q => n_2021, QN 
                           => n20083);
   clk_r_REG5031_S1 : DFF_X1 port map( D => n13815, CK => CLK, Q => n_2022, QN 
                           => n20082);
   clk_r_REG6218_S1 : DFF_X1 port map( D => n13816, CK => CLK, Q => n_2023, QN 
                           => n20081);
   clk_r_REG6095_S1 : DFF_X1 port map( D => n13817, CK => CLK, Q => n_2024, QN 
                           => n20080);
   clk_r_REG6476_S1 : DFF_X1 port map( D => n13818, CK => CLK, Q => n_2025, QN 
                           => n20079);
   clk_r_REG4882_S1 : DFF_X1 port map( D => n13819, CK => CLK, Q => n_2026, QN 
                           => n20078);
   clk_r_REG5477_S1 : DFF_X1 port map( D => n13820, CK => CLK, Q => n_2027, QN 
                           => n20077);
   clk_r_REG5540_S1 : DFF_X1 port map( D => n13821, CK => CLK, Q => n_2028, QN 
                           => n20076);
   clk_r_REG5475_S1 : DFF_X1 port map( D => n13822, CK => CLK, Q => n_2029, QN 
                           => n20075);
   clk_r_REG5347_S1 : DFF_X1 port map( D => n13823, CK => CLK, Q => n_2030, QN 
                           => n20074);
   clk_r_REG5895_S1 : DFF_X1 port map( D => n13824, CK => CLK, Q => n_2031, QN 
                           => n20073);
   clk_r_REG5473_S1 : DFF_X1 port map( D => n13825, CK => CLK, Q => n_2032, QN 
                           => n20072);
   clk_r_REG6474_S1 : DFF_X1 port map( D => n13826, CK => CLK, Q => n_2033, QN 
                           => n20071);
   clk_r_REG5091_S1 : DFF_X1 port map( D => n13827, CK => CLK, Q => n_2034, QN 
                           => n20070);
   clk_r_REG6413_S1 : DFF_X1 port map( D => n13828, CK => CLK, Q => n_2035, QN 
                           => n20069);
   clk_r_REG6411_S1 : DFF_X1 port map( D => n13829, CK => CLK, Q => n_2036, QN 
                           => n20068);
   clk_r_REG6093_S1 : DFF_X1 port map( D => n13830, CK => CLK, Q => n_2037, QN 
                           => n20067);
   clk_r_REG5538_S1 : DFF_X1 port map( D => n13831, CK => CLK, Q => n_2038, QN 
                           => n20066);
   clk_r_REG6544_S1 : DFF_X1 port map( D => n13832, CK => CLK, Q => n_2039, QN 
                           => n20065);
   clk_r_REG4279_S1 : DFF_X1 port map( D => n13833, CK => CLK, Q => n_2040, QN 
                           => n20064);
   clk_r_REG5893_S1 : DFF_X1 port map( D => n13834, CK => CLK, Q => n_2041, QN 
                           => n20063);
   clk_r_REG6216_S1 : DFF_X1 port map( D => n13835, CK => CLK, Q => n_2042, QN 
                           => n20062);
   clk_r_REG5029_S1 : DFF_X1 port map( D => n13836, CK => CLK, Q => n_2043, QN 
                           => n20061);
   clk_r_REG6542_S1 : DFF_X1 port map( D => n13837, CK => CLK, Q => n_2044, QN 
                           => n20060);
   clk_r_REG5027_S1 : DFF_X1 port map( D => n13838, CK => CLK, Q => n_2045, QN 
                           => n20059);
   clk_r_REG5345_S1 : DFF_X1 port map( D => n13839, CK => CLK, Q => n_2046, QN 
                           => n20058);
   clk_r_REG5222_S1 : DFF_X1 port map( D => n13840, CK => CLK, Q => n_2047, QN 
                           => n20057);
   clk_r_REG5220_S1 : DFF_X1 port map( D => n13841, CK => CLK, Q => n_2048, QN 
                           => n20056);
   clk_r_REG4229_S1 : DFF_X1 port map( D => n13843, CK => CLK, Q => n_2049, QN 
                           => n20055);
   clk_r_REG4227_S1 : DFF_X1 port map( D => n13845, CK => CLK, Q => n_2050, QN 
                           => n20054);
   clk_r_REG4225_S1 : DFF_X1 port map( D => n13847, CK => CLK, Q => n_2051, QN 
                           => n20053);
   clk_r_REG4223_S1 : DFF_X1 port map( D => n13849, CK => CLK, Q => n_2052, QN 
                           => n20052);
   clk_r_REG4221_S1 : DFF_X1 port map( D => n13851, CK => CLK, Q => n_2053, QN 
                           => n20051);
   clk_r_REG4219_S1 : DFF_X1 port map( D => n13853, CK => CLK, Q => n_2054, QN 
                           => n20050);
   clk_r_REG6320_S1 : DFF_X1 port map( D => n13854, CK => CLK, Q => n_2055, QN 
                           => n20049);
   clk_r_REG6385_S1 : DFF_X1 port map( D => n13855, CK => CLK, Q => n_2056, QN 
                           => n20048);
   clk_r_REG5719_S1 : DFF_X1 port map( D => n13856, CK => CLK, Q => n_2057, QN 
                           => n20047);
   clk_r_REG5319_S1 : DFF_X1 port map( D => n13857, CK => CLK, Q => n_2058, QN 
                           => n20046);
   clk_r_REG5783_S1 : DFF_X1 port map( D => n13858, CK => CLK, Q => n_2059, QN 
                           => n20045);
   clk_r_REG5717_S1 : DFF_X1 port map( D => n13859, CK => CLK, Q => n_2060, QN 
                           => n20044);
   clk_r_REG5781_S1 : DFF_X1 port map( D => n13860, CK => CLK, Q => n_2061, QN 
                           => n20043);
   clk_r_REG6318_S1 : DFF_X1 port map( D => n13861, CK => CLK, Q => n_2062, QN 
                           => n20042);
   clk_r_REG5845_S1 : DFF_X1 port map( D => n13862, CK => CLK, Q => n_2063, QN 
                           => n20041);
   clk_r_REG6383_S1 : DFF_X1 port map( D => n13863, CK => CLK, Q => n_2064, QN 
                           => n20040);
   clk_r_REG5317_S1 : DFF_X1 port map( D => n13864, CK => CLK, Q => n_2065, QN 
                           => n20039);
   clk_r_REG5715_S1 : DFF_X1 port map( D => n13865, CK => CLK, Q => n_2066, QN 
                           => n20038);
   clk_r_REG5779_S1 : DFF_X1 port map( D => n13866, CK => CLK, Q => n_2067, QN 
                           => n20037);
   clk_r_REG5713_S1 : DFF_X1 port map( D => n13867, CK => CLK, Q => n_2068, QN 
                           => n20036);
   clk_r_REG6316_S1 : DFF_X1 port map( D => n13868, CK => CLK, Q => n_2069, QN 
                           => n20035);
   clk_r_REG5843_S1 : DFF_X1 port map( D => n13869, CK => CLK, Q => n_2070, QN 
                           => n20034);
   clk_r_REG6381_S1 : DFF_X1 port map( D => n13870, CK => CLK, Q => n_2071, QN 
                           => n20033);
   clk_r_REG5315_S1 : DFF_X1 port map( D => n13871, CK => CLK, Q => n_2072, QN 
                           => n20032);
   clk_r_REG5711_S1 : DFF_X1 port map( D => n13872, CK => CLK, Q => n_2073, QN 
                           => n20031);
   clk_r_REG5777_S1 : DFF_X1 port map( D => n13873, CK => CLK, Q => n_2074, QN 
                           => n20030);
   clk_r_REG5775_S1 : DFF_X1 port map( D => n13874, CK => CLK, Q => n_2075, QN 
                           => n20029);
   clk_r_REG5445_S1 : DFF_X1 port map( D => n13875, CK => CLK, Q => n_2076, QN 
                           => n20028);
   clk_r_REG6314_S1 : DFF_X1 port map( D => n13876, CK => CLK, Q => n_2077, QN 
                           => n20027);
   clk_r_REG5841_S1 : DFF_X1 port map( D => n13877, CK => CLK, Q => n_2078, QN 
                           => n20026);
   clk_r_REG6379_S1 : DFF_X1 port map( D => n13878, CK => CLK, Q => n_2079, QN 
                           => n20025);
   clk_r_REG5313_S1 : DFF_X1 port map( D => n13879, CK => CLK, Q => n_2080, QN 
                           => n20024);
   clk_r_REG6312_S1 : DFF_X1 port map( D => n13880, CK => CLK, Q => n_2081, QN 
                           => n20023);
   clk_r_REG5839_S1 : DFF_X1 port map( D => n13881, CK => CLK, Q => n_2082, QN 
                           => n20022);
   clk_r_REG6377_S1 : DFF_X1 port map( D => n13882, CK => CLK, Q => n_2083, QN 
                           => n20021);
   clk_r_REG5311_S1 : DFF_X1 port map( D => n13883, CK => CLK, Q => n_2084, QN 
                           => n20020);
   clk_r_REG5837_S1 : DFF_X1 port map( D => n13884, CK => CLK, Q => n_2085, QN 
                           => n20019);
   clk_r_REG6375_S1 : DFF_X1 port map( D => n13885, CK => CLK, Q => n_2086, QN 
                           => n20018);
   clk_r_REG5773_S1 : DFF_X1 port map( D => n13886, CK => CLK, Q => n_2087, QN 
                           => n20017);
   clk_r_REG5771_S1 : DFF_X1 port map( D => n13887, CK => CLK, Q => n_2088, QN 
                           => n20016);
   clk_r_REG5443_S1 : DFF_X1 port map( D => n13888, CK => CLK, Q => n_2089, QN 
                           => n20015);
   clk_r_REG6310_S1 : DFF_X1 port map( D => n13889, CK => CLK, Q => n_2090, QN 
                           => n20014);
   clk_r_REG5835_S1 : DFF_X1 port map( D => n13890, CK => CLK, Q => n_2091, QN 
                           => n20013);
   clk_r_REG6373_S1 : DFF_X1 port map( D => n13891, CK => CLK, Q => n_2092, QN 
                           => n20012);
   clk_r_REG5309_S1 : DFF_X1 port map( D => n13892, CK => CLK, Q => n_2093, QN 
                           => n20011);
   clk_r_REG6371_S1 : DFF_X1 port map( D => n13893, CK => CLK, Q => n_2094, QN 
                           => n20010);
   clk_r_REG5307_S1 : DFF_X1 port map( D => n13894, CK => CLK, Q => n_2095, QN 
                           => n20009);
   clk_r_REG5709_S1 : DFF_X1 port map( D => n13895, CK => CLK, Q => n_2096, QN 
                           => n20008);
   clk_r_REG5769_S1 : DFF_X1 port map( D => n13896, CK => CLK, Q => n_2097, QN 
                           => n20007);
   clk_r_REG5833_S1 : DFF_X1 port map( D => n13897, CK => CLK, Q => n_2098, QN 
                           => n20006);
   clk_r_REG5831_S1 : DFF_X1 port map( D => n13898, CK => CLK, Q => n_2099, QN 
                           => n20005);
   clk_r_REG6369_S1 : DFF_X1 port map( D => n13899, CK => CLK, Q => n_2100, QN 
                           => n20004);
   clk_r_REG5441_S1 : DFF_X1 port map( D => n13901, CK => CLK, Q => n_2101, QN 
                           => n20003);
   clk_r_REG6308_S1 : DFF_X1 port map( D => n13902, CK => CLK, Q => n_2102, QN 
                           => n20002);
   clk_r_REG5829_S1 : DFF_X1 port map( D => n13903, CK => CLK, Q => n_2103, QN 
                           => n20001);
   clk_r_REG5767_S1 : DFF_X1 port map( D => n13904, CK => CLK, Q => n_2104, QN 
                           => n20000);
   clk_r_REG5305_S1 : DFF_X1 port map( D => n13905, CK => CLK, Q => n_2105, QN 
                           => n19999);
   clk_r_REG6306_S1 : DFF_X1 port map( D => n13906, CK => CLK, Q => n_2106, QN 
                           => n19998);
   clk_r_REG5707_S1 : DFF_X1 port map( D => n13907, CK => CLK, Q => n_2107, QN 
                           => n19997);
   clk_r_REG5705_S1 : DFF_X1 port map( D => n13908, CK => CLK, Q => n_2108, QN 
                           => n19996);
   clk_r_REG5827_S1 : DFF_X1 port map( D => n13909, CK => CLK, Q => n_2109, QN 
                           => n19995);
   clk_r_REG5703_S1 : DFF_X1 port map( D => n13910, CK => CLK, Q => n_2110, QN 
                           => n19994);
   clk_r_REG6367_S1 : DFF_X1 port map( D => n13911, CK => CLK, Q => n_2111, QN 
                           => n19993);
   clk_r_REG5303_S1 : DFF_X1 port map( D => n13913, CK => CLK, Q => n_2112, QN 
                           => n19992);
   clk_r_REG6304_S1 : DFF_X1 port map( D => n13914, CK => CLK, Q => n_2113, QN 
                           => n19991);
   clk_r_REG5439_S1 : DFF_X1 port map( D => n13915, CK => CLK, Q => n_2114, QN 
                           => n19990);
   clk_r_REG5437_S1 : DFF_X1 port map( D => n13917, CK => CLK, Q => n_2115, QN 
                           => n19989);
   clk_r_REG5435_S1 : DFF_X1 port map( D => n13919, CK => CLK, Q => n_2116, QN 
                           => n19988);
   clk_r_REG5301_S1 : DFF_X1 port map( D => n13920, CK => CLK, Q => n_2117, QN 
                           => n19987);
   clk_r_REG6302_S1 : DFF_X1 port map( D => n13922, CK => CLK, Q => n_2118, QN 
                           => n19986);
   clk_r_REG6300_S1 : DFF_X1 port map( D => n13923, CK => CLK, Q => n_2119, QN 
                           => n19985);
   clk_r_REG6365_S1 : DFF_X1 port map( D => n13924, CK => CLK, Q => n_2120, QN 
                           => n19984);
   clk_r_REG5471_S1 : DFF_X1 port map( D => n13925, CK => CLK, Q => n_2121, QN 
                           => n19983);
   clk_r_REG5955_S1 : DFF_X1 port map( D => n13926, CK => CLK, Q => n_2122, QN 
                           => n19982);
   clk_r_REG5299_S1 : DFF_X1 port map( D => n13927, CK => CLK, Q => n_2123, QN 
                           => n19981);
   clk_r_REG5218_S1 : DFF_X1 port map( D => n13928, CK => CLK, Q => n_2124, QN 
                           => n19980);
   clk_r_REG5089_S1 : DFF_X1 port map( D => n13929, CK => CLK, Q => n_2125, QN 
                           => n19979);
   clk_r_REG5343_S1 : DFF_X1 port map( D => n13930, CK => CLK, Q => n_2126, QN 
                           => n19978);
   clk_r_REG5891_S1 : DFF_X1 port map( D => n13931, CK => CLK, Q => n_2127, QN 
                           => n19977);
   clk_r_REG5765_S1 : DFF_X1 port map( D => n13932, CK => CLK, Q => n_2128, QN 
                           => n19976);
   clk_r_REG6472_S1 : DFF_X1 port map( D => n13933, CK => CLK, Q => n_2129, QN 
                           => n19975);
   clk_r_REG6409_S1 : DFF_X1 port map( D => n13934, CK => CLK, Q => n_2130, QN 
                           => n19974);
   clk_r_REG6091_S1 : DFF_X1 port map( D => n13935, CK => CLK, Q => n_2131, QN 
                           => n19973);
   clk_r_REG4880_S1 : DFF_X1 port map( D => n13936, CK => CLK, Q => n_2132, QN 
                           => n19972);
   clk_r_REG5536_S1 : DFF_X1 port map( D => n13937, CK => CLK, Q => n_2133, QN 
                           => n19971);
   clk_r_REG5825_S1 : DFF_X1 port map( D => n13938, CK => CLK, Q => n_2134, QN 
                           => n19970);
   clk_r_REG6540_S1 : DFF_X1 port map( D => n13939, CK => CLK, Q => n_2135, QN 
                           => n19969);
   clk_r_REG5701_S1 : DFF_X1 port map( D => n13940, CK => CLK, Q => n_2136, QN 
                           => n19968);
   clk_r_REG4277_S1 : DFF_X1 port map( D => n13941, CK => CLK, Q => n_2137, QN 
                           => n19967);
   clk_r_REG6214_S1 : DFF_X1 port map( D => n13942, CK => CLK, Q => n_2138, QN 
                           => n19966);
   clk_r_REG5025_S1 : DFF_X1 port map( D => n13943, CK => CLK, Q => n_2139, QN 
                           => n19965);
   clk_r_REG5023_S1 : DFF_X1 port map( D => n13944, CK => CLK, Q => n_2140, QN 
                           => n19964);
   clk_r_REG5433_S1 : DFF_X1 port map( D => n13945, CK => CLK, Q => n_2141, QN 
                           => n19963);
   clk_r_REG5431_S1 : DFF_X1 port map( D => n13946, CK => CLK, Q => n_2142, QN 
                           => n19962);
   clk_r_REG5021_S1 : DFF_X1 port map( D => n13947, CK => CLK, Q => n_2143, QN 
                           => n19961);
   clk_r_REG5469_S1 : DFF_X1 port map( D => n13948, CK => CLK, Q => n_2144, QN 
                           => n19960);
   clk_r_REG5467_S1 : DFF_X1 port map( D => n13949, CK => CLK, Q => n_2145, QN 
                           => n19959);
   clk_r_REG5465_S1 : DFF_X1 port map( D => n13950, CK => CLK, Q => n_2146, QN 
                           => n19958);
   clk_r_REG5429_S1 : DFF_X1 port map( D => n13951, CK => CLK, Q => n_2147, QN 
                           => n19957);
   clk_r_REG5699_S1 : DFF_X1 port map( D => n13952, CK => CLK, Q => n_2148, QN 
                           => n19956);
   clk_r_REG5697_S1 : DFF_X1 port map( D => n13953, CK => CLK, Q => n_2149, QN 
                           => n19955);
   clk_r_REG5695_S1 : DFF_X1 port map( D => n13954, CK => CLK, Q => n_2150, QN 
                           => n19954);
   clk_r_REG5763_S1 : DFF_X1 port map( D => n13955, CK => CLK, Q => n_2151, QN 
                           => n19953);
   clk_r_REG5761_S1 : DFF_X1 port map( D => n13956, CK => CLK, Q => n_2152, QN 
                           => n19952);
   clk_r_REG5759_S1 : DFF_X1 port map( D => n13957, CK => CLK, Q => n_2153, QN 
                           => n19951);
   clk_r_REG5534_S1 : DFF_X1 port map( D => n13958, CK => CLK, Q => n_2154, QN 
                           => n19950);
   clk_r_REG5532_S1 : DFF_X1 port map( D => n13959, CK => CLK, Q => n_2155, QN 
                           => n19949);
   clk_r_REG5530_S1 : DFF_X1 port map( D => n13960, CK => CLK, Q => n_2156, QN 
                           => n19948);
   clk_r_REG5019_S1 : DFF_X1 port map( D => n13961, CK => CLK, Q => n_2157, QN 
                           => n19947);
   clk_r_REG5528_S1 : DFF_X1 port map( D => n13962, CK => CLK, Q => n_2158, QN 
                           => n19946);
   clk_r_REG5463_S1 : DFF_X1 port map( D => n13963, CK => CLK, Q => n_2159, QN 
                           => n19945);
   clk_r_REG5427_S1 : DFF_X1 port map( D => n13964, CK => CLK, Q => n_2160, QN 
                           => n19944);
   clk_r_REG5757_S1 : DFF_X1 port map( D => n13965, CK => CLK, Q => n_2161, QN 
                           => n19943);
   clk_r_REG5693_S1 : DFF_X1 port map( D => n13966, CK => CLK, Q => n_2162, QN 
                           => n19942);
   clk_r_REG6486_S1 : DFF_X1 port map( D => n13967, CK => CLK, Q => n_2163, QN 
                           => n19941);
   clk_r_REG5017_S1 : DFF_X1 port map( D => n13968, CK => CLK, Q => n_2164, QN 
                           => n19940);
   clk_r_REG5526_S1 : DFF_X1 port map( D => n13969, CK => CLK, Q => n_2165, QN 
                           => n19939);
   clk_r_REG5461_S1 : DFF_X1 port map( D => n13970, CK => CLK, Q => n_2166, QN 
                           => n19938);
   clk_r_REG5425_S1 : DFF_X1 port map( D => n13971, CK => CLK, Q => n_2167, QN 
                           => n19937);
   clk_r_REG5755_S1 : DFF_X1 port map( D => n13972, CK => CLK, Q => n_2168, QN 
                           => n19936);
   clk_r_REG5691_S1 : DFF_X1 port map( D => n13973, CK => CLK, Q => n_2169, QN 
                           => n19935);
   clk_r_REG6538_S1 : DFF_X1 port map( D => n13974, CK => CLK, Q => n_2170, QN 
                           => n19934);
   clk_r_REG6536_S1 : DFF_X1 port map( D => n13975, CK => CLK, Q => n_2171, QN 
                           => n19933);
   clk_r_REG6534_S1 : DFF_X1 port map( D => n13976, CK => CLK, Q => n_2172, QN 
                           => n19932);
   clk_r_REG5015_S1 : DFF_X1 port map( D => n13977, CK => CLK, Q => n_2173, QN 
                           => n19931);
   clk_r_REG6532_S1 : DFF_X1 port map( D => n13978, CK => CLK, Q => n_2174, QN 
                           => n19930);
   clk_r_REG6530_S1 : DFF_X1 port map( D => n13979, CK => CLK, Q => n_2175, QN 
                           => n19929);
   clk_r_REG6528_S1 : DFF_X1 port map( D => n13980, CK => CLK, Q => n_2176, QN 
                           => n19928);
   clk_r_REG5524_S1 : DFF_X1 port map( D => n13981, CK => CLK, Q => n_2177, QN 
                           => n19927);
   clk_r_REG5459_S1 : DFF_X1 port map( D => n13982, CK => CLK, Q => n_2178, QN 
                           => n19926);
   clk_r_REG5423_S1 : DFF_X1 port map( D => n13983, CK => CLK, Q => n_2179, QN 
                           => n19925);
   clk_r_REG5753_S1 : DFF_X1 port map( D => n13984, CK => CLK, Q => n_2180, QN 
                           => n19924);
   clk_r_REG5689_S1 : DFF_X1 port map( D => n13985, CK => CLK, Q => n_2181, QN 
                           => n19923);
   clk_r_REG4275_S1 : DFF_X1 port map( D => n13986, CK => CLK, Q => n_2182, QN 
                           => n19922);
   clk_r_REG4273_S1 : DFF_X1 port map( D => n13987, CK => CLK, Q => n_2183, QN 
                           => n19921);
   clk_r_REG4271_S1 : DFF_X1 port map( D => n13988, CK => CLK, Q => n_2184, QN 
                           => n19920);
   clk_r_REG4269_S1 : DFF_X1 port map( D => n13989, CK => CLK, Q => n_2185, QN 
                           => n19919);
   clk_r_REG4289_S1 : DFF_X1 port map( D => n13990, CK => CLK, Q => n_2186, QN 
                           => n19918);
   clk_r_REG5889_S1 : DFF_X1 port map( D => n13991, CK => CLK, Q => n_2187, QN 
                           => n19917);
   clk_r_REG5160_S1 : DFF_X1 port map( D => n13992, CK => CLK, Q => n_2188, QN 
                           => n19916);
   clk_r_REG5158_S1 : DFF_X1 port map( D => n13993, CK => CLK, Q => n_2189, QN 
                           => n19915);
   clk_r_REG5156_S1 : DFF_X1 port map( D => n13994, CK => CLK, Q => n_2190, QN 
                           => n19914);
   clk_r_REG5154_S1 : DFF_X1 port map( D => n13995, CK => CLK, Q => n_2191, QN 
                           => n19913);
   clk_r_REG5152_S1 : DFF_X1 port map( D => n13996, CK => CLK, Q => n_2192, QN 
                           => n19912);
   clk_r_REG5150_S1 : DFF_X1 port map( D => n13997, CK => CLK, Q => n_2193, QN 
                           => n19911);
   clk_r_REG5013_S1 : DFF_X1 port map( D => n13998, CK => CLK, Q => n_2194, QN 
                           => n19910);
   clk_r_REG4267_S1 : DFF_X1 port map( D => n13999, CK => CLK, Q => n_2195, QN 
                           => n19909);
   clk_r_REG6526_S1 : DFF_X1 port map( D => n14000, CK => CLK, Q => n_2196, QN 
                           => n19908);
   clk_r_REG4878_S1 : DFF_X1 port map( D => n14001, CK => CLK, Q => n_2197, QN 
                           => n19907);
   clk_r_REG4876_S1 : DFF_X1 port map( D => n14002, CK => CLK, Q => n_2198, QN 
                           => n19906);
   clk_r_REG4874_S1 : DFF_X1 port map( D => n14003, CK => CLK, Q => n_2199, QN 
                           => n19905);
   clk_r_REG4872_S1 : DFF_X1 port map( D => n14004, CK => CLK, Q => n_2200, QN 
                           => n19904);
   clk_r_REG4870_S1 : DFF_X1 port map( D => n14005, CK => CLK, Q => n_2201, QN 
                           => n19903);
   clk_r_REG4868_S1 : DFF_X1 port map( D => n14006, CK => CLK, Q => n_2202, QN 
                           => n19902);
   clk_r_REG5687_S1 : DFF_X1 port map( D => n14007, CK => CLK, Q => n_2203, QN 
                           => n19901);
   clk_r_REG5216_S1 : DFF_X1 port map( D => n14008, CK => CLK, Q => n_2204, QN 
                           => n19900);
   clk_r_REG5214_S1 : DFF_X1 port map( D => n14009, CK => CLK, Q => n_2205, QN 
                           => n19899);
   clk_r_REG5212_S1 : DFF_X1 port map( D => n14010, CK => CLK, Q => n_2206, QN 
                           => n19898);
   clk_r_REG5210_S1 : DFF_X1 port map( D => n14011, CK => CLK, Q => n_2207, QN 
                           => n19897);
   clk_r_REG5208_S1 : DFF_X1 port map( D => n14012, CK => CLK, Q => n_2208, QN 
                           => n19896);
   clk_r_REG5206_S1 : DFF_X1 port map( D => n14013, CK => CLK, Q => n_2209, QN 
                           => n19895);
   clk_r_REG5751_S1 : DFF_X1 port map( D => n14014, CK => CLK, Q => n_2210, QN 
                           => n19894);
   clk_r_REG5421_S1 : DFF_X1 port map( D => n14015, CK => CLK, Q => n_2211, QN 
                           => n19893);
   clk_r_REG5457_S1 : DFF_X1 port map( D => n14016, CK => CLK, Q => n_2212, QN 
                           => n19892);
   clk_r_REG5522_S1 : DFF_X1 port map( D => n14017, CK => CLK, Q => n_2213, QN 
                           => n19891);
   clk_r_REG5148_S1 : DFF_X1 port map( D => n14018, CK => CLK, Q => n_2214, QN 
                           => n19890);
   clk_r_REG5011_S1 : DFF_X1 port map( D => n14019, CK => CLK, Q => n_2215, QN 
                           => n19889);
   clk_r_REG4866_S1 : DFF_X1 port map( D => n14020, CK => CLK, Q => n_2216, QN 
                           => n19888);
   clk_r_REG5204_S1 : DFF_X1 port map( D => n14021, CK => CLK, Q => n_2217, QN 
                           => n19887);
   clk_r_REG5087_S1 : DFF_X1 port map( D => n14022, CK => CLK, Q => n_2218, QN 
                           => n19886);
   clk_r_REG5085_S1 : DFF_X1 port map( D => n14023, CK => CLK, Q => n_2219, QN 
                           => n19885);
   clk_r_REG5083_S1 : DFF_X1 port map( D => n14024, CK => CLK, Q => n_2220, QN 
                           => n19884);
   clk_r_REG5081_S1 : DFF_X1 port map( D => n14025, CK => CLK, Q => n_2221, QN 
                           => n19883);
   clk_r_REG5079_S1 : DFF_X1 port map( D => n14026, CK => CLK, Q => n_2222, QN 
                           => n19882);
   clk_r_REG5077_S1 : DFF_X1 port map( D => n14027, CK => CLK, Q => n_2223, QN 
                           => n19881);
   clk_r_REG5075_S1 : DFF_X1 port map( D => n14028, CK => CLK, Q => n_2224, QN 
                           => n19880);
   clk_r_REG4265_S1 : DFF_X1 port map( D => n14029, CK => CLK, Q => n_2225, QN 
                           => n19879);
   clk_r_REG6524_S1 : DFF_X1 port map( D => n14030, CK => CLK, Q => n_2226, QN 
                           => n19878);
   clk_r_REG5887_S1 : DFF_X1 port map( D => n14031, CK => CLK, Q => n_2227, QN 
                           => n19877);
   clk_r_REG5885_S1 : DFF_X1 port map( D => n14032, CK => CLK, Q => n_2228, QN 
                           => n19876);
   clk_r_REG5883_S1 : DFF_X1 port map( D => n14033, CK => CLK, Q => n_2229, QN 
                           => n19875);
   clk_r_REG5881_S1 : DFF_X1 port map( D => n14034, CK => CLK, Q => n_2230, QN 
                           => n19874);
   clk_r_REG5879_S1 : DFF_X1 port map( D => n14035, CK => CLK, Q => n_2231, QN 
                           => n19873);
   clk_r_REG5877_S1 : DFF_X1 port map( D => n14036, CK => CLK, Q => n_2232, QN 
                           => n19872);
   clk_r_REG4263_S1 : DFF_X1 port map( D => n14037, CK => CLK, Q => n_2233, QN 
                           => n19871);
   clk_r_REG5297_S1 : DFF_X1 port map( D => n14038, CK => CLK, Q => n_2234, QN 
                           => n19870);
   clk_r_REG5295_S1 : DFF_X1 port map( D => n14039, CK => CLK, Q => n_2235, QN 
                           => n19869);
   clk_r_REG5293_S1 : DFF_X1 port map( D => n14040, CK => CLK, Q => n_2236, QN 
                           => n19868);
   clk_r_REG5291_S1 : DFF_X1 port map( D => n14041, CK => CLK, Q => n_2237, QN 
                           => n19867);
   clk_r_REG6522_S1 : DFF_X1 port map( D => n14042, CK => CLK, Q => n_2238, QN 
                           => n19866);
   clk_r_REG4261_S1 : DFF_X1 port map( D => n14043, CK => CLK, Q => n_2239, QN 
                           => n19865);
   clk_r_REG5875_S1 : DFF_X1 port map( D => n14044, CK => CLK, Q => n_2240, QN 
                           => n19864);
   clk_r_REG5073_S1 : DFF_X1 port map( D => n14045, CK => CLK, Q => n_2241, QN 
                           => n19863);
   clk_r_REG5202_S1 : DFF_X1 port map( D => n14046, CK => CLK, Q => n_2242, QN 
                           => n19862);
   clk_r_REG4864_S1 : DFF_X1 port map( D => n14047, CK => CLK, Q => n_2243, QN 
                           => n19861);
   clk_r_REG5009_S1 : DFF_X1 port map( D => n14048, CK => CLK, Q => n_2244, QN 
                           => n19860);
   clk_r_REG6407_S1 : DFF_X1 port map( D => n14049, CK => CLK, Q => n_2245, QN 
                           => n19859);
   clk_r_REG5146_S1 : DFF_X1 port map( D => n14050, CK => CLK, Q => n_2246, QN 
                           => n19858);
   clk_r_REG5520_S1 : DFF_X1 port map( D => n14051, CK => CLK, Q => n_2247, QN 
                           => n19857);
   clk_r_REG6405_S1 : DFF_X1 port map( D => n14052, CK => CLK, Q => n_2248, QN 
                           => n19856);
   clk_r_REG6421_S1 : DFF_X1 port map( D => n14053, CK => CLK, Q => n_2249, QN 
                           => n19855);
   clk_r_REG6403_S1 : DFF_X1 port map( D => n14054, CK => CLK, Q => n_2250, QN 
                           => n19854);
   clk_r_REG6401_S1 : DFF_X1 port map( D => n14055, CK => CLK, Q => n_2251, QN 
                           => n19853);
   clk_r_REG6399_S1 : DFF_X1 port map( D => n14056, CK => CLK, Q => n_2252, QN 
                           => n19852);
   clk_r_REG6419_S1 : DFF_X1 port map( D => n14057, CK => CLK, Q => n_2253, QN 
                           => n19851);
   clk_r_REG6397_S1 : DFF_X1 port map( D => n14058, CK => CLK, Q => n_2254, QN 
                           => n19850);
   clk_r_REG5685_S1 : DFF_X1 port map( D => n14059, CK => CLK, Q => n_2255, QN 
                           => n19849);
   clk_r_REG6395_S1 : DFF_X1 port map( D => n14060, CK => CLK, Q => n_2256, QN 
                           => n19848);
   clk_r_REG5455_S1 : DFF_X1 port map( D => n14061, CK => CLK, Q => n_2257, QN 
                           => n19847);
   clk_r_REG5419_S1 : DFF_X1 port map( D => n14062, CK => CLK, Q => n_2258, QN 
                           => n19846);
   clk_r_REG5749_S1 : DFF_X1 port map( D => n14063, CK => CLK, Q => n_2259, QN 
                           => n19845);
   clk_r_REG5683_S1 : DFF_X1 port map( D => n14064, CK => CLK, Q => n_2260, QN 
                           => n19844);
   clk_r_REG5747_S1 : DFF_X1 port map( D => n14065, CK => CLK, Q => n_2261, QN 
                           => n19843);
   clk_r_REG5417_S1 : DFF_X1 port map( D => n14066, CK => CLK, Q => n_2262, QN 
                           => n19842);
   clk_r_REG5453_S1 : DFF_X1 port map( D => n14067, CK => CLK, Q => n_2263, QN 
                           => n19841);
   clk_r_REG6393_S1 : DFF_X1 port map( D => n14068, CK => CLK, Q => n_2264, QN 
                           => n19840);
   clk_r_REG5518_S1 : DFF_X1 port map( D => n14069, CK => CLK, Q => n_2265, QN 
                           => n19839);
   clk_r_REG5144_S1 : DFF_X1 port map( D => n14070, CK => CLK, Q => n_2266, QN 
                           => n19838);
   clk_r_REG5823_S1 : DFF_X1 port map( D => n14071, CK => CLK, Q => n_2267, QN 
                           => n19837);
   clk_r_REG5821_S1 : DFF_X1 port map( D => n14072, CK => CLK, Q => n_2268, QN 
                           => n19836);
   clk_r_REG5007_S1 : DFF_X1 port map( D => n14073, CK => CLK, Q => n_2269, QN 
                           => n19835);
   clk_r_REG4862_S1 : DFF_X1 port map( D => n14074, CK => CLK, Q => n_2270, QN 
                           => n19834);
   clk_r_REG5200_S1 : DFF_X1 port map( D => n14075, CK => CLK, Q => n_2271, QN 
                           => n19833);
   clk_r_REG5071_S1 : DFF_X1 port map( D => n14076, CK => CLK, Q => n_2272, QN 
                           => n19832);
   clk_r_REG5819_S1 : DFF_X1 port map( D => n14077, CK => CLK, Q => n_2273, QN 
                           => n19831);
   clk_r_REG5817_S1 : DFF_X1 port map( D => n14078, CK => CLK, Q => n_2274, QN 
                           => n19830);
   clk_r_REG5873_S1 : DFF_X1 port map( D => n14079, CK => CLK, Q => n_2275, QN 
                           => n19829);
   clk_r_REG5815_S1 : DFF_X1 port map( D => n14080, CK => CLK, Q => n_2276, QN 
                           => n19828);
   clk_r_REG4259_S1 : DFF_X1 port map( D => n14081, CK => CLK, Q => n_2277, QN 
                           => n19827);
   clk_r_REG5813_S1 : DFF_X1 port map( D => n14082, CK => CLK, Q => n_2278, QN 
                           => n19826);
   clk_r_REG6520_S1 : DFF_X1 port map( D => n14083, CK => CLK, Q => n_2279, QN 
                           => n19825);
   clk_r_REG5811_S1 : DFF_X1 port map( D => n14084, CK => CLK, Q => n_2280, QN 
                           => n19824);
   clk_r_REG6363_S1 : DFF_X1 port map( D => n14085, CK => CLK, Q => n_2281, QN 
                           => n19823);
   clk_r_REG6361_S1 : DFF_X1 port map( D => n14086, CK => CLK, Q => n_2282, QN 
                           => n19822);
   clk_r_REG6359_S1 : DFF_X1 port map( D => n14087, CK => CLK, Q => n_2283, QN 
                           => n19821);
   clk_r_REG6357_S1 : DFF_X1 port map( D => n14088, CK => CLK, Q => n_2284, QN 
                           => n19820);
   clk_r_REG6355_S1 : DFF_X1 port map( D => n14089, CK => CLK, Q => n_2285, QN 
                           => n19819);
   clk_r_REG6353_S1 : DFF_X1 port map( D => n14090, CK => CLK, Q => n_2286, QN 
                           => n19818);
   clk_r_REG6351_S1 : DFF_X1 port map( D => n14091, CK => CLK, Q => n_2287, QN 
                           => n19817);
   clk_r_REG6349_S1 : DFF_X1 port map( D => n14092, CK => CLK, Q => n_2288, QN 
                           => n19816);
   clk_r_REG6417_S1 : DFF_X1 port map( D => n14094, CK => CLK, Q => n_2289, QN 
                           => n19815);
   clk_r_REG6298_S1 : DFF_X1 port map( D => n14095, CK => CLK, Q => n_2290, QN 
                           => n19814);
   clk_r_REG6296_S1 : DFF_X1 port map( D => n14096, CK => CLK, Q => n_2291, QN 
                           => n19813);
   clk_r_REG5289_S1 : DFF_X1 port map( D => n14097, CK => CLK, Q => n_2292, QN 
                           => n19812);
   clk_r_REG6294_S1 : DFF_X1 port map( D => n14098, CK => CLK, Q => n_2293, QN 
                           => n19811);
   clk_r_REG6292_S1 : DFF_X1 port map( D => n14099, CK => CLK, Q => n_2294, QN 
                           => n19810);
   clk_r_REG6290_S1 : DFF_X1 port map( D => n14100, CK => CLK, Q => n_2295, QN 
                           => n19809);
   clk_r_REG6288_S1 : DFF_X1 port map( D => n14101, CK => CLK, Q => n_2296, QN 
                           => n19808);
   clk_r_REG5809_S1 : DFF_X1 port map( D => n14102, CK => CLK, Q => n_2297, QN 
                           => n19807);
   clk_r_REG6286_S1 : DFF_X1 port map( D => n14103, CK => CLK, Q => n_2298, QN 
                           => n19806);
   clk_r_REG6284_S1 : DFF_X1 port map( D => n14104, CK => CLK, Q => n_2299, QN 
                           => n19805);
   clk_r_REG5481_S1 : DFF_X1 port map( D => n14105, CK => CLK, Q => n_2300, QN 
                           => n19804);
   clk_r_REG5546_S1 : DFF_X1 port map( D => n14106, CK => CLK, Q => n_2301, QN 
                           => n19803);
   clk_r_REG5164_S1 : DFF_X1 port map( D => n14107, CK => CLK, Q => n_2302, QN 
                           => n19802);
   clk_r_REG5953_S1 : DFF_X1 port map( D => n14108, CK => CLK, Q => n_2303, QN 
                           => n19801);
   clk_r_REG5951_S1 : DFF_X1 port map( D => n14109, CK => CLK, Q => n_2304, QN 
                           => n19800);
   clk_r_REG5949_S1 : DFF_X1 port map( D => n14110, CK => CLK, Q => n_2305, QN 
                           => n19799);
   clk_r_REG5967_S1 : DFF_X1 port map( D => n14111, CK => CLK, Q => n_2306, QN 
                           => n19798);
   clk_r_REG5947_S1 : DFF_X1 port map( D => n14112, CK => CLK, Q => n_2307, QN 
                           => n19797);
   clk_r_REG5945_S1 : DFF_X1 port map( D => n14113, CK => CLK, Q => n_2308, QN 
                           => n19796);
   clk_r_REG5035_S1 : DFF_X1 port map( D => n14114, CK => CLK, Q => n_2309, QN 
                           => n19795);
   clk_r_REG5943_S1 : DFF_X1 port map( D => n14115, CK => CLK, Q => n_2310, QN 
                           => n19794);
   clk_r_REG5965_S1 : DFF_X1 port map( D => n14116, CK => CLK, Q => n_2311, QN 
                           => n19793);
   clk_r_REG4890_S1 : DFF_X1 port map( D => n14117, CK => CLK, Q => n_2312, QN 
                           => n19792);
   clk_r_REG5228_S1 : DFF_X1 port map( D => n14118, CK => CLK, Q => n_2313, QN 
                           => n19791);
   clk_r_REG6550_S1 : DFF_X1 port map( D => n14119, CK => CLK, Q => n_2314, QN 
                           => n19790);
   clk_r_REG4287_S1 : DFF_X1 port map( D => n14120, CK => CLK, Q => n_2315, QN 
                           => n19789);
   clk_r_REG5941_S1 : DFF_X1 port map( D => n14121, CK => CLK, Q => n_2316, QN 
                           => n19788);
   clk_r_REG5963_S1 : DFF_X1 port map( D => n14123, CK => CLK, Q => n_2317, QN 
                           => n19787);
   clk_r_REG5099_S1 : DFF_X1 port map( D => n14124, CK => CLK, Q => n_2318, QN 
                           => n19786);
   clk_r_REG4285_S1 : DFF_X1 port map( D => n14126, CK => CLK, Q => n_2319, QN 
                           => n19785);
   clk_r_REG6548_S1 : DFF_X1 port map( D => n14128, CK => CLK, Q => n_2320, QN 
                           => n19784);
   clk_r_REG5097_S1 : DFF_X1 port map( D => n14130, CK => CLK, Q => n_2321, QN 
                           => n19783);
   clk_r_REG5226_S1 : DFF_X1 port map( D => n14132, CK => CLK, Q => n_2322, QN 
                           => n19782);
   clk_r_REG4860_S1 : DFF_X1 port map( D => n14133, CK => CLK, Q => n_2323, QN 
                           => n19781);
   clk_r_REG6282_S1 : DFF_X1 port map( D => n14134, CK => CLK, Q => n_2324, QN 
                           => n19780);
   clk_r_REG5939_S1 : DFF_X1 port map( D => n14135, CK => CLK, Q => n_2325, QN 
                           => n19779);
   clk_r_REG5807_S1 : DFF_X1 port map( D => n14136, CK => CLK, Q => n_2326, QN 
                           => n19778);
   clk_r_REG6347_S1 : DFF_X1 port map( D => n14137, CK => CLK, Q => n_2327, QN 
                           => n19777);
   clk_r_REG6391_S1 : DFF_X1 port map( D => n14138, CK => CLK, Q => n_2328, QN 
                           => n19776);
   clk_r_REG5005_S1 : DFF_X1 port map( D => n14139, CK => CLK, Q => n_2329, QN 
                           => n19775);
   clk_r_REG5142_S1 : DFF_X1 port map( D => n14140, CK => CLK, Q => n_2330, QN 
                           => n19774);
   clk_r_REG5516_S1 : DFF_X1 port map( D => n14141, CK => CLK, Q => n_2331, QN 
                           => n19773);
   clk_r_REG5451_S1 : DFF_X1 port map( D => n14142, CK => CLK, Q => n_2332, QN 
                           => n19772);
   clk_r_REG5415_S1 : DFF_X1 port map( D => n14143, CK => CLK, Q => n_2333, QN 
                           => n19771);
   clk_r_REG5745_S1 : DFF_X1 port map( D => n14144, CK => CLK, Q => n_2334, QN 
                           => n19770);
   clk_r_REG6212_S1 : DFF_X1 port map( D => n14145, CK => CLK, Q => n_2335, QN 
                           => n19769);
   clk_r_REG6210_S1 : DFF_X1 port map( D => n14146, CK => CLK, Q => n_2336, QN 
                           => n19768);
   clk_r_REG6208_S1 : DFF_X1 port map( D => n14147, CK => CLK, Q => n_2337, QN 
                           => n19767);
   clk_r_REG5681_S1 : DFF_X1 port map( D => n14148, CK => CLK, Q => n_2338, QN 
                           => n19766);
   clk_r_REG6389_S1 : DFF_X1 port map( D => n14149, CK => CLK, Q => n_2339, QN 
                           => n19765);
   clk_r_REG6228_S1 : DFF_X1 port map( D => n14150, CK => CLK, Q => n_2340, QN 
                           => n19764);
   clk_r_REG6226_S1 : DFF_X1 port map( D => n14151, CK => CLK, Q => n_2341, QN 
                           => n19763);
   clk_r_REG6206_S1 : DFF_X1 port map( D => n14152, CK => CLK, Q => n_2342, QN 
                           => n19762);
   clk_r_REG6204_S1 : DFF_X1 port map( D => n14153, CK => CLK, Q => n_2343, QN 
                           => n19761);
   clk_r_REG6202_S1 : DFF_X1 port map( D => n14154, CK => CLK, Q => n_2344, QN 
                           => n19760);
   clk_r_REG6200_S1 : DFF_X1 port map( D => n14155, CK => CLK, Q => n_2345, QN 
                           => n19759);
   clk_r_REG6198_S1 : DFF_X1 port map( D => n14156, CK => CLK, Q => n_2346, QN 
                           => n19758);
   clk_r_REG6196_S1 : DFF_X1 port map( D => n14157, CK => CLK, Q => n_2347, QN 
                           => n19757);
   clk_r_REG6224_S1 : DFF_X1 port map( D => n14158, CK => CLK, Q => n_2348, QN 
                           => n19756);
   clk_r_REG6345_S1 : DFF_X1 port map( D => n14159, CK => CLK, Q => n_2349, QN 
                           => n19755);
   clk_r_REG5805_S1 : DFF_X1 port map( D => n14160, CK => CLK, Q => n_2350, QN 
                           => n19754);
   clk_r_REG5937_S1 : DFF_X1 port map( D => n14161, CK => CLK, Q => n_2351, QN 
                           => n19753);
   clk_r_REG6280_S1 : DFF_X1 port map( D => n14162, CK => CLK, Q => n_2352, QN 
                           => n19752);
   clk_r_REG3579_S1 : DFF_X1 port map( D => n14164, CK => CLK, Q => n_2353, QN 
                           => n19751);
   clk_r_REG5479_S1 : DFF_X1 port map( D => n14166, CK => CLK, Q => n_2354, QN 
                           => n19750);
   clk_r_REG5544_S1 : DFF_X1 port map( D => n14168, CK => CLK, Q => n_2355, QN 
                           => n19749);
   clk_r_REG5162_S1 : DFF_X1 port map( D => n14170, CK => CLK, Q => n_2356, QN 
                           => n19748);
   clk_r_REG5033_S1 : DFF_X1 port map( D => n14172, CK => CLK, Q => n_2357, QN 
                           => n19747);
   clk_r_REG4888_S1 : DFF_X1 port map( D => n14174, CK => CLK, Q => n_2358, QN 
                           => n19746);
   clk_r_REG5198_S1 : DFF_X1 port map( D => n14175, CK => CLK, Q => n_2359, QN 
                           => n19745);
   clk_r_REG5069_S1 : DFF_X1 port map( D => n14176, CK => CLK, Q => n_2360, QN 
                           => n19744);
   clk_r_REG6518_S1 : DFF_X1 port map( D => n14177, CK => CLK, Q => n_2361, QN 
                           => n19743);
   clk_r_REG4257_S1 : DFF_X1 port map( D => n14178, CK => CLK, Q => n_2362, QN 
                           => n19742);
   clk_r_REG5871_S1 : DFF_X1 port map( D => n14179, CK => CLK, Q => n_2363, QN 
                           => n19741);
   clk_r_REG5287_S1 : DFF_X1 port map( D => n14180, CK => CLK, Q => n_2364, QN 
                           => n19740);
   clk_r_REG5285_S1 : DFF_X1 port map( D => n14181, CK => CLK, Q => n_2365, QN 
                           => n19739);
   clk_r_REG5283_S1 : DFF_X1 port map( D => n14182, CK => CLK, Q => n_2366, QN 
                           => n19738);
   clk_r_REG5341_S1 : DFF_X1 port map( D => n14183, CK => CLK, Q => n_2367, QN 
                           => n19737);
   clk_r_REG5339_S1 : DFF_X1 port map( D => n14184, CK => CLK, Q => n_2368, QN 
                           => n19736);
   clk_r_REG5337_S1 : DFF_X1 port map( D => n14185, CK => CLK, Q => n_2369, QN 
                           => n19735);
   clk_r_REG5335_S1 : DFF_X1 port map( D => n14186, CK => CLK, Q => n_2370, QN 
                           => n19734);
   clk_r_REG5333_S1 : DFF_X1 port map( D => n14187, CK => CLK, Q => n_2371, QN 
                           => n19733);
   clk_r_REG5331_S1 : DFF_X1 port map( D => n14188, CK => CLK, Q => n_2372, QN 
                           => n19732);
   clk_r_REG5679_S1 : DFF_X1 port map( D => n14189, CK => CLK, Q => n_2373, QN 
                           => n19731);
   clk_r_REG5743_S1 : DFF_X1 port map( D => n14190, CK => CLK, Q => n_2374, QN 
                           => n19730);
   clk_r_REG5413_S1 : DFF_X1 port map( D => n14191, CK => CLK, Q => n_2375, QN 
                           => n19729);
   clk_r_REG5449_S1 : DFF_X1 port map( D => n14192, CK => CLK, Q => n_2376, QN 
                           => n19728);
   clk_r_REG5329_S1 : DFF_X1 port map( D => n14193, CK => CLK, Q => n_2377, QN 
                           => n19727);
   clk_r_REG5353_S1 : DFF_X1 port map( D => n14194, CK => CLK, Q => n_2378, QN 
                           => n19726);
   clk_r_REG5351_S1 : DFF_X1 port map( D => n14196, CK => CLK, Q => n_2379, QN 
                           => n19725);
   clk_r_REG5327_S1 : DFF_X1 port map( D => n14197, CK => CLK, Q => n_2380, QN 
                           => n19724);
   clk_r_REG5325_S1 : DFF_X1 port map( D => n14198, CK => CLK, Q => n_2381, QN 
                           => n19723);
   clk_r_REG5323_S1 : DFF_X1 port map( D => n14199, CK => CLK, Q => n_2382, QN 
                           => n19722);
   clk_r_REG5321_S1 : DFF_X1 port map( D => n14200, CK => CLK, Q => n_2383, QN 
                           => n19721);
   clk_r_REG5514_S1 : DFF_X1 port map( D => n14201, CK => CLK, Q => n_2384, QN 
                           => n19720);
   clk_r_REG5140_S1 : DFF_X1 port map( D => n14202, CK => CLK, Q => n_2385, QN 
                           => n19719);
   clk_r_REG5003_S1 : DFF_X1 port map( D => n14203, CK => CLK, Q => n_2386, QN 
                           => n19718);
   clk_r_REG5281_S1 : DFF_X1 port map( D => n14204, CK => CLK, Q => n_2387, QN 
                           => n19717);
   clk_r_REG4858_S1 : DFF_X1 port map( D => n14205, CK => CLK, Q => n_2388, QN 
                           => n19716);
   clk_r_REG5196_S1 : DFF_X1 port map( D => n14206, CK => CLK, Q => n_2389, QN 
                           => n19715);
   clk_r_REG5067_S1 : DFF_X1 port map( D => n14207, CK => CLK, Q => n_2390, QN 
                           => n19714);
   clk_r_REG5869_S1 : DFF_X1 port map( D => n14208, CK => CLK, Q => n_2391, QN 
                           => n19713);
   clk_r_REG6032_S1 : DFF_X1 port map( D => n14209, CK => CLK, Q => n_2392, QN 
                           => n19712);
   clk_r_REG3854_S1 : DFF_X1 port map( D => n14211, CK => CLK, Q => n_2393, QN 
                           => n19711);
   clk_r_REG6030_S1 : DFF_X1 port map( D => n14212, CK => CLK, Q => n_2394, QN 
                           => n19710);
   clk_r_REG6028_S1 : DFF_X1 port map( D => n14213, CK => CLK, Q => n_2395, QN 
                           => n19709);
   clk_r_REG6026_S1 : DFF_X1 port map( D => n14214, CK => CLK, Q => n_2396, QN 
                           => n19708);
   clk_r_REG6024_S1 : DFF_X1 port map( D => n14215, CK => CLK, Q => n_2397, QN 
                           => n19707);
   clk_r_REG6022_S1 : DFF_X1 port map( D => n14216, CK => CLK, Q => n_2398, QN 
                           => n19706);
   clk_r_REG6020_S1 : DFF_X1 port map( D => n14217, CK => CLK, Q => n_2399, QN 
                           => n19705);
   clk_r_REG4060_S1 : DFF_X1 port map( D => n14219, CK => CLK, Q => n_2400, QN 
                           => n19704);
   clk_r_REG3530_S1 : DFF_X1 port map( D => n14221, CK => CLK, Q => n_2401, QN 
                           => n19703);
   clk_r_REG6018_S1 : DFF_X1 port map( D => n14222, CK => CLK, Q => n_2402, QN 
                           => n19702);
   clk_r_REG6036_S1 : DFF_X1 port map( D => n14223, CK => CLK, Q => n_2403, QN 
                           => n19701);
   clk_r_REG6034_S1 : DFF_X1 port map( D => n14225, CK => CLK, Q => n_2404, QN 
                           => n19700);
   clk_r_REG6016_S1 : DFF_X1 port map( D => n14226, CK => CLK, Q => n_2405, QN 
                           => n19699);
   clk_r_REG6014_S1 : DFF_X1 port map( D => n14227, CK => CLK, Q => n_2406, QN 
                           => n19698);
   clk_r_REG6012_S1 : DFF_X1 port map( D => n14228, CK => CLK, Q => n_2407, QN 
                           => n19697);
   clk_r_REG6222_S1 : DFF_X1 port map( D => n14230, CK => CLK, Q => n_2408, QN 
                           => n19696);
   clk_r_REG6278_S1 : DFF_X1 port map( D => n14231, CK => CLK, Q => n_2409, QN 
                           => n19695);
   clk_r_REG5935_S1 : DFF_X1 port map( D => n14232, CK => CLK, Q => n_2410, QN 
                           => n19694);
   clk_r_REG6484_S1 : DFF_X1 port map( D => n14233, CK => CLK, Q => n_2411, QN 
                           => n19693);
   clk_r_REG6470_S1 : DFF_X1 port map( D => n14234, CK => CLK, Q => n_2412, QN 
                           => n19692);
   clk_r_REG6468_S1 : DFF_X1 port map( D => n14235, CK => CLK, Q => n_2413, QN 
                           => n19691);
   clk_r_REG6466_S1 : DFF_X1 port map( D => n14236, CK => CLK, Q => n_2414, QN 
                           => n19690);
   clk_r_REG6482_S1 : DFF_X1 port map( D => n14237, CK => CLK, Q => n_2415, QN 
                           => n19689);
   clk_r_REG6464_S1 : DFF_X1 port map( D => n14238, CK => CLK, Q => n_2416, QN 
                           => n19688);
   clk_r_REG5803_S1 : DFF_X1 port map( D => n14239, CK => CLK, Q => n_2417, QN 
                           => n19687);
   clk_r_REG6343_S1 : DFF_X1 port map( D => n14240, CK => CLK, Q => n_2418, QN 
                           => n19686);
   clk_r_REG3552_S1 : DFF_X1 port map( D => n14242, CK => CLK, Q => n_2419, QN 
                           => n19685);
   clk_r_REG5279_S1 : DFF_X1 port map( D => n14243, CK => CLK, Q => n_2420, QN 
                           => n19684);
   clk_r_REG6462_S1 : DFF_X1 port map( D => n14244, CK => CLK, Q => n_2421, QN 
                           => n19683);
   clk_r_REG6089_S1 : DFF_X1 port map( D => n14245, CK => CLK, Q => n_2422, QN 
                           => n19682);
   clk_r_REG6101_S1 : DFF_X1 port map( D => n14246, CK => CLK, Q => n_2423, QN 
                           => n19681);
   clk_r_REG6099_S1 : DFF_X1 port map( D => n14248, CK => CLK, Q => n_2424, QN 
                           => n19680);
   clk_r_REG6087_S1 : DFF_X1 port map( D => n14249, CK => CLK, Q => n_2425, QN 
                           => n19679);
   clk_r_REG6085_S1 : DFF_X1 port map( D => n14250, CK => CLK, Q => n_2426, QN 
                           => n19678);
   clk_r_REG6083_S1 : DFF_X1 port map( D => n14251, CK => CLK, Q => n_2427, QN 
                           => n19677);
   clk_r_REG6081_S1 : DFF_X1 port map( D => n14252, CK => CLK, Q => n_2428, QN 
                           => n19676);
   clk_r_REG6480_S1 : DFF_X1 port map( D => n14254, CK => CLK, Q => n_2429, QN 
                           => n19675);
   clk_r_REG6460_S1 : DFF_X1 port map( D => n14255, CK => CLK, Q => n_2430, QN 
                           => n19674);
   clk_r_REG6458_S1 : DFF_X1 port map( D => n14256, CK => CLK, Q => n_2431, QN 
                           => n19673);
   clk_r_REG6079_S1 : DFF_X1 port map( D => n14257, CK => CLK, Q => n_2432, QN 
                           => n19672);
   clk_r_REG6456_S1 : DFF_X1 port map( D => n14258, CK => CLK, Q => n_2433, QN 
                           => n19671);
   clk_r_REG6454_S1 : DFF_X1 port map( D => n14259, CK => CLK, Q => n_2434, QN 
                           => n19670);
   clk_r_REG6010_S1 : DFF_X1 port map( D => n14260, CK => CLK, Q => n_2435, QN 
                           => n19669);
   clk_r_REG3627_S1 : DFF_X1 port map( D => n14262, CK => CLK, Q => n_2436, QN 
                           => n19668);
   clk_r_REG6077_S1 : DFF_X1 port map( D => n14263, CK => CLK, Q => n_2437, QN 
                           => n19667);
   clk_r_REG6075_S1 : DFF_X1 port map( D => n14264, CK => CLK, Q => n_2438, QN 
                           => n19666);
   clk_r_REG5277_S1 : DFF_X1 port map( D => n14265, CK => CLK, Q => n_2439, QN 
                           => n19665);
   clk_r_REG6073_S1 : DFF_X1 port map( D => n14266, CK => CLK, Q => n_2440, QN 
                           => n19664);
   clk_r_REG3544_S1 : DFF_X1 port map( D => n14268, CK => CLK, Q => n_2441, QN 
                           => n19663);
   clk_r_REG5677_S1 : DFF_X1 port map( D => n14269, CK => CLK, Q => n_2442, QN 
                           => n19662);
   clk_r_REG5741_S1 : DFF_X1 port map( D => n14270, CK => CLK, Q => n_2443, QN 
                           => n19661);
   clk_r_REG3752_S1 : DFF_X1 port map( D => n14272, CK => CLK, Q => n_2444, QN 
                           => n19660);
   clk_r_REG5411_S1 : DFF_X1 port map( D => n14273, CK => CLK, Q => n_2445, QN 
                           => n19659);
   clk_r_REG3738_S1 : DFF_X1 port map( D => n14275, CK => CLK, Q => n_2446, QN 
                           => n19658);
   clk_r_REG3731_S1 : DFF_X1 port map( D => n14277, CK => CLK, Q => n_2447, QN 
                           => n19657);
   clk_r_REG5138_S1 : DFF_X1 port map( D => n14278, CK => CLK, Q => n_2448, QN 
                           => n19656);
   clk_r_REG6071_S1 : DFF_X1 port map( D => n14279, CK => CLK, Q => n_2449, QN 
                           => n19655);
   clk_r_REG3948_S1 : DFF_X1 port map( D => n14281, CK => CLK, Q => n_2450, QN 
                           => n19654);
   clk_r_REG3879_S1 : DFF_X1 port map( D => n14283, CK => CLK, Q => n_2451, QN 
                           => n19653);
   clk_r_REG6069_S1 : DFF_X1 port map( D => n14284, CK => CLK, Q => n_2452, QN 
                           => n19652);
   clk_r_REG3608_S1 : DFF_X1 port map( D => n14286, CK => CLK, Q => n_2453, QN 
                           => n19651);
   clk_r_REG3783_S1 : DFF_X1 port map( D => n14288, CK => CLK, Q => n_2454, QN 
                           => n19650);
   clk_r_REG6158_S1 : DFF_X1 port map( D => n14290, CK => CLK, Q => n_2455, QN 
                           => n19649);
   clk_r_REG6156_S1 : DFF_X1 port map( D => n14292, CK => CLK, Q => n_2456, QN 
                           => n19648);
   clk_r_REG6154_S1 : DFF_X1 port map( D => n14294, CK => CLK, Q => n_2457, QN 
                           => n19647);
   clk_r_REG5867_S1 : DFF_X1 port map( D => n14296, CK => CLK, Q => n_2458, QN 
                           => n19646);
   clk_r_REG5865_S1 : DFF_X1 port map( D => n14297, CK => CLK, Q => n_2459, QN 
                           => n19645);
   clk_r_REG5863_S1 : DFF_X1 port map( D => n14298, CK => CLK, Q => n_2460, QN 
                           => n19644);
   clk_r_REG5861_S1 : DFF_X1 port map( D => n14299, CK => CLK, Q => n_2461, QN 
                           => n19643);
   clk_r_REG5859_S1 : DFF_X1 port map( D => n14300, CK => CLK, Q => n_2462, QN 
                           => n19642);
   clk_r_REG5857_S1 : DFF_X1 port map( D => n14301, CK => CLK, Q => n_2463, QN 
                           => n19641);
   clk_r_REG5855_S1 : DFF_X1 port map( D => n14302, CK => CLK, Q => n_2464, QN 
                           => n19640);
   clk_r_REG5853_S1 : DFF_X1 port map( D => n14303, CK => CLK, Q => n_2465, QN 
                           => n19639);
   clk_r_REG5851_S1 : DFF_X1 port map( D => n14304, CK => CLK, Q => n_2466, QN 
                           => n19638);
   clk_r_REG5849_S1 : DFF_X1 port map( D => n14305, CK => CLK, Q => n_2467, QN 
                           => n19637);
   clk_r_REG3657_S1 : DFF_X1 port map( D => n14307, CK => CLK, Q => n_2468, QN 
                           => n19636);
   clk_r_REG6152_S1 : DFF_X1 port map( D => n14309, CK => CLK, Q => n_2469, QN 
                           => n19635);
   clk_r_REG4217_S1 : DFF_X1 port map( D => n14310, CK => CLK, Q => n_2470, QN 
                           => n19634);
   clk_r_REG4215_S1 : DFF_X1 port map( D => n14311, CK => CLK, Q => n_2471, QN 
                           => n19633);
   clk_r_REG4213_S1 : DFF_X1 port map( D => n14312, CK => CLK, Q => n_2472, QN 
                           => n19632);
   clk_r_REG4211_S1 : DFF_X1 port map( D => n14313, CK => CLK, Q => n_2473, QN 
                           => n19631);
   clk_r_REG5409_S1 : DFF_X1 port map( D => n14315, CK => CLK, Q => n_2474, QN 
                           => n19630);
   clk_r_REG5407_S1 : DFF_X1 port map( D => n14317, CK => CLK, Q => n_2475, QN 
                           => n19629);
   clk_r_REG5405_S1 : DFF_X1 port map( D => n14319, CK => CLK, Q => n_2476, QN 
                           => n19628);
   clk_r_REG5403_S1 : DFF_X1 port map( D => n14321, CK => CLK, Q => n_2477, QN 
                           => n19627);
   clk_r_REG4209_S1 : DFF_X1 port map( D => n14322, CK => CLK, Q => n_2478, QN 
                           => n19626);
   clk_r_REG5401_S1 : DFF_X1 port map( D => n14324, CK => CLK, Q => n_2479, QN 
                           => n19625);
   clk_r_REG4207_S1 : DFF_X1 port map( D => n14325, CK => CLK, Q => n_2480, QN 
                           => n19624);
   clk_r_REG4205_S1 : DFF_X1 port map( D => n14326, CK => CLK, Q => n_2481, QN 
                           => n19623);
   clk_r_REG5399_S1 : DFF_X1 port map( D => n14328, CK => CLK, Q => n_2482, QN 
                           => n19622);
   clk_r_REG5397_S1 : DFF_X1 port map( D => n14329, CK => CLK, Q => n_2483, QN 
                           => n19621);
   clk_r_REG4203_S1 : DFF_X1 port map( D => n14331, CK => CLK, Q => n_2484, QN 
                           => n19620);
   clk_r_REG5395_S1 : DFF_X1 port map( D => n14333, CK => CLK, Q => n_2485, QN 
                           => n19619);
   clk_r_REG5675_S1 : DFF_X1 port map( D => n14335, CK => CLK, Q => n_2486, QN 
                           => n19618);
   clk_r_REG5673_S1 : DFF_X1 port map( D => n14336, CK => CLK, Q => n_2487, QN 
                           => n19617);
   clk_r_REG5739_S1 : DFF_X1 port map( D => n14338, CK => CLK, Q => n_2488, QN 
                           => n19616);
   clk_r_REG5671_S1 : DFF_X1 port map( D => n14339, CK => CLK, Q => n_2489, QN 
                           => n19615);
   clk_r_REG5737_S1 : DFF_X1 port map( D => n14340, CK => CLK, Q => n_2490, QN 
                           => n19614);
   clk_r_REG5669_S1 : DFF_X1 port map( D => n14341, CK => CLK, Q => n_2491, QN 
                           => n19613);
   clk_r_REG5667_S1 : DFF_X1 port map( D => n14342, CK => CLK, Q => n_2492, QN 
                           => n19612);
   clk_r_REG5735_S1 : DFF_X1 port map( D => n14343, CK => CLK, Q => n_2493, QN 
                           => n19611);
   clk_r_REG5275_S1 : DFF_X1 port map( D => n14345, CK => CLK, Q => n_2494, QN 
                           => n19610);
   clk_r_REG5733_S1 : DFF_X1 port map( D => n14346, CK => CLK, Q => n_2495, QN 
                           => n19609);
   clk_r_REG5665_S1 : DFF_X1 port map( D => n14347, CK => CLK, Q => n_2496, QN 
                           => n19608);
   clk_r_REG5731_S1 : DFF_X1 port map( D => n14348, CK => CLK, Q => n_2497, QN 
                           => n19607);
   clk_r_REG5729_S1 : DFF_X1 port map( D => n14349, CK => CLK, Q => n_2498, QN 
                           => n19606);
   clk_r_REG5727_S1 : DFF_X1 port map( D => n14350, CK => CLK, Q => n_2499, QN 
                           => n19605);
   clk_r_REG5725_S1 : DFF_X1 port map( D => n14351, CK => CLK, Q => n_2500, QN 
                           => n19604);
   clk_r_REG5723_S1 : DFF_X1 port map( D => n14352, CK => CLK, Q => n_2501, QN 
                           => n19603);
   clk_r_REG6164_S1 : DFF_X1 port map( D => n14354, CK => CLK, Q => n_2502, QN 
                           => n19602);
   clk_r_REG3693_S1 : DFF_X1 port map( D => n14356, CK => CLK, Q => n_2503, QN 
                           => n19601);
   clk_r_REG5273_S1 : DFF_X1 port map( D => n14357, CK => CLK, Q => n_2504, QN 
                           => n19600);
   clk_r_REG5663_S1 : DFF_X1 port map( D => n14359, CK => CLK, Q => n_2505, QN 
                           => n19599);
   clk_r_REG5393_S1 : DFF_X1 port map( D => n14360, CK => CLK, Q => n_2506, QN 
                           => n19598);
   clk_r_REG6162_S1 : DFF_X1 port map( D => n14362, CK => CLK, Q => n_2507, QN 
                           => n19597);
   clk_r_REG6276_S1 : DFF_X1 port map( D => n14364, CK => CLK, Q => n_2508, QN 
                           => n19596);
   clk_r_REG5661_S1 : DFF_X1 port map( D => n14366, CK => CLK, Q => n_2509, QN 
                           => n19595);
   clk_r_REG5659_S1 : DFF_X1 port map( D => n14367, CK => CLK, Q => n_2510, QN 
                           => n19594);
   clk_r_REG6274_S1 : DFF_X1 port map( D => n14368, CK => CLK, Q => n_2511, QN 
                           => n19593);
   clk_r_REG6272_S1 : DFF_X1 port map( D => n14369, CK => CLK, Q => n_2512, QN 
                           => n19592);
   clk_r_REG6270_S1 : DFF_X1 port map( D => n14370, CK => CLK, Q => n_2513, QN 
                           => n19591);
   clk_r_REG6268_S1 : DFF_X1 port map( D => n14371, CK => CLK, Q => n_2514, QN 
                           => n19590);
   clk_r_REG6266_S1 : DFF_X1 port map( D => n14372, CK => CLK, Q => n_2515, QN 
                           => n19589);
   clk_r_REG6160_S1 : DFF_X1 port map( D => n14374, CK => CLK, Q => n_2516, QN 
                           => n19588);
   clk_r_REG5801_S1 : DFF_X1 port map( D => n14376, CK => CLK, Q => n_2517, QN 
                           => n19587);
   clk_r_REG6264_S1 : DFF_X1 port map( D => n14377, CK => CLK, Q => n_2518, QN 
                           => n19586);
   clk_r_REG5799_S1 : DFF_X1 port map( D => n14378, CK => CLK, Q => n_2519, QN 
                           => n19585);
   clk_r_REG5797_S1 : DFF_X1 port map( D => n14379, CK => CLK, Q => n_2520, QN 
                           => n19584);
   clk_r_REG5795_S1 : DFF_X1 port map( D => n14380, CK => CLK, Q => n_2521, QN 
                           => n19583);
   clk_r_REG3700_S1 : DFF_X1 port map( D => n14382, CK => CLK, Q => n_2522, QN 
                           => n19582);
   clk_r_REG6262_S1 : DFF_X1 port map( D => n14383, CK => CLK, Q => n_2523, QN 
                           => n19581);
   clk_r_REG6341_S1 : DFF_X1 port map( D => n14385, CK => CLK, Q => n_2524, QN 
                           => n19580);
   clk_r_REG5271_S1 : DFF_X1 port map( D => n14386, CK => CLK, Q => n_2525, QN 
                           => n19579);
   clk_r_REG5793_S1 : DFF_X1 port map( D => n14387, CK => CLK, Q => n_2526, QN 
                           => n19578);
   clk_r_REG5791_S1 : DFF_X1 port map( D => n14388, CK => CLK, Q => n_2527, QN 
                           => n19577);
   clk_r_REG6260_S1 : DFF_X1 port map( D => n14389, CK => CLK, Q => n_2528, QN 
                           => n19576);
   clk_r_REG6339_S1 : DFF_X1 port map( D => n14390, CK => CLK, Q => n_2529, QN 
                           => n19575);
   clk_r_REG6337_S1 : DFF_X1 port map( D => n14391, CK => CLK, Q => n_2530, QN 
                           => n19574);
   clk_r_REG5789_S1 : DFF_X1 port map( D => n14392, CK => CLK, Q => n_2531, QN 
                           => n19573);
   clk_r_REG5787_S1 : DFF_X1 port map( D => n14393, CK => CLK, Q => n_2532, QN 
                           => n19572);
   clk_r_REG5785_S1 : DFF_X1 port map( D => n14394, CK => CLK, Q => n_2533, QN 
                           => n19571);
   clk_r_REG3675_S1 : DFF_X1 port map( D => n14396, CK => CLK, Q => n_2534, QN 
                           => n19570);
   clk_r_REG6335_S1 : DFF_X1 port map( D => n14397, CK => CLK, Q => n_2535, QN 
                           => n19569);
   clk_r_REG6333_S1 : DFF_X1 port map( D => n14398, CK => CLK, Q => n_2536, QN 
                           => n19568);
   clk_r_REG6331_S1 : DFF_X1 port map( D => n14399, CK => CLK, Q => n_2537, QN 
                           => n19567);
   clk_r_REG3571_S1 : DFF_X1 port map( D => n14401, CK => CLK, Q => n_2538, QN 
                           => n19566);
   clk_r_REG6329_S1 : DFF_X1 port map( D => n14402, CK => CLK, Q => n_2539, QN 
                           => n19565);
   clk_r_REG6327_S1 : DFF_X1 port map( D => n14403, CK => CLK, Q => n_2540, QN 
                           => n19564);
   clk_r_REG5269_S1 : DFF_X1 port map( D => n14405, CK => CLK, Q => n_2541, QN 
                           => n19563);
   clk_r_REG6325_S1 : DFF_X1 port map( D => n14407, CK => CLK, Q => n_2542, QN 
                           => n19562);
   clk_r_REG5267_S1 : DFF_X1 port map( D => n14409, CK => CLK, Q => n_2543, QN 
                           => n19561);
   clk_r_REG5265_S1 : DFF_X1 port map( D => n14411, CK => CLK, Q => n_2544, QN 
                           => n19560);
   clk_r_REG5391_S1 : DFF_X1 port map( D => n14413, CK => CLK, Q => n_2545, QN 
                           => n19559);
   clk_r_REG5263_S1 : DFF_X1 port map( D => n14415, CK => CLK, Q => n_2546, QN 
                           => n19558);
   clk_r_REG5261_S1 : DFF_X1 port map( D => n14416, CK => CLK, Q => n_2547, QN 
                           => n19557);
   clk_r_REG5259_S1 : DFF_X1 port map( D => n14418, CK => CLK, Q => n_2548, QN 
                           => n19556);
   clk_r_REG3767_S1 : DFF_X1 port map( D => n14421, CK => CLK, Q => n_2549, QN 
                           => n19555);
   clk_r_REG3561_S1 : DFF_X1 port map( D => n14424, CK => CLK, Q => n_2550, QN 
                           => n19554);
   clk_r_REG4964_S1 : DFF_X1 port map( D => n14425, CK => CLK, Q => n_2551, QN 
                           => n19553);
   clk_r_REG4962_S1 : DFF_X1 port map( D => n14426, CK => CLK, Q => n_2552, QN 
                           => n19552);
   clk_r_REG5389_S1 : DFF_X1 port map( D => n14427, CK => CLK, Q => n_2553, QN 
                           => n19551);
   clk_r_REG6008_S1 : DFF_X1 port map( D => n14428, CK => CLK, Q => n_2554, QN 
                           => n19550);
   clk_r_REG5136_S1 : DFF_X1 port map( D => n14429, CK => CLK, Q => n_2555, QN 
                           => n19549);
   clk_r_REG5387_S1 : DFF_X1 port map( D => n14430, CK => CLK, Q => n_2556, QN 
                           => n19548);
   clk_r_REG6006_S1 : DFF_X1 port map( D => n14431, CK => CLK, Q => n_2557, QN 
                           => n19547);
   clk_r_REG4960_S1 : DFF_X1 port map( D => n14432, CK => CLK, Q => n_2558, QN 
                           => n19546);
   clk_r_REG4818_S1 : DFF_X1 port map( D => n14433, CK => CLK, Q => n_2559, QN 
                           => n19545);
   clk_r_REG5385_S1 : DFF_X1 port map( D => n14434, CK => CLK, Q => n_2560, QN 
                           => n19544);
   clk_r_REG6610_S1 : DFF_X1 port map( D => n14435, CK => CLK, Q => n_2561, QN 
                           => n19543);
   clk_r_REG4197_S1 : DFF_X1 port map( D => n14436, CK => CLK, Q => n_2562, QN 
                           => n19542);
   clk_r_REG4816_S1 : DFF_X1 port map( D => n14437, CK => CLK, Q => n_2563, QN 
                           => n19541);
   clk_r_REG4534_S1 : DFF_X1 port map( D => n14438, CK => CLK, Q => n_2564, QN 
                           => n19540);
   clk_r_REG4195_S1 : DFF_X1 port map( D => n14439, CK => CLK, Q => n_2565, QN 
                           => n19539);
   clk_r_REG4736_S1 : DFF_X1 port map( D => n14440, CK => CLK, Q => n_2566, QN 
                           => n19538);
   clk_r_REG4193_S1 : DFF_X1 port map( D => n14441, CK => CLK, Q => n_2567, QN 
                           => n19537);
   clk_r_REG5620_S1 : DFF_X1 port map( D => n14442, CK => CLK, Q => n_2568, QN 
                           => n19536);
   clk_r_REG5134_S1 : DFF_X1 port map( D => n14443, CK => CLK, Q => n_2569, QN 
                           => n19535);
   clk_r_REG4814_S1 : DFF_X1 port map( D => n14444, CK => CLK, Q => n_2570, QN 
                           => n19534);
   clk_r_REG5132_S1 : DFF_X1 port map( D => n14445, CK => CLK, Q => n_2571, QN 
                           => n19533);
   clk_r_REG6004_S1 : DFF_X1 port map( D => n14446, CK => CLK, Q => n_2572, QN 
                           => n19532);
   clk_r_REG4532_S1 : DFF_X1 port map( D => n14447, CK => CLK, Q => n_2573, QN 
                           => n19531);
   clk_r_REG5618_S1 : DFF_X1 port map( D => n14448, CK => CLK, Q => n_2574, QN 
                           => n19530);
   clk_r_REG4530_S1 : DFF_X1 port map( D => n14449, CK => CLK, Q => n_2575, QN 
                           => n19529);
   clk_r_REG6608_S1 : DFF_X1 port map( D => n14451, CK => CLK, Q => n_2576, QN 
                           => n19528);
   clk_r_REG6606_S1 : DFF_X1 port map( D => n14452, CK => CLK, Q => n_2577, QN 
                           => n19527);
   clk_r_REG5616_S1 : DFF_X1 port map( D => n14453, CK => CLK, Q => n_2578, QN 
                           => n19526);
   clk_r_REG4734_S1 : DFF_X1 port map( D => n14455, CK => CLK, Q => n_2579, QN 
                           => n19525);
   clk_r_REG4732_S1 : DFF_X1 port map( D => n14457, CK => CLK, Q => n_2580, QN 
                           => n19524);
   clk_r_REG6150_S1 : DFF_X1 port map( D => n14459, CK => CLK, Q => n_2581, QN 
                           => n19523);
   clk_r_REG6148_S1 : DFF_X1 port map( D => n14461, CK => CLK, Q => n_2582, QN 
                           => n19522);
   clk_r_REG6146_S1 : DFF_X1 port map( D => n14463, CK => CLK, Q => n_2583, QN 
                           => n19521);
   clk_r_REG6144_S1 : DFF_X1 port map( D => n14465, CK => CLK, Q => n_2584, QN 
                           => n19520);
   clk_r_REG6142_S1 : DFF_X1 port map( D => n14467, CK => CLK, Q => n_2585, QN 
                           => n19519);
   clk_r_REG6140_S1 : DFF_X1 port map( D => n14469, CK => CLK, Q => n_2586, QN 
                           => n19518);
   clk_r_REG6138_S1 : DFF_X1 port map( D => n14471, CK => CLK, Q => n_2587, QN 
                           => n19517);
   clk_r_REG6136_S1 : DFF_X1 port map( D => n14473, CK => CLK, Q => n_2588, QN 
                           => n19516);
   clk_r_REG6134_S1 : DFF_X1 port map( D => n14475, CK => CLK, Q => n_2589, QN 
                           => n19515);
   clk_r_REG6132_S1 : DFF_X1 port map( D => n14477, CK => CLK, Q => n_2590, QN 
                           => n19514);
   clk_r_REG3588_S1 : DFF_X1 port map( D => n14480, CK => CLK, Q => n_2591, QN 
                           => n19513);
   clk_r_REG4812_S1 : DFF_X1 port map( D => n14481, CK => CLK, Q => n_2592, QN 
                           => n19512);
   clk_r_REG4191_S1 : DFF_X1 port map( D => n14482, CK => CLK, Q => n_2593, QN 
                           => n19511);
   clk_r_REG4958_S1 : DFF_X1 port map( D => n14483, CK => CLK, Q => n_2594, QN 
                           => n19510);
   clk_r_REG3829_S1 : DFF_X1 port map( D => n14485, CK => CLK, Q => n_2595, QN 
                           => n19509);
   clk_r_REG4730_S1 : DFF_X1 port map( D => n14486, CK => CLK, Q => n_2596, QN 
                           => n19508);
   clk_r_REG6604_S1 : DFF_X1 port map( D => n14487, CK => CLK, Q => n_2597, QN 
                           => n19507);
   clk_r_REG3745_S1 : DFF_X1 port map( D => n14489, CK => CLK, Q => n_2598, QN 
                           => n19506);
   clk_r_REG3615_S1 : DFF_X1 port map( D => n14491, CK => CLK, Q => n_2599, QN 
                           => n19505);
   clk_r_REG4528_S1 : DFF_X1 port map( D => n14492, CK => CLK, Q => n_2600, QN 
                           => n19504);
   clk_r_REG5614_S1 : DFF_X1 port map( D => n14494, CK => CLK, Q => n_2601, QN 
                           => n19503);
   clk_r_REG6626_S1 : DFF_X1 port map( D => n14495, CK => CLK, Q => n_2602, QN 
                           => n19502);
   clk_r_REG4201_S1 : DFF_X1 port map( D => n14496, CK => CLK, Q => n_2603, QN 
                           => n19501);
   clk_r_REG4980_S1 : DFF_X1 port map( D => n14497, CK => CLK, Q => n_2604, QN 
                           => n19500);
   clk_r_REG4550_S1 : DFF_X1 port map( D => n14498, CK => CLK, Q => n_2605, QN 
                           => n19499);
   clk_r_REG4199_S1 : DFF_X1 port map( D => n14500, CK => CLK, Q => n_2606, QN 
                           => n19498);
   clk_r_REG4752_S1 : DFF_X1 port map( D => n14501, CK => CLK, Q => n_2607, QN 
                           => n19497);
   clk_r_REG4750_S1 : DFF_X1 port map( D => n14503, CK => CLK, Q => n_2608, QN 
                           => n19496);
   clk_r_REG5636_S1 : DFF_X1 port map( D => n14504, CK => CLK, Q => n_2609, QN 
                           => n19495);
   clk_r_REG4978_S1 : DFF_X1 port map( D => n14506, CK => CLK, Q => n_2610, QN 
                           => n19494);
   clk_r_REG4834_S1 : DFF_X1 port map( D => n14507, CK => CLK, Q => n_2611, QN 
                           => n19493);
   clk_r_REG6624_S1 : DFF_X1 port map( D => n14509, CK => CLK, Q => n_2612, QN 
                           => n19492);
   clk_r_REG4832_S1 : DFF_X1 port map( D => n14512, CK => CLK, Q => n_2613, QN 
                           => n19491);
   clk_r_REG5634_S1 : DFF_X1 port map( D => n14514, CK => CLK, Q => n_2614, QN 
                           => n19490);
   clk_r_REG4548_S1 : DFF_X1 port map( D => n14517, CK => CLK, Q => n_2615, QN 
                           => n19489);
   clk_r_REG4526_S1 : DFF_X1 port map( D => n14518, CK => CLK, Q => n_2616, QN 
                           => n19488);
   clk_r_REG4524_S1 : DFF_X1 port map( D => n14519, CK => CLK, Q => n_2617, QN 
                           => n19487);
   clk_r_REG5612_S1 : DFF_X1 port map( D => n14520, CK => CLK, Q => n_2618, QN 
                           => n19486);
   clk_r_REG5610_S1 : DFF_X1 port map( D => n14521, CK => CLK, Q => n_2619, QN 
                           => n19485);
   clk_r_REG5608_S1 : DFF_X1 port map( D => n14522, CK => CLK, Q => n_2620, QN 
                           => n19484);
   clk_r_REG4522_S1 : DFF_X1 port map( D => n14523, CK => CLK, Q => n_2621, QN 
                           => n19483);
   clk_r_REG5606_S1 : DFF_X1 port map( D => n14524, CK => CLK, Q => n_2622, QN 
                           => n19482);
   clk_r_REG4810_S1 : DFF_X1 port map( D => n14525, CK => CLK, Q => n_2623, QN 
                           => n19481);
   clk_r_REG4956_S1 : DFF_X1 port map( D => n14526, CK => CLK, Q => n_2624, QN 
                           => n19480);
   clk_r_REG4808_S1 : DFF_X1 port map( D => n14527, CK => CLK, Q => n_2625, QN 
                           => n19479);
   clk_r_REG4806_S1 : DFF_X1 port map( D => n14528, CK => CLK, Q => n_2626, QN 
                           => n19478);
   clk_r_REG4954_S1 : DFF_X1 port map( D => n14529, CK => CLK, Q => n_2627, QN 
                           => n19477);
   clk_r_REG4804_S1 : DFF_X1 port map( D => n14530, CK => CLK, Q => n_2628, QN 
                           => n19476);
   clk_r_REG4802_S1 : DFF_X1 port map( D => n14531, CK => CLK, Q => n_2629, QN 
                           => n19475);
   clk_r_REG5604_S1 : DFF_X1 port map( D => n14532, CK => CLK, Q => n_2630, QN 
                           => n19474);
   clk_r_REG4189_S1 : DFF_X1 port map( D => n14533, CK => CLK, Q => n_2631, QN 
                           => n19473);
   clk_r_REG4520_S1 : DFF_X1 port map( D => n14534, CK => CLK, Q => n_2632, QN 
                           => n19472);
   clk_r_REG5602_S1 : DFF_X1 port map( D => n14535, CK => CLK, Q => n_2633, QN 
                           => n19471);
   clk_r_REG5600_S1 : DFF_X1 port map( D => n14536, CK => CLK, Q => n_2634, QN 
                           => n19470);
   clk_r_REG4800_S1 : DFF_X1 port map( D => n14537, CK => CLK, Q => n_2635, QN 
                           => n19469);
   clk_r_REG4798_S1 : DFF_X1 port map( D => n14538, CK => CLK, Q => n_2636, QN 
                           => n19468);
   clk_r_REG4518_S1 : DFF_X1 port map( D => n14539, CK => CLK, Q => n_2637, QN 
                           => n19467);
   clk_r_REG4516_S1 : DFF_X1 port map( D => n14540, CK => CLK, Q => n_2638, QN 
                           => n19466);
   clk_r_REG4514_S1 : DFF_X1 port map( D => n14541, CK => CLK, Q => n_2639, QN 
                           => n19465);
   clk_r_REG4512_S1 : DFF_X1 port map( D => n14542, CK => CLK, Q => n_2640, QN 
                           => n19464);
   clk_r_REG4796_S1 : DFF_X1 port map( D => n14543, CK => CLK, Q => n_2641, QN 
                           => n19463);
   clk_r_REG4952_S1 : DFF_X1 port map( D => n14544, CK => CLK, Q => n_2642, QN 
                           => n19462);
   clk_r_REG5598_S1 : DFF_X1 port map( D => n14545, CK => CLK, Q => n_2643, QN 
                           => n19461);
   clk_r_REG4728_S1 : DFF_X1 port map( D => n14546, CK => CLK, Q => n_2644, QN 
                           => n19460);
   clk_r_REG5596_S1 : DFF_X1 port map( D => n14547, CK => CLK, Q => n_2645, QN 
                           => n19459);
   clk_r_REG4726_S1 : DFF_X1 port map( D => n14548, CK => CLK, Q => n_2646, QN 
                           => n19458);
   clk_r_REG4950_S1 : DFF_X1 port map( D => n14549, CK => CLK, Q => n_2647, QN 
                           => n19457);
   clk_r_REG4724_S1 : DFF_X1 port map( D => n14550, CK => CLK, Q => n_2648, QN 
                           => n19456);
   clk_r_REG4722_S1 : DFF_X1 port map( D => n14551, CK => CLK, Q => n_2649, QN 
                           => n19455);
   clk_r_REG4794_S1 : DFF_X1 port map( D => n14552, CK => CLK, Q => n_2650, QN 
                           => n19454);
   clk_r_REG4510_S1 : DFF_X1 port map( D => n14553, CK => CLK, Q => n_2651, QN 
                           => n19453);
   clk_r_REG4720_S1 : DFF_X1 port map( D => n14554, CK => CLK, Q => n_2652, QN 
                           => n19452);
   clk_r_REG5594_S1 : DFF_X1 port map( D => n14555, CK => CLK, Q => n_2653, QN 
                           => n19451);
   clk_r_REG4718_S1 : DFF_X1 port map( D => n14556, CK => CLK, Q => n_2654, QN 
                           => n19450);
   clk_r_REG5592_S1 : DFF_X1 port map( D => n14557, CK => CLK, Q => n_2655, QN 
                           => n19449);
   clk_r_REG4716_S1 : DFF_X1 port map( D => n14558, CK => CLK, Q => n_2656, QN 
                           => n19448);
   clk_r_REG4714_S1 : DFF_X1 port map( D => n14559, CK => CLK, Q => n_2657, QN 
                           => n19447);
   clk_r_REG4792_S1 : DFF_X1 port map( D => n14560, CK => CLK, Q => n_2658, QN 
                           => n19446);
   clk_r_REG4712_S1 : DFF_X1 port map( D => n14561, CK => CLK, Q => n_2659, QN 
                           => n19445);
   clk_r_REG4710_S1 : DFF_X1 port map( D => n14562, CK => CLK, Q => n_2660, QN 
                           => n19444);
   clk_r_REG4508_S1 : DFF_X1 port map( D => n14563, CK => CLK, Q => n_2661, QN 
                           => n19443);
   clk_r_REG4790_S1 : DFF_X1 port map( D => n14564, CK => CLK, Q => n_2662, QN 
                           => n19442);
   clk_r_REG6602_S1 : DFF_X1 port map( D => n14565, CK => CLK, Q => n_2663, QN 
                           => n19441);
   clk_r_REG4506_S1 : DFF_X1 port map( D => n14566, CK => CLK, Q => n_2664, QN 
                           => n19440);
   clk_r_REG4708_S1 : DFF_X1 port map( D => n14567, CK => CLK, Q => n_2665, QN 
                           => n19439);
   clk_r_REG6600_S1 : DFF_X1 port map( D => n14568, CK => CLK, Q => n_2666, QN 
                           => n19438);
   clk_r_REG6598_S1 : DFF_X1 port map( D => n14569, CK => CLK, Q => n_2667, QN 
                           => n19437);
   clk_r_REG6596_S1 : DFF_X1 port map( D => n14570, CK => CLK, Q => n_2668, QN 
                           => n19436);
   clk_r_REG6594_S1 : DFF_X1 port map( D => n14571, CK => CLK, Q => n_2669, QN 
                           => n19435);
   clk_r_REG4187_S1 : DFF_X1 port map( D => n14572, CK => CLK, Q => n_2670, QN 
                           => n19434);
   clk_r_REG3992_S1 : DFF_X1 port map( D => n14574, CK => CLK, Q => n_2671, QN 
                           => n19433);
   clk_r_REG4948_S1 : DFF_X1 port map( D => n14575, CK => CLK, Q => n_2672, QN 
                           => n19432);
   clk_r_REG6592_S1 : DFF_X1 port map( D => n14576, CK => CLK, Q => n_2673, QN 
                           => n19431);
   clk_r_REG4946_S1 : DFF_X1 port map( D => n14577, CK => CLK, Q => n_2674, QN 
                           => n19430);
   clk_r_REG4944_S1 : DFF_X1 port map( D => n14578, CK => CLK, Q => n_2675, QN 
                           => n19429);
   clk_r_REG6590_S1 : DFF_X1 port map( D => n14579, CK => CLK, Q => n_2676, QN 
                           => n19428);
   clk_r_REG6588_S1 : DFF_X1 port map( D => n14581, CK => CLK, Q => n_2677, QN 
                           => n19427);
   clk_r_REG6586_S1 : DFF_X1 port map( D => n14582, CK => CLK, Q => n_2678, QN 
                           => n19426);
   clk_r_REG4185_S1 : DFF_X1 port map( D => n14584, CK => CLK, Q => n_2679, QN 
                           => n19425);
   clk_r_REG4942_S1 : DFF_X1 port map( D => n14585, CK => CLK, Q => n_2680, QN 
                           => n19424);
   clk_r_REG4940_S1 : DFF_X1 port map( D => n14586, CK => CLK, Q => n_2681, QN 
                           => n19423);
   clk_r_REG4183_S1 : DFF_X1 port map( D => n14587, CK => CLK, Q => n_2682, QN 
                           => n19422);
   clk_r_REG4938_S1 : DFF_X1 port map( D => n14589, CK => CLK, Q => n_2683, QN 
                           => n19421);
   clk_r_REG4181_S1 : DFF_X1 port map( D => n14590, CK => CLK, Q => n_2684, QN 
                           => n19420);
   clk_r_REG3714_S1 : DFF_X1 port map( D => n14592, CK => CLK, Q => n_2685, QN 
                           => n19419);
   clk_r_REG4936_S1 : DFF_X1 port map( D => n14593, CK => CLK, Q => n_2686, QN 
                           => n19418);
   clk_r_REG3935_S1 : DFF_X1 port map( D => n14595, CK => CLK, Q => n_2687, QN 
                           => n19417);
   clk_r_REG6584_S1 : DFF_X1 port map( D => n14596, CK => CLK, Q => n_2688, QN 
                           => n19416);
   clk_r_REG4179_S1 : DFF_X1 port map( D => n14598, CK => CLK, Q => n_2689, QN 
                           => n19415);
   clk_r_REG3978_S1 : DFF_X1 port map( D => n14600, CK => CLK, Q => n_2690, QN 
                           => n19414);
   clk_r_REG6582_S1 : DFF_X1 port map( D => n14602, CK => CLK, Q => n_2691, QN 
                           => n19413);
   clk_r_REG4047_S1 : DFF_X1 port map( D => n14605, CK => CLK, Q => n_2692, QN 
                           => n19412);
   clk_r_REG4177_S1 : DFF_X1 port map( D => n14607, CK => CLK, Q => n_2693, QN 
                           => n19411);
   clk_r_REG4175_S1 : DFF_X1 port map( D => n14609, CK => CLK, Q => n_2694, QN 
                           => n19410);
   clk_r_REG3517_S1 : DFF_X1 port map( D => n14611, CK => CLK, Q => n_2695, QN 
                           => n19409);
   clk_r_REG4173_S1 : DFF_X1 port map( D => n14613, CK => CLK, Q => n_2696, QN 
                           => n19408);
   clk_r_REG4171_S1 : DFF_X1 port map( D => n14615, CK => CLK, Q => n_2697, QN 
                           => n19407);
   clk_r_REG4169_S1 : DFF_X1 port map( D => n14617, CK => CLK, Q => n_2698, QN 
                           => n19406);
   clk_r_REG4127_S1 : DFF_X1 port map( D => n14620, CK => CLK, Q => n_2699, QN 
                           => n19405);
   clk_r_REG6737_S5 : DFFS_X1 port map( D => n1513, CK => CLK, SN => RESET_BAR,
                           Q => n19404, QN => n_2700);
   clk_r_REG6731_S5 : DFFS_X1 port map( D => n1512, CK => CLK, SN => RESET_BAR,
                           Q => n19403, QN => n_2701);
   clk_r_REG6793_S6 : DFFR_X1 port map( D => n11226, CK => CLK, RN => RESET_BAR
                           , Q => n19402, QN => n_2702);
   clk_r_REG6812_S6 : DFFS_X1 port map( D => n11227, CK => CLK, SN => RESET_BAR
                           , Q => n19401, QN => n_2703);
   clk_r_REG6899_S6 : DFFR_X1 port map( D => n11229, CK => CLK, RN => RESET_BAR
                           , Q => n19395, QN => n_2704);
   clk_r_REG6513_S1 : DFF_X1 port map( D => n13480, CK => CLK, Q => n19394, QN 
                           => n_2705);
   clk_r_REG6045_S1 : DFF_X1 port map( D => n13742, CK => CLK, Q => n19393, QN 
                           => n_2706);
   clk_r_REG6185_S1 : DFF_X1 port map( D => n13681, CK => CLK, Q => n19392, QN 
                           => n_2707);
   clk_r_REG5629_S1 : DFF_X1 port map( D => n13764, CK => CLK, Q => n19391, QN 
                           => n_2708);
   clk_r_REG4977_S1 : DFF_X1 port map( D => n13762, CK => CLK, Q => n19390, QN 
                           => n_2709);
   clk_r_REG4829_S1 : DFF_X1 port map( D => n13761, CK => CLK, Q => n19389, QN 
                           => n_2710);
   clk_r_REG4547_S1 : DFF_X1 port map( D => n13760, CK => CLK, Q => n19388, QN 
                           => n_2711);
   clk_r_REG4747_S1 : DFF_X1 port map( D => n13759, CK => CLK, Q => n19387, QN 
                           => n_2712);
   clk_r_REG6623_S1 : DFF_X1 port map( D => n13756, CK => CLK, Q => n19386, QN 
                           => n_2713);
   clk_r_REG4224_S1 : DFF_X1 port map( D => n13849, CK => CLK, Q => n19385, QN 
                           => n_2714);
   clk_r_REG6569_S1 : DFF_X1 port map( D => n13562, CK => CLK, Q => n19384, QN 
                           => n_2715);
   clk_r_REG4308_S1 : DFF_X1 port map( D => n13560, CK => CLK, Q => n19383, QN 
                           => n_2716);
   clk_r_REG5906_S1 : DFF_X1 port map( D => n13793, CK => CLK, Q => n19382, QN 
                           => n_2717);
   clk_r_REG5120_S1 : DFF_X1 port map( D => n13559, CK => CLK, Q => n19381, QN 
                           => n_2718);
   clk_r_REG5249_S1 : DFF_X1 port map( D => n13555, CK => CLK, Q => n19380, QN 
                           => n_2719);
   clk_r_REG4911_S1 : DFF_X1 port map( D => n13552, CK => CLK, Q => n19379, QN 
                           => n_2720);
   clk_r_REG5064_S1 : DFF_X1 port map( D => n13490, CK => CLK, Q => n19378, QN 
                           => n_2721);
   clk_r_REG5193_S1 : DFF_X1 port map( D => n13483, CK => CLK, Q => n19377, QN 
                           => n_2722);
   clk_r_REG6124_S1 : DFF_X1 port map( D => n13535, CK => CLK, Q => n19376, QN 
                           => n_2723);
   clk_r_REG6065_S1 : DFF_X1 port map( D => n13484, CK => CLK, Q => n19375, QN 
                           => n_2724);
   clk_r_REG5575_S1 : DFF_X1 port map( D => n13486, CK => CLK, Q => n19374, QN 
                           => n_2725);
   clk_r_REG5510_S1 : DFF_X1 port map( D => n13489, CK => CLK, Q => n19373, QN 
                           => n_2726);
   clk_r_REG5440_S1 : DFF_X1 port map( D => n13915, CK => CLK, Q => n19372, QN 
                           => n_2727);
   clk_r_REG5382_S1 : DFF_X1 port map( D => n13491, CK => CLK, Q => n19371, QN 
                           => n_2728);
   clk_r_REG5768_S1 : DFF_X1 port map( D => n13904, CK => CLK, Q => n19370, QN 
                           => n_2729);
   clk_r_REG5706_S1 : DFF_X1 port map( D => n13908, CK => CLK, Q => n19369, QN 
                           => n_2730);
   clk_r_REG6509_S1 : DFF_X1 port map( D => n13492, CK => CLK, Q => n19368, QN 
                           => n_2731);
   clk_r_REG5302_S1 : DFF_X1 port map( D => n13920, CK => CLK, Q => n19367, QN 
                           => n_2732);
   clk_r_REG6444_S1 : DFF_X1 port map( D => n13493, CK => CLK, Q => n19366, QN 
                           => n_2733);
   clk_r_REG6370_S1 : DFF_X1 port map( D => n13899, CK => CLK, Q => n19365, QN 
                           => n_2734);
   clk_r_REG5828_S1 : DFF_X1 port map( D => n13909, CK => CLK, Q => n19364, QN 
                           => n_2735);
   clk_r_REG5990_S1 : DFF_X1 port map( D => n13500, CK => CLK, Q => n19363, QN 
                           => n_2736);
   clk_r_REG6303_S1 : DFF_X1 port map( D => n13922, CK => CLK, Q => n19362, QN 
                           => n_2737);
   clk_r_REG6233_S1 : DFF_X1 port map( D => n13630, CK => CLK, Q => n19361, QN 
                           => n_2738);
   clk_r_REG6191_S1 : DFF_X1 port map( D => n13678, CK => CLK, Q => n19360, QN 
                           => n_2739);
   clk_r_REG5633_S1 : DFF_X1 port map( D => n13757, CK => CLK, Q => n19359, QN 
                           => n_2740);
   clk_r_REG4975_S1 : DFF_X1 port map( D => n13767, CK => CLK, Q => n19358, QN 
                           => n_2741);
   clk_r_REG4827_S1 : DFF_X1 port map( D => n13770, CK => CLK, Q => n19357, QN 
                           => n_2742);
   clk_r_REG4545_S1 : DFF_X1 port map( D => n13772, CK => CLK, Q => n19356, QN 
                           => n_2743);
   clk_r_REG4745_S1 : DFF_X1 port map( D => n13773, CK => CLK, Q => n19355, QN 
                           => n_2744);
   clk_r_REG6617_S1 : DFF_X1 port map( D => n13774, CK => CLK, Q => n19354, QN 
                           => n_2745);
   clk_r_REG4226_S1 : DFF_X1 port map( D => n13847, CK => CLK, Q => n19353, QN 
                           => n_2746);
   clk_r_REG6577_S1 : DFF_X1 port map( D => n13517, CK => CLK, Q => n19352, QN 
                           => n_2747);
   clk_r_REG4314_S1 : DFF_X1 port map( D => n13518, CK => CLK, Q => n19351, QN 
                           => n_2748);
   clk_r_REG5908_S1 : DFF_X1 port map( D => n13792, CK => CLK, Q => n19350, QN 
                           => n_2749);
   clk_r_REG5124_S1 : DFF_X1 port map( D => n13520, CK => CLK, Q => n19349, QN 
                           => n_2750);
   clk_r_REG5253_S1 : DFF_X1 port map( D => n13521, CK => CLK, Q => n19348, QN 
                           => n_2751);
   clk_r_REG4915_S1 : DFF_X1 port map( D => n13523, CK => CLK, Q => n19347, QN 
                           => n_2752);
   clk_r_REG5058_S1 : DFF_X1 port map( D => n13524, CK => CLK, Q => n19346, QN 
                           => n_2753);
   clk_r_REG5187_S1 : DFF_X1 port map( D => n13532, CK => CLK, Q => n19345, QN 
                           => n_2754);
   clk_r_REG6126_S1 : DFF_X1 port map( D => n13533, CK => CLK, Q => n19344, QN 
                           => n_2755);
   clk_r_REG6057_S1 : DFF_X1 port map( D => n13534, CK => CLK, Q => n19343, QN 
                           => n_2756);
   clk_r_REG5567_S1 : DFF_X1 port map( D => n13536, CK => CLK, Q => n19342, QN 
                           => n_2757);
   clk_r_REG5502_S1 : DFF_X1 port map( D => n13538, CK => CLK, Q => n19341, QN 
                           => n_2758);
   clk_r_REG5438_S1 : DFF_X1 port map( D => n13917, CK => CLK, Q => n19340, QN 
                           => n_2759);
   clk_r_REG5374_S1 : DFF_X1 port map( D => n13544, CK => CLK, Q => n19339, QN 
                           => n_2760);
   clk_r_REG5770_S1 : DFF_X1 port map( D => n13896, CK => CLK, Q => n19338, QN 
                           => n_2761);
   clk_r_REG5710_S1 : DFF_X1 port map( D => n13895, CK => CLK, Q => n19337, QN 
                           => n_2762);
   clk_r_REG6505_S1 : DFF_X1 port map( D => n13550, CK => CLK, Q => n19336, QN 
                           => n_2763);
   clk_r_REG5308_S1 : DFF_X1 port map( D => n13894, CK => CLK, Q => n19335, QN 
                           => n_2764);
   clk_r_REG6438_S1 : DFF_X1 port map( D => n13565, CK => CLK, Q => n19334, QN 
                           => n_2765);
   clk_r_REG6372_S1 : DFF_X1 port map( D => n13893, CK => CLK, Q => n19333, QN 
                           => n_2766);
   clk_r_REG5834_S1 : DFF_X1 port map( D => n13897, CK => CLK, Q => n19332, QN 
                           => n_2767);
   clk_r_REG5986_S1 : DFF_X1 port map( D => n13553, CK => CLK, Q => n19331, QN 
                           => n_2768);
   clk_r_REG6305_S1 : DFF_X1 port map( D => n13914, CK => CLK, Q => n19330, QN 
                           => n_2769);
   clk_r_REG6241_S1 : DFF_X1 port map( D => n13596, CK => CLK, Q => n19329, QN 
                           => n_2770);
   clk_r_REG6189_S1 : DFF_X1 port map( D => n13679, CK => CLK, Q => n19328, QN 
                           => n_2771);
   clk_r_REG5627_S1 : DFF_X1 port map( D => n13768, CK => CLK, Q => n19327, QN 
                           => n_2772);
   clk_r_REG4973_S1 : DFF_X1 port map( D => n13769, CK => CLK, Q => n19326, QN 
                           => n_2773);
   clk_r_REG4831_S1 : DFF_X1 port map( D => n13755, CK => CLK, Q => n19325, QN 
                           => n_2774);
   clk_r_REG4537_S1 : DFF_X1 port map( D => n13781, CK => CLK, Q => n19324, QN 
                           => n_2775);
   clk_r_REG4741_S1 : DFF_X1 port map( D => n13778, CK => CLK, Q => n19323, QN 
                           => n_2776);
   clk_r_REG6621_S1 : DFF_X1 port map( D => n13765, CK => CLK, Q => n19322, QN 
                           => n_2777);
   clk_r_REG4222_S1 : DFF_X1 port map( D => n13851, CK => CLK, Q => n19321, QN 
                           => n_2778);
   clk_r_REG6573_S1 : DFF_X1 port map( D => n13537, CK => CLK, Q => n19320, QN 
                           => n_2779);
   clk_r_REG4310_S1 : DFF_X1 port map( D => n13548, CK => CLK, Q => n19319, QN 
                           => n_2780);
   clk_r_REG5902_S1 : DFF_X1 port map( D => n13795, CK => CLK, Q => n19318, QN 
                           => n_2781);
   clk_r_REG5118_S1 : DFF_X1 port map( D => n13567, CK => CLK, Q => n19317, QN 
                           => n_2782);
   clk_r_REG5251_S1 : DFF_X1 port map( D => n13551, CK => CLK, Q => n19316, QN 
                           => n_2783);
   clk_r_REG4909_S1 : DFF_X1 port map( D => n13569, CK => CLK, Q => n19315, QN 
                           => n_2784);
   clk_r_REG5054_S1 : DFF_X1 port map( D => n13568, CK => CLK, Q => n19314, QN 
                           => n_2785);
   clk_r_REG5183_S1 : DFF_X1 port map( D => n13556, CK => CLK, Q => n19313, QN 
                           => n_2786);
   clk_r_REG6120_S1 : DFF_X1 port map( D => n13561, CK => CLK, Q => n19312, QN 
                           => n_2787);
   clk_r_REG6063_S1 : DFF_X1 port map( D => n13502, CK => CLK, Q => n19311, QN 
                           => n_2788);
   clk_r_REG5565_S1 : DFF_X1 port map( D => n13554, CK => CLK, Q => n19310, QN 
                           => n_2789);
   clk_r_REG5500_S1 : DFF_X1 port map( D => n13557, CK => CLK, Q => n19309, QN 
                           => n_2790);
   clk_r_REG5436_S1 : DFF_X1 port map( D => n13919, CK => CLK, Q => n19308, QN 
                           => n_2791);
   clk_r_REG5372_S1 : DFF_X1 port map( D => n13564, CK => CLK, Q => n19307, QN 
                           => n_2792);
   clk_r_REG5772_S1 : DFF_X1 port map( D => n13887, CK => CLK, Q => n19306, QN 
                           => n_2793);
   clk_r_REG5704_S1 : DFF_X1 port map( D => n13910, CK => CLK, Q => n19305, QN 
                           => n_2794);
   clk_r_REG6503_S1 : DFF_X1 port map( D => n13558, CK => CLK, Q => n19304, QN 
                           => n_2795);
   clk_r_REG5314_S1 : DFF_X1 port map( D => n13879, CK => CLK, Q => n19303, QN 
                           => n_2796);
   clk_r_REG6440_S1 : DFF_X1 port map( D => n13546, CK => CLK, Q => n19302, QN 
                           => n_2797);
   clk_r_REG6380_S1 : DFF_X1 port map( D => n13878, CK => CLK, Q => n19301, QN 
                           => n_2798);
   clk_r_REG5842_S1 : DFF_X1 port map( D => n13877, CK => CLK, Q => n19300, QN 
                           => n_2799);
   clk_r_REG5984_S1 : DFF_X1 port map( D => n13566, CK => CLK, Q => n19299, QN 
                           => n_2800);
   clk_r_REG6315_S1 : DFF_X1 port map( D => n13876, CK => CLK, Q => n19298, QN 
                           => n_2801);
   clk_r_REG6235_S1 : DFF_X1 port map( D => n13619, CK => CLK, Q => n19297, QN 
                           => n_2802);
   clk_r_REG6183_S1 : DFF_X1 port map( D => n13682, CK => CLK, Q => n19296, QN 
                           => n_2803);
   clk_r_REG5625_S1 : DFF_X1 port map( D => n13771, CK => CLK, Q => n19295, QN 
                           => n_2804);
   clk_r_REG4967_S1 : DFF_X1 port map( D => n13790, CK => CLK, Q => n19294, QN 
                           => n_2805);
   clk_r_REG4821_S1 : DFF_X1 port map( D => n13789, CK => CLK, Q => n19293, QN 
                           => n_2806);
   clk_r_REG4543_S1 : DFF_X1 port map( D => n13775, CK => CLK, Q => n19292, QN 
                           => n_2807);
   clk_r_REG4743_S1 : DFF_X1 port map( D => n13776, CK => CLK, Q => n19291, QN 
                           => n_2808);
   clk_r_REG6619_S1 : DFF_X1 port map( D => n13766, CK => CLK, Q => n19290, QN 
                           => n_2809);
   clk_r_REG4230_S1 : DFF_X1 port map( D => n13843, CK => CLK, Q => n19289, QN 
                           => n_2810);
   clk_r_REG6571_S1 : DFF_X1 port map( D => n13542, CK => CLK, Q => n19288, QN 
                           => n_2811);
   clk_r_REG4312_S1 : DFF_X1 port map( D => n13540, CK => CLK, Q => n19287, QN 
                           => n_2812);
   clk_r_REG5900_S1 : DFF_X1 port map( D => n13796, CK => CLK, Q => n19286, QN 
                           => n_2813);
   clk_r_REG5122_S1 : DFF_X1 port map( D => n13539, CK => CLK, Q => n19285, QN 
                           => n_2814);
   clk_r_REG5247_S1 : DFF_X1 port map( D => n13563, CK => CLK, Q => n19284, QN 
                           => n_2815);
   clk_r_REG4913_S1 : DFF_X1 port map( D => n13549, CK => CLK, Q => n19283, QN 
                           => n_2816);
   clk_r_REG5056_S1 : DFF_X1 port map( D => n13547, CK => CLK, Q => n19282, QN 
                           => n_2817);
   clk_r_REG5185_S1 : DFF_X1 port map( D => n13545, CK => CLK, Q => n19281, QN 
                           => n_2818);
   clk_r_REG6122_S1 : DFF_X1 port map( D => n13543, CK => CLK, Q => n19280, QN 
                           => n_2819);
   clk_r_REG6055_S1 : DFF_X1 port map( D => n13541, CK => CLK, Q => n19279, QN 
                           => n_2820);
   clk_r_REG5569_S1 : DFF_X1 port map( D => n13531, CK => CLK, Q => n19278, QN 
                           => n_2821);
   clk_r_REG5504_S1 : DFF_X1 port map( D => n13530, CK => CLK, Q => n19277, QN 
                           => n_2822);
   clk_r_REG5446_S1 : DFF_X1 port map( D => n13875, CK => CLK, Q => n19276, QN 
                           => n_2823);
   clk_r_REG5376_S1 : DFF_X1 port map( D => n13529, CK => CLK, Q => n19275, QN 
                           => n_2824);
   clk_r_REG5776_S1 : DFF_X1 port map( D => n13874, CK => CLK, Q => n19274, QN 
                           => n_2825);
   clk_r_REG5708_S1 : DFF_X1 port map( D => n13907, CK => CLK, Q => n19273, QN 
                           => n_2826);
   clk_r_REG6507_S1 : DFF_X1 port map( D => n13528, CK => CLK, Q => n19272, QN 
                           => n_2827);
   clk_r_REG5304_S1 : DFF_X1 port map( D => n13913, CK => CLK, Q => n19271, QN 
                           => n_2828);
   clk_r_REG6442_S1 : DFF_X1 port map( D => n13527, CK => CLK, Q => n19270, QN 
                           => n_2829);
   clk_r_REG6368_S1 : DFF_X1 port map( D => n13911, CK => CLK, Q => n19269, QN 
                           => n_2830);
   clk_r_REG5832_S1 : DFF_X1 port map( D => n13898, CK => CLK, Q => n19268, QN 
                           => n_2831);
   clk_r_REG5988_S1 : DFF_X1 port map( D => n13526, CK => CLK, Q => n19267, QN 
                           => n_2832);
   clk_r_REG6307_S1 : DFF_X1 port map( D => n13906, CK => CLK, Q => n19266, QN 
                           => n_2833);
   clk_r_REG6239_S1 : DFF_X1 port map( D => n13610, CK => CLK, Q => n19265, QN 
                           => n_2834);
   clk_r_REG6187_S1 : DFF_X1 port map( D => n13680, CK => CLK, Q => n19264, QN 
                           => n_2835);
   clk_r_REG5623_S1 : DFF_X1 port map( D => n13788, CK => CLK, Q => n19263, QN 
                           => n_2836);
   clk_r_REG4971_S1 : DFF_X1 port map( D => n13779, CK => CLK, Q => n19262, QN 
                           => n_2837);
   clk_r_REG4825_S1 : DFF_X1 port map( D => n13783, CK => CLK, Q => n19261, QN 
                           => n_2838);
   clk_r_REG4541_S1 : DFF_X1 port map( D => n13777, CK => CLK, Q => n19260, QN 
                           => n_2839);
   clk_r_REG4739_S1 : DFF_X1 port map( D => n13787, CK => CLK, Q => n19259, QN 
                           => n_2840);
   clk_r_REG6613_S1 : DFF_X1 port map( D => n13784, CK => CLK, Q => n19258, QN 
                           => n_2841);
   clk_r_REG4220_S1 : DFF_X1 port map( D => n13853, CK => CLK, Q => n19257, QN 
                           => n_2842);
   clk_r_REG6575_S1 : DFF_X1 port map( D => n13525, CK => CLK, Q => n19256, QN 
                           => n_2843);
   clk_r_REG4316_S1 : DFF_X1 port map( D => n13516, CK => CLK, Q => n19255, QN 
                           => n_2844);
   clk_r_REG5904_S1 : DFF_X1 port map( D => n13794, CK => CLK, Q => n19254, QN 
                           => n_2845);
   clk_r_REG5126_S1 : DFF_X1 port map( D => n13514, CK => CLK, Q => n19253, QN 
                           => n_2846);
   clk_r_REG5255_S1 : DFF_X1 port map( D => n13513, CK => CLK, Q => n19252, QN 
                           => n_2847);
   clk_r_REG4917_S1 : DFF_X1 port map( D => n13512, CK => CLK, Q => n19251, QN 
                           => n_2848);
   clk_r_REG5060_S1 : DFF_X1 port map( D => n13510, CK => CLK, Q => n19250, QN 
                           => n_2849);
   clk_r_REG5189_S1 : DFF_X1 port map( D => n13508, CK => CLK, Q => n19249, QN 
                           => n_2850);
   clk_r_REG6130_S1 : DFF_X1 port map( D => n13501, CK => CLK, Q => n19248, QN 
                           => n_2851);
   clk_r_REG6059_S1 : DFF_X1 port map( D => n13509, CK => CLK, Q => n19247, QN 
                           => n_2852);
   clk_r_REG5571_S1 : DFF_X1 port map( D => n13515, CK => CLK, Q => n19246, QN 
                           => n_2853);
   clk_r_REG5506_S1 : DFF_X1 port map( D => n13519, CK => CLK, Q => n19245, QN 
                           => n_2854);
   clk_r_REG5442_S1 : DFF_X1 port map( D => n13901, CK => CLK, Q => n19244, QN 
                           => n_2855);
   clk_r_REG5378_S1 : DFF_X1 port map( D => n13522, CK => CLK, Q => n19243, QN 
                           => n_2856);
   clk_r_REG5784_S1 : DFF_X1 port map( D => n13858, CK => CLK, Q => n19242, QN 
                           => n_2857);
   clk_r_REG5720_S1 : DFF_X1 port map( D => n13856, CK => CLK, Q => n19241, QN 
                           => n_2858);
   clk_r_REG6511_S1 : DFF_X1 port map( D => n13485, CK => CLK, Q => n19240, QN 
                           => n_2859);
   clk_r_REG5310_S1 : DFF_X1 port map( D => n13892, CK => CLK, Q => n19239, QN 
                           => n_2860);
   clk_r_REG6446_S1 : DFF_X1 port map( D => n13487, CK => CLK, Q => n19238, QN 
                           => n_2861);
   clk_r_REG6374_S1 : DFF_X1 port map( D => n13891, CK => CLK, Q => n19237, QN 
                           => n_2862);
   clk_r_REG5836_S1 : DFF_X1 port map( D => n13890, CK => CLK, Q => n19236, QN 
                           => n_2863);
   clk_r_REG5992_S1 : DFF_X1 port map( D => n13488, CK => CLK, Q => n19235, QN 
                           => n_2864);
   clk_r_REG6311_S1 : DFF_X1 port map( D => n13889, CK => CLK, Q => n19234, QN 
                           => n_2865);
   clk_r_REG6237_S1 : DFF_X1 port map( D => n13615, CK => CLK, Q => n19233, QN 
                           => n_2866);
   clk_r_REG6193_S1 : DFF_X1 port map( D => n13677, CK => CLK, Q => n19232, QN 
                           => n_2867);
   clk_r_REG5631_S1 : DFF_X1 port map( D => n13763, CK => CLK, Q => n19231, QN 
                           => n_2868);
   clk_r_REG4969_S1 : DFF_X1 port map( D => n13785, CK => CLK, Q => n19230, QN 
                           => n_2869);
   clk_r_REG4823_S1 : DFF_X1 port map( D => n13786, CK => CLK, Q => n19229, QN 
                           => n_2870);
   clk_r_REG4539_S1 : DFF_X1 port map( D => n13780, CK => CLK, Q => n19228, QN 
                           => n_2871);
   clk_r_REG4749_S1 : DFF_X1 port map( D => n13758, CK => CLK, Q => n19227, QN 
                           => n_2872);
   clk_r_REG6615_S1 : DFF_X1 port map( D => n13782, CK => CLK, Q => n19226, QN 
                           => n_2873);
   clk_r_REG4228_S1 : DFF_X1 port map( D => n13845, CK => CLK, Q => n19225, QN 
                           => n_2874);
   clk_r_REG6579_S1 : DFF_X1 port map( D => n13494, CK => CLK, Q => n19224, QN 
                           => n_2875);
   clk_r_REG4318_S1 : DFF_X1 port map( D => n13495, CK => CLK, Q => n19223, QN 
                           => n_2876);
   clk_r_REG5910_S1 : DFF_X1 port map( D => n13791, CK => CLK, Q => n19222, QN 
                           => n_2877);
   clk_r_REG5128_S1 : DFF_X1 port map( D => n13496, CK => CLK, Q => n19221, QN 
                           => n_2878);
   clk_r_REG5257_S1 : DFF_X1 port map( D => n13497, CK => CLK, Q => n19220, QN 
                           => n_2879);
   clk_r_REG4919_S1 : DFF_X1 port map( D => n13498, CK => CLK, Q => n19219, QN 
                           => n_2880);
   clk_r_REG5062_S1 : DFF_X1 port map( D => n13499, CK => CLK, Q => n19218, QN 
                           => n_2881);
   clk_r_REG5191_S1 : DFF_X1 port map( D => n13503, CK => CLK, Q => n19217, QN 
                           => n_2882);
   clk_r_REG6128_S1 : DFF_X1 port map( D => n13504, CK => CLK, Q => n19216, QN 
                           => n_2883);
   clk_r_REG6061_S1 : DFF_X1 port map( D => n13505, CK => CLK, Q => n19215, QN 
                           => n_2884);
   clk_r_REG5573_S1 : DFF_X1 port map( D => n13506, CK => CLK, Q => n19214, QN 
                           => n_2885);
   clk_r_REG5508_S1 : DFF_X1 port map( D => n13507, CK => CLK, Q => n19213, QN 
                           => n_2886);
   clk_r_REG5444_S1 : DFF_X1 port map( D => n13888, CK => CLK, Q => n19212, QN 
                           => n_2887);
   clk_r_REG5380_S1 : DFF_X1 port map( D => n13511, CK => CLK, Q => n19211, QN 
                           => n_2888);
   clk_r_REG5774_S1 : DFF_X1 port map( D => n13886, CK => CLK, Q => n19210, QN 
                           => n_2889);
   clk_r_REG5714_S1 : DFF_X1 port map( D => n13867, CK => CLK, Q => n19209, QN 
                           => n_2890);
   clk_r_REG6497_S1 : DFF_X1 port map( D => n13580, CK => CLK, Q => n19208, QN 
                           => n_2891);
   clk_r_REG5264_S1 : DFF_X1 port map( D => n14415, CK => CLK, Q => n19207, QN 
                           => n_2892);
   clk_r_REG6424_S1 : DFF_X1 port map( D => n13620, CK => CLK, Q => n19206, QN 
                           => n_2893);
   clk_r_REG6338_S1 : DFF_X1 port map( D => n14391, CK => CLK, Q => n19205, QN 
                           => n_2894);
   clk_r_REG5786_S1 : DFF_X1 port map( D => n14394, CK => CLK, Q => n19204, QN 
                           => n_2895);
   clk_r_REG5970_S1 : DFF_X1 port map( D => n13621, CK => CLK, Q => n19203, QN 
                           => n_2896);
   clk_r_REG6277_S1 : DFF_X1 port map( D => n14364, CK => CLK, Q => n19202, QN 
                           => n_2897);
   clk_r_REG6231_S1 : DFF_X1 port map( D => n13638, CK => CLK, Q => n19201, QN 
                           => n_2898);
   clk_r_REG6135_S1 : DFF_X1 port map( D => n14475, CK => CLK, Q => n19200, QN 
                           => n_2899);
   clk_r_REG5605_S1 : DFF_X1 port map( D => n14532, CK => CLK, Q => n19199, QN 
                           => n_2900);
   clk_r_REG4943_S1 : DFF_X1 port map( D => n14585, CK => CLK, Q => n19198, QN 
                           => n_2901);
   clk_r_REG4803_S1 : DFF_X1 port map( D => n14531, CK => CLK, Q => n19197, QN 
                           => n_2902);
   clk_r_REG4513_S1 : DFF_X1 port map( D => n14542, CK => CLK, Q => n19196, QN 
                           => n_2903);
   clk_r_REG4715_S1 : DFF_X1 port map( D => n14559, CK => CLK, Q => n19195, QN 
                           => n_2904);
   clk_r_REG6585_S1 : DFF_X1 port map( D => n14596, CK => CLK, Q => n19194, QN 
                           => n_2905);
   clk_r_REG4176_S1 : DFF_X1 port map( D => n14609, CK => CLK, Q => n19193, QN 
                           => n_2906);
   clk_r_REG6533_S1 : DFF_X1 port map( D => n13978, CK => CLK, Q => n19192, QN 
                           => n_2907);
   clk_r_REG4264_S1 : DFF_X1 port map( D => n14037, CK => CLK, Q => n19191, QN 
                           => n_2908);
   clk_r_REG5878_S1 : DFF_X1 port map( D => n14036, CK => CLK, Q => n19190, QN 
                           => n_2909);
   clk_r_REG5076_S1 : DFF_X1 port map( D => n14028, CK => CLK, Q => n19189, QN 
                           => n_2910);
   clk_r_REG5207_S1 : DFF_X1 port map( D => n14013, CK => CLK, Q => n19188, QN 
                           => n_2911);
   clk_r_REG4869_S1 : DFF_X1 port map( D => n14006, CK => CLK, Q => n19187, QN 
                           => n_2912);
   clk_r_REG5020_S1 : DFF_X1 port map( D => n13961, CK => CLK, Q => n19186, QN 
                           => n_2913);
   clk_r_REG5153_S1 : DFF_X1 port map( D => n13996, CK => CLK, Q => n19185, QN 
                           => n_2914);
   clk_r_REG6074_S1 : DFF_X1 port map( D => n14266, CK => CLK, Q => n19184, QN 
                           => n_2915);
   clk_r_REG6021_S1 : DFF_X1 port map( D => n14217, CK => CLK, Q => n19183, QN 
                           => n_2916);
   clk_r_REG5529_S1 : DFF_X1 port map( D => n13962, CK => CLK, Q => n19182, QN 
                           => n_2917);
   clk_r_REG5464_S1 : DFF_X1 port map( D => n13963, CK => CLK, Q => n19181, QN 
                           => n_2918);
   clk_r_REG5428_S1 : DFF_X1 port map( D => n13964, CK => CLK, Q => n19180, QN 
                           => n_2919);
   clk_r_REG5332_S1 : DFF_X1 port map( D => n14188, CK => CLK, Q => n19179, QN 
                           => n_2920);
   clk_r_REG5758_S1 : DFF_X1 port map( D => n13965, CK => CLK, Q => n19178, QN 
                           => n_2921);
   clk_r_REG5694_S1 : DFF_X1 port map( D => n13966, CK => CLK, Q => n19177, QN 
                           => n_2922);
   clk_r_REG6465_S1 : DFF_X1 port map( D => n14238, CK => CLK, Q => n19176, QN 
                           => n_2923);
   clk_r_REG5298_S1 : DFF_X1 port map( D => n14038, CK => CLK, Q => n19175, QN 
                           => n_2924);
   clk_r_REG6406_S1 : DFF_X1 port map( D => n14052, CK => CLK, Q => n19174, QN 
                           => n_2925);
   clk_r_REG6354_S1 : DFF_X1 port map( D => n14090, CK => CLK, Q => n19173, QN 
                           => n_2926);
   clk_r_REG5814_S1 : DFF_X1 port map( D => n14082, CK => CLK, Q => n19172, QN 
                           => n_2927);
   clk_r_REG5942_S1 : DFF_X1 port map( D => n14121, CK => CLK, Q => n19171, QN 
                           => n_2928);
   clk_r_REG6287_S1 : DFF_X1 port map( D => n14103, CK => CLK, Q => n19170, QN 
                           => n_2929);
   clk_r_REG6229_S1 : DFF_X1 port map( D => n14150, CK => CLK, Q => n19169, QN 
                           => n_2930);
   clk_r_REG6133_S1 : DFF_X1 port map( D => n14477, CK => CLK, Q => n19168, QN 
                           => n_2931);
   clk_r_REG5603_S1 : DFF_X1 port map( D => n14535, CK => CLK, Q => n19167, QN 
                           => n_2932);
   clk_r_REG3936_S1 : DFF_X1 port map( D => n14595, CK => CLK, Q => n19166, QN 
                           => n_2933);
   clk_r_REG4801_S1 : DFF_X1 port map( D => n14537, CK => CLK, Q => n19165, QN 
                           => n_2934);
   clk_r_REG4519_S1 : DFF_X1 port map( D => n14539, CK => CLK, Q => n19164, QN 
                           => n_2935);
   clk_r_REG4713_S1 : DFF_X1 port map( D => n14561, CK => CLK, Q => n19163, QN 
                           => n_2936);
   clk_r_REG6599_S1 : DFF_X1 port map( D => n14569, CK => CLK, Q => n19162, QN 
                           => n_2937);
   clk_r_REG4178_S1 : DFF_X1 port map( D => n14607, CK => CLK, Q => n19161, QN 
                           => n_2938);
   clk_r_REG6531_S1 : DFF_X1 port map( D => n13979, CK => CLK, Q => n19160, QN 
                           => n_2939);
   clk_r_REG4272_S1 : DFF_X1 port map( D => n13988, CK => CLK, Q => n19159, QN 
                           => n_2940);
   clk_r_REG5880_S1 : DFF_X1 port map( D => n14035, CK => CLK, Q => n19158, QN 
                           => n_2941);
   clk_r_REG5078_S1 : DFF_X1 port map( D => n14027, CK => CLK, Q => n19157, QN 
                           => n_2942);
   clk_r_REG5209_S1 : DFF_X1 port map( D => n14012, CK => CLK, Q => n19156, QN 
                           => n_2943);
   clk_r_REG4871_S1 : DFF_X1 port map( D => n14005, CK => CLK, Q => n19155, QN 
                           => n_2944);
   clk_r_REG5018_S1 : DFF_X1 port map( D => n13968, CK => CLK, Q => n19154, QN 
                           => n_2945);
   clk_r_REG5155_S1 : DFF_X1 port map( D => n13995, CK => CLK, Q => n19153, QN 
                           => n_2946);
   clk_r_REG6076_S1 : DFF_X1 port map( D => n14264, CK => CLK, Q => n19152, QN 
                           => n_2947);
   clk_r_REG6023_S1 : DFF_X1 port map( D => n14216, CK => CLK, Q => n19151, QN 
                           => n_2948);
   clk_r_REG5527_S1 : DFF_X1 port map( D => n13969, CK => CLK, Q => n19150, QN 
                           => n_2949);
   clk_r_REG5462_S1 : DFF_X1 port map( D => n13970, CK => CLK, Q => n19149, QN 
                           => n_2950);
   clk_r_REG5426_S1 : DFF_X1 port map( D => n13971, CK => CLK, Q => n19148, QN 
                           => n_2951);
   clk_r_REG5334_S1 : DFF_X1 port map( D => n14187, CK => CLK, Q => n19147, QN 
                           => n_2952);
   clk_r_REG5756_S1 : DFF_X1 port map( D => n13972, CK => CLK, Q => n19146, QN 
                           => n_2953);
   clk_r_REG5692_S1 : DFF_X1 port map( D => n13973, CK => CLK, Q => n19145, QN 
                           => n_2954);
   clk_r_REG6483_S1 : DFF_X1 port map( D => n14237, CK => CLK, Q => n19144, QN 
                           => n_2955);
   clk_r_REG5262_S1 : DFF_X1 port map( D => n14416, CK => CLK, Q => n19143, QN 
                           => n_2956);
   clk_r_REG6422_S1 : DFF_X1 port map( D => n14053, CK => CLK, Q => n19142, QN 
                           => n_2957);
   clk_r_REG6340_S1 : DFF_X1 port map( D => n14390, CK => CLK, Q => n19141, QN 
                           => n_2958);
   clk_r_REG3676_S1 : DFF_X1 port map( D => n14396, CK => CLK, Q => n19140, QN 
                           => n_2959);
   clk_r_REG5964_S1 : DFF_X1 port map( D => n14123, CK => CLK, Q => n19139, QN 
                           => n_2960);
   clk_r_REG6275_S1 : DFF_X1 port map( D => n14368, CK => CLK, Q => n19138, QN 
                           => n_2961);
   clk_r_REG6227_S1 : DFF_X1 port map( D => n14151, CK => CLK, Q => n19137, QN 
                           => n_2962);
   clk_r_REG6149_S1 : DFF_X1 port map( D => n14461, CK => CLK, Q => n19136, QN 
                           => n_2963);
   clk_r_REG3715_S1 : DFF_X1 port map( D => n14592, CK => CLK, Q => n19135, QN 
                           => n_2964);
   clk_r_REG4937_S1 : DFF_X1 port map( D => n14593, CK => CLK, Q => n19134, QN 
                           => n_2965);
   clk_r_REG4791_S1 : DFF_X1 port map( D => n14564, CK => CLK, Q => n19133, QN 
                           => n_2966);
   clk_r_REG4509_S1 : DFF_X1 port map( D => n14563, CK => CLK, Q => n19132, QN 
                           => n_2967);
   clk_r_REG4711_S1 : DFF_X1 port map( D => n14562, CK => CLK, Q => n19131, QN 
                           => n_2968);
   clk_r_REG6583_S1 : DFF_X1 port map( D => n14602, CK => CLK, Q => n19130, QN 
                           => n_2969);
   clk_r_REG4182_S1 : DFF_X1 port map( D => n14590, CK => CLK, Q => n19129, QN 
                           => n_2970);
   clk_r_REG6529_S1 : DFF_X1 port map( D => n13980, CK => CLK, Q => n19128, QN 
                           => n_2971);
   clk_r_REG4270_S1 : DFF_X1 port map( D => n13989, CK => CLK, Q => n19127, QN 
                           => n_2972);
   clk_r_REG5882_S1 : DFF_X1 port map( D => n14034, CK => CLK, Q => n19126, QN 
                           => n_2973);
   clk_r_REG5080_S1 : DFF_X1 port map( D => n14026, CK => CLK, Q => n19125, QN 
                           => n_2974);
   clk_r_REG5211_S1 : DFF_X1 port map( D => n14011, CK => CLK, Q => n19124, QN 
                           => n_2975);
   clk_r_REG4873_S1 : DFF_X1 port map( D => n14004, CK => CLK, Q => n19123, QN 
                           => n_2976);
   clk_r_REG5016_S1 : DFF_X1 port map( D => n13977, CK => CLK, Q => n19122, QN 
                           => n_2977);
   clk_r_REG5157_S1 : DFF_X1 port map( D => n13994, CK => CLK, Q => n19121, QN 
                           => n_2978);
   clk_r_REG6078_S1 : DFF_X1 port map( D => n14263, CK => CLK, Q => n19120, QN 
                           => n_2979);
   clk_r_REG6025_S1 : DFF_X1 port map( D => n14215, CK => CLK, Q => n19119, QN 
                           => n_2980);
   clk_r_REG5525_S1 : DFF_X1 port map( D => n13981, CK => CLK, Q => n19118, QN 
                           => n_2981);
   clk_r_REG5460_S1 : DFF_X1 port map( D => n13982, CK => CLK, Q => n19117, QN 
                           => n_2982);
   clk_r_REG5424_S1 : DFF_X1 port map( D => n13983, CK => CLK, Q => n19116, QN 
                           => n_2983);
   clk_r_REG5336_S1 : DFF_X1 port map( D => n14186, CK => CLK, Q => n19115, QN 
                           => n_2984);
   clk_r_REG5754_S1 : DFF_X1 port map( D => n13984, CK => CLK, Q => n19114, QN 
                           => n_2985);
   clk_r_REG5690_S1 : DFF_X1 port map( D => n13985, CK => CLK, Q => n19113, QN 
                           => n_2986);
   clk_r_REG6467_S1 : DFF_X1 port map( D => n14236, CK => CLK, Q => n19112, QN 
                           => n_2987);
   clk_r_REG5296_S1 : DFF_X1 port map( D => n14039, CK => CLK, Q => n19111, QN 
                           => n_2988);
   clk_r_REG6404_S1 : DFF_X1 port map( D => n14054, CK => CLK, Q => n19110, QN 
                           => n_2989);
   clk_r_REG6352_S1 : DFF_X1 port map( D => n14091, CK => CLK, Q => n19109, QN 
                           => n_2990);
   clk_r_REG5812_S1 : DFF_X1 port map( D => n14084, CK => CLK, Q => n19108, QN 
                           => n_2991);
   clk_r_REG5954_S1 : DFF_X1 port map( D => n14108, CK => CLK, Q => n19107, QN 
                           => n_2992);
   clk_r_REG6297_S1 : DFF_X1 port map( D => n14096, CK => CLK, Q => n19106, QN 
                           => n_2993);
   clk_r_REG6207_S1 : DFF_X1 port map( D => n14152, CK => CLK, Q => n19105, QN 
                           => n_2994);
   clk_r_REG3589_S1 : DFF_X1 port map( D => n14480, CK => CLK, Q => n19104, QN 
                           => n_2995);
   clk_r_REG5601_S1 : DFF_X1 port map( D => n14536, CK => CLK, Q => n19103, QN 
                           => n_2996);
   clk_r_REG4939_S1 : DFF_X1 port map( D => n14589, CK => CLK, Q => n19102, QN 
                           => n_2997);
   clk_r_REG4799_S1 : DFF_X1 port map( D => n14538, CK => CLK, Q => n19101, QN 
                           => n_2998);
   clk_r_REG4517_S1 : DFF_X1 port map( D => n14540, CK => CLK, Q => n19100, QN 
                           => n_2999);
   clk_r_REG4729_S1 : DFF_X1 port map( D => n14546, CK => CLK, Q => n19099, QN 
                           => n_3000);
   clk_r_REG6603_S1 : DFF_X1 port map( D => n14565, CK => CLK, Q => n19098, QN 
                           => n_3001);
   clk_r_REG4184_S1 : DFF_X1 port map( D => n14587, CK => CLK, Q => n19097, QN 
                           => n_3002);
   clk_r_REG6525_S1 : DFF_X1 port map( D => n14030, CK => CLK, Q => n19096, QN 
                           => n_3003);
   clk_r_REG4266_S1 : DFF_X1 port map( D => n14029, CK => CLK, Q => n19095, QN 
                           => n_3004);
   clk_r_REG5884_S1 : DFF_X1 port map( D => n14033, CK => CLK, Q => n19094, QN 
                           => n_3005);
   clk_r_REG5082_S1 : DFF_X1 port map( D => n14025, CK => CLK, Q => n19093, QN 
                           => n_3006);
   clk_r_REG5205_S1 : DFF_X1 port map( D => n14021, CK => CLK, Q => n19092, QN 
                           => n_3007);
   clk_r_REG4867_S1 : DFF_X1 port map( D => n14020, CK => CLK, Q => n19091, QN 
                           => n_3008);
   clk_r_REG5012_S1 : DFF_X1 port map( D => n14019, CK => CLK, Q => n19090, QN 
                           => n_3009);
   clk_r_REG5149_S1 : DFF_X1 port map( D => n14018, CK => CLK, Q => n19089, QN 
                           => n_3010);
   clk_r_REG6086_S1 : DFF_X1 port map( D => n14250, CK => CLK, Q => n19088, QN 
                           => n_3011);
   clk_r_REG6027_S1 : DFF_X1 port map( D => n14214, CK => CLK, Q => n19087, QN 
                           => n_3012);
   clk_r_REG5523_S1 : DFF_X1 port map( D => n14017, CK => CLK, Q => n19086, QN 
                           => n_3013);
   clk_r_REG5458_S1 : DFF_X1 port map( D => n14016, CK => CLK, Q => n19085, QN 
                           => n_3014);
   clk_r_REG5422_S1 : DFF_X1 port map( D => n14015, CK => CLK, Q => n19084, QN 
                           => n_3015);
   clk_r_REG5338_S1 : DFF_X1 port map( D => n14185, CK => CLK, Q => n19083, QN 
                           => n_3016);
   clk_r_REG5752_S1 : DFF_X1 port map( D => n14014, CK => CLK, Q => n19082, QN 
                           => n_3017);
   clk_r_REG5688_S1 : DFF_X1 port map( D => n14007, CK => CLK, Q => n19081, QN 
                           => n_3018);
   clk_r_REG6469_S1 : DFF_X1 port map( D => n14235, CK => CLK, Q => n19080, QN 
                           => n_3019);
   clk_r_REG5294_S1 : DFF_X1 port map( D => n14040, CK => CLK, Q => n19079, QN 
                           => n_3020);
   clk_r_REG6402_S1 : DFF_X1 port map( D => n14055, CK => CLK, Q => n19078, QN 
                           => n_3021);
   clk_r_REG6350_S1 : DFF_X1 port map( D => n14092, CK => CLK, Q => n19077, QN 
                           => n_3022);
   clk_r_REG5824_S1 : DFF_X1 port map( D => n14071, CK => CLK, Q => n19076, QN 
                           => n_3023);
   clk_r_REG5952_S1 : DFF_X1 port map( D => n14109, CK => CLK, Q => n19075, QN 
                           => n_3024);
   clk_r_REG6295_S1 : DFF_X1 port map( D => n14098, CK => CLK, Q => n19074, QN 
                           => n_3025);
   clk_r_REG6205_S1 : DFF_X1 port map( D => n14153, CK => CLK, Q => n19073, QN 
                           => n_3026);
   clk_r_REG6143_S1 : DFF_X1 port map( D => n14467, CK => CLK, Q => n19072, QN 
                           => n_3027);
   clk_r_REG5595_S1 : DFF_X1 port map( D => n14555, CK => CLK, Q => n19071, QN 
                           => n_3028);
   clk_r_REG4941_S1 : DFF_X1 port map( D => n14586, CK => CLK, Q => n19070, QN 
                           => n_3029);
   clk_r_REG4793_S1 : DFF_X1 port map( D => n14560, CK => CLK, Q => n19069, QN 
                           => n_3030);
   clk_r_REG4507_S1 : DFF_X1 port map( D => n14566, CK => CLK, Q => n19068, QN 
                           => n_3031);
   clk_r_REG4709_S1 : DFF_X1 port map( D => n14567, CK => CLK, Q => n19067, QN 
                           => n_3032);
   clk_r_REG6601_S1 : DFF_X1 port map( D => n14568, CK => CLK, Q => n19066, QN 
                           => n_3033);
   clk_r_REG4170_S1 : DFF_X1 port map( D => n14617, CK => CLK, Q => n19065, QN 
                           => n_3034);
   clk_r_REG6527_S1 : DFF_X1 port map( D => n14000, CK => CLK, Q => n19064, QN 
                           => n_3035);
   clk_r_REG4268_S1 : DFF_X1 port map( D => n13999, CK => CLK, Q => n19063, QN 
                           => n_3036);
   clk_r_REG5886_S1 : DFF_X1 port map( D => n14032, CK => CLK, Q => n19062, QN 
                           => n_3037);
   clk_r_REG5084_S1 : DFF_X1 port map( D => n14024, CK => CLK, Q => n19061, QN 
                           => n_3038);
   clk_r_REG5213_S1 : DFF_X1 port map( D => n14010, CK => CLK, Q => n19060, QN 
                           => n_3039);
   clk_r_REG4875_S1 : DFF_X1 port map( D => n14003, CK => CLK, Q => n19059, QN 
                           => n_3040);
   clk_r_REG5014_S1 : DFF_X1 port map( D => n13998, CK => CLK, Q => n19058, QN 
                           => n_3041);
   clk_r_REG5151_S1 : DFF_X1 port map( D => n13997, CK => CLK, Q => n19057, QN 
                           => n_3042);
   clk_r_REG6080_S1 : DFF_X1 port map( D => n14257, CK => CLK, Q => n19056, QN 
                           => n_3043);
   clk_r_REG6029_S1 : DFF_X1 port map( D => n14213, CK => CLK, Q => n19055, QN 
                           => n_3044);
   clk_r_REG5531_S1 : DFF_X1 port map( D => n13960, CK => CLK, Q => n19054, QN 
                           => n_3045);
   clk_r_REG5470_S1 : DFF_X1 port map( D => n13948, CK => CLK, Q => n19053, QN 
                           => n_3046);
   clk_r_REG5434_S1 : DFF_X1 port map( D => n13945, CK => CLK, Q => n19052, QN 
                           => n_3047);
   clk_r_REG5340_S1 : DFF_X1 port map( D => n14184, CK => CLK, Q => n19051, QN 
                           => n_3048);
   clk_r_REG5760_S1 : DFF_X1 port map( D => n13957, CK => CLK, Q => n19050, QN 
                           => n_3049);
   clk_r_REG5700_S1 : DFF_X1 port map( D => n13952, CK => CLK, Q => n19049, QN 
                           => n_3050);
   clk_r_REG6471_S1 : DFF_X1 port map( D => n14234, CK => CLK, Q => n19048, QN 
                           => n_3051);
   clk_r_REG5292_S1 : DFF_X1 port map( D => n14041, CK => CLK, Q => n19047, QN 
                           => n_3052);
   clk_r_REG6400_S1 : DFF_X1 port map( D => n14056, CK => CLK, Q => n19046, QN 
                           => n_3053);
   clk_r_REG6364_S1 : DFF_X1 port map( D => n14085, CK => CLK, Q => n19045, QN 
                           => n_3054);
   clk_r_REG5822_S1 : DFF_X1 port map( D => n14072, CK => CLK, Q => n19044, QN 
                           => n_3055);
   clk_r_REG5950_S1 : DFF_X1 port map( D => n14110, CK => CLK, Q => n19043, QN 
                           => n_3056);
   clk_r_REG6293_S1 : DFF_X1 port map( D => n14099, CK => CLK, Q => n19042, QN 
                           => n_3057);
   clk_r_REG6203_S1 : DFF_X1 port map( D => n14154, CK => CLK, Q => n19041, QN 
                           => n_3058);
   clk_r_REG6161_S1 : DFF_X1 port map( D => n14374, CK => CLK, Q => n19040, QN 
                           => n_3059);
   clk_r_REG5607_S1 : DFF_X1 port map( D => n14524, CK => CLK, Q => n19039, QN 
                           => n_3060);
   clk_r_REG4945_S1 : DFF_X1 port map( D => n14578, CK => CLK, Q => n19038, QN 
                           => n_3061);
   clk_r_REG4807_S1 : DFF_X1 port map( D => n14528, CK => CLK, Q => n19037, QN 
                           => n_3062);
   clk_r_REG4523_S1 : DFF_X1 port map( D => n14523, CK => CLK, Q => n19036, QN 
                           => n_3063);
   clk_r_REG4727_S1 : DFF_X1 port map( D => n14548, CK => CLK, Q => n19035, QN 
                           => n_3064);
   clk_r_REG6597_S1 : DFF_X1 port map( D => n14570, CK => CLK, Q => n19034, QN 
                           => n_3065);
   clk_r_REG4128_S1 : DFF_X1 port map( D => n14620, CK => CLK, Q => n19033, QN 
                           => n_3066);
   clk_r_REG6539_S1 : DFF_X1 port map( D => n13974, CK => CLK, Q => n19032, QN 
                           => n_3067);
   clk_r_REG4290_S1 : DFF_X1 port map( D => n13990, CK => CLK, Q => n19031, QN 
                           => n_3068);
   clk_r_REG5852_S1 : DFF_X1 port map( D => n14304, CK => CLK, Q => n19030, QN 
                           => n_3069);
   clk_r_REG5086_S1 : DFF_X1 port map( D => n14023, CK => CLK, Q => n19029, QN 
                           => n_3070);
   clk_r_REG5215_S1 : DFF_X1 port map( D => n14009, CK => CLK, Q => n19028, QN 
                           => n_3071);
   clk_r_REG4877_S1 : DFF_X1 port map( D => n14002, CK => CLK, Q => n19027, QN 
                           => n_3072);
   clk_r_REG5024_S1 : DFF_X1 port map( D => n13944, CK => CLK, Q => n19026, QN 
                           => n_3073);
   clk_r_REG5159_S1 : DFF_X1 port map( D => n13993, CK => CLK, Q => n19025, QN 
                           => n_3074);
   clk_r_REG6070_S1 : DFF_X1 port map( D => n14284, CK => CLK, Q => n19024, QN 
                           => n_3075);
   clk_r_REG6031_S1 : DFF_X1 port map( D => n14212, CK => CLK, Q => n19023, QN 
                           => n_3076);
   clk_r_REG5535_S1 : DFF_X1 port map( D => n13958, CK => CLK, Q => n19022, QN 
                           => n_3077);
   clk_r_REG5468_S1 : DFF_X1 port map( D => n13949, CK => CLK, Q => n19021, QN 
                           => n_3078);
   clk_r_REG5432_S1 : DFF_X1 port map( D => n13946, CK => CLK, Q => n19020, QN 
                           => n_3079);
   clk_r_REG5342_S1 : DFF_X1 port map( D => n14183, CK => CLK, Q => n19019, QN 
                           => n_3080);
   clk_r_REG5764_S1 : DFF_X1 port map( D => n13955, CK => CLK, Q => n19018, QN 
                           => n_3081);
   clk_r_REG5698_S1 : DFF_X1 port map( D => n13953, CK => CLK, Q => n19017, QN 
                           => n_3082);
   clk_r_REG6487_S1 : DFF_X1 port map( D => n13967, CK => CLK, Q => n19016, QN 
                           => n_3083);
   clk_r_REG5260_S1 : DFF_X1 port map( D => n14418, CK => CLK, Q => n19015, QN 
                           => n_3084);
   clk_r_REG6420_S1 : DFF_X1 port map( D => n14057, CK => CLK, Q => n19014, QN 
                           => n_3085);
   clk_r_REG6342_S1 : DFF_X1 port map( D => n14385, CK => CLK, Q => n19013, QN 
                           => n_3086);
   clk_r_REG5790_S1 : DFF_X1 port map( D => n14392, CK => CLK, Q => n19012, QN 
                           => n_3087);
   clk_r_REG5968_S1 : DFF_X1 port map( D => n14111, CK => CLK, Q => n19011, QN 
                           => n_3088);
   clk_r_REG6263_S1 : DFF_X1 port map( D => n14383, CK => CLK, Q => n19010, QN 
                           => n_3089);
   clk_r_REG6201_S1 : DFF_X1 port map( D => n14155, CK => CLK, Q => n19009, QN 
                           => n_3090);
   clk_r_REG6151_S1 : DFF_X1 port map( D => n14459, CK => CLK, Q => n19008, QN 
                           => n_3091);
   clk_r_REG5609_S1 : DFF_X1 port map( D => n14522, CK => CLK, Q => n19007, QN 
                           => n_3092);
   clk_r_REG4947_S1 : DFF_X1 port map( D => n14577, CK => CLK, Q => n19006, QN 
                           => n_3093);
   clk_r_REG4809_S1 : DFF_X1 port map( D => n14527, CK => CLK, Q => n19005, QN 
                           => n_3094);
   clk_r_REG4525_S1 : DFF_X1 port map( D => n14519, CK => CLK, Q => n19004, QN 
                           => n_3095);
   clk_r_REG4725_S1 : DFF_X1 port map( D => n14550, CK => CLK, Q => n19003, QN 
                           => n_3096);
   clk_r_REG6595_S1 : DFF_X1 port map( D => n14571, CK => CLK, Q => n19002, QN 
                           => n_3097);
   clk_r_REG4180_S1 : DFF_X1 port map( D => n14598, CK => CLK, Q => n19001, QN 
                           => n_3098);
   clk_r_REG6537_S1 : DFF_X1 port map( D => n13975, CK => CLK, Q => n19000, QN 
                           => n_3099);
   clk_r_REG4276_S1 : DFF_X1 port map( D => n13986, CK => CLK, Q => n18999, QN 
                           => n_3100);
   clk_r_REG5888_S1 : DFF_X1 port map( D => n14031, CK => CLK, Q => n18998, QN 
                           => n_3101);
   clk_r_REG5088_S1 : DFF_X1 port map( D => n14022, CK => CLK, Q => n18997, QN 
                           => n_3102);
   clk_r_REG5217_S1 : DFF_X1 port map( D => n14008, CK => CLK, Q => n18996, QN 
                           => n_3103);
   clk_r_REG4879_S1 : DFF_X1 port map( D => n14001, CK => CLK, Q => n18995, QN 
                           => n_3104);
   clk_r_REG5022_S1 : DFF_X1 port map( D => n13947, CK => CLK, Q => n18994, QN 
                           => n_3105);
   clk_r_REG5161_S1 : DFF_X1 port map( D => n13992, CK => CLK, Q => n18993, QN 
                           => n_3106);
   clk_r_REG3609_S1 : DFF_X1 port map( D => n14286, CK => CLK, Q => n18992, QN 
                           => n_3107);
   clk_r_REG6033_S1 : DFF_X1 port map( D => n14209, CK => CLK, Q => n18991, QN 
                           => n_3108);
   clk_r_REG5533_S1 : DFF_X1 port map( D => n13959, CK => CLK, Q => n18990, QN 
                           => n_3109);
   clk_r_REG5466_S1 : DFF_X1 port map( D => n13950, CK => CLK, Q => n18989, QN 
                           => n_3110);
   clk_r_REG5430_S1 : DFF_X1 port map( D => n13951, CK => CLK, Q => n18988, QN 
                           => n_3111);
   clk_r_REG5322_S1 : DFF_X1 port map( D => n14200, CK => CLK, Q => n18987, QN 
                           => n_3112);
   clk_r_REG5762_S1 : DFF_X1 port map( D => n13956, CK => CLK, Q => n18986, QN 
                           => n_3113);
   clk_r_REG5696_S1 : DFF_X1 port map( D => n13954, CK => CLK, Q => n18985, QN 
                           => n_3114);
   clk_r_REG6485_S1 : DFF_X1 port map( D => n14233, CK => CLK, Q => n18984, QN 
                           => n_3115);
   clk_r_REG5284_S1 : DFF_X1 port map( D => n14182, CK => CLK, Q => n18983, QN 
                           => n_3116);
   clk_r_REG6398_S1 : DFF_X1 port map( D => n14058, CK => CLK, Q => n18982, QN 
                           => n_3117);
   clk_r_REG6362_S1 : DFF_X1 port map( D => n14086, CK => CLK, Q => n18981, QN 
                           => n_3118);
   clk_r_REG5820_S1 : DFF_X1 port map( D => n14077, CK => CLK, Q => n18980, QN 
                           => n_3119);
   clk_r_REG5948_S1 : DFF_X1 port map( D => n14112, CK => CLK, Q => n18979, QN 
                           => n_3120);
   clk_r_REG6291_S1 : DFF_X1 port map( D => n14100, CK => CLK, Q => n18978, QN 
                           => n_3121);
   clk_r_REG6199_S1 : DFF_X1 port map( D => n14156, CK => CLK, Q => n18977, QN 
                           => n_3122);
   clk_r_REG6139_S1 : DFF_X1 port map( D => n14471, CK => CLK, Q => n18976, QN 
                           => n_3123);
   clk_r_REG5593_S1 : DFF_X1 port map( D => n14557, CK => CLK, Q => n18975, QN 
                           => n_3124);
   clk_r_REG4949_S1 : DFF_X1 port map( D => n14575, CK => CLK, Q => n18974, QN 
                           => n_3125);
   clk_r_REG4805_S1 : DFF_X1 port map( D => n14530, CK => CLK, Q => n18973, QN 
                           => n_3126);
   clk_r_REG4515_S1 : DFF_X1 port map( D => n14541, CK => CLK, Q => n18972, QN 
                           => n_3127);
   clk_r_REG4717_S1 : DFF_X1 port map( D => n14558, CK => CLK, Q => n18971, QN 
                           => n_3128);
   clk_r_REG3518_S1 : DFF_X1 port map( D => n14611, CK => CLK, Q => n18970, QN 
                           => n_3129);
   clk_r_REG4172_S1 : DFF_X1 port map( D => n14615, CK => CLK, Q => n18969, QN 
                           => n_3130);
   clk_r_REG6535_S1 : DFF_X1 port map( D => n13976, CK => CLK, Q => n18968, QN 
                           => n_3131);
   clk_r_REG4274_S1 : DFF_X1 port map( D => n13987, CK => CLK, Q => n18967, QN 
                           => n_3132);
   clk_r_REG5890_S1 : DFF_X1 port map( D => n13991, CK => CLK, Q => n18966, QN 
                           => n_3133);
   clk_r_REG3855_S1 : DFF_X1 port map( D => n14211, CK => CLK, Q => n18965, QN 
                           => n_3134);
   clk_r_REG3784_S1 : DFF_X1 port map( D => n14288, CK => CLK, Q => n18964, QN 
                           => n_3135);
   clk_r_REG3949_S1 : DFF_X1 port map( D => n14281, CK => CLK, Q => n18963, QN 
                           => n_3136);
   clk_r_REG3880_S1 : DFF_X1 port map( D => n14283, CK => CLK, Q => n18962, QN 
                           => n_3137);
   clk_r_REG5139_S1 : DFF_X1 port map( D => n14278, CK => CLK, Q => n18961, QN 
                           => n_3138);
   clk_r_REG6072_S1 : DFF_X1 port map( D => n14279, CK => CLK, Q => n18960, QN 
                           => n_3139);
   clk_r_REG6011_S1 : DFF_X1 port map( D => n14260, CK => CLK, Q => n18959, QN 
                           => n_3140);
   clk_r_REG3732_S1 : DFF_X1 port map( D => n14277, CK => CLK, Q => n18958, QN 
                           => n_3141);
   clk_r_REG3739_S1 : DFF_X1 port map( D => n14275, CK => CLK, Q => n18957, QN 
                           => n_3142);
   clk_r_REG5412_S1 : DFF_X1 port map( D => n14273, CK => CLK, Q => n18956, QN 
                           => n_3143);
   clk_r_REG3753_S1 : DFF_X1 port map( D => n14272, CK => CLK, Q => n18955, QN 
                           => n_3144);
   clk_r_REG5742_S1 : DFF_X1 port map( D => n14270, CK => CLK, Q => n18954, QN 
                           => n_3145);
   clk_r_REG5678_S1 : DFF_X1 port map( D => n14269, CK => CLK, Q => n18953, QN 
                           => n_3146);
   clk_r_REG3545_S1 : DFF_X1 port map( D => n14268, CK => CLK, Q => n18952, QN 
                           => n_3147);
   clk_r_REG5280_S1 : DFF_X1 port map( D => n14243, CK => CLK, Q => n18951, QN 
                           => n_3148);
   clk_r_REG3553_S1 : DFF_X1 port map( D => n14242, CK => CLK, Q => n18950, QN 
                           => n_3149);
   clk_r_REG6344_S1 : DFF_X1 port map( D => n14240, CK => CLK, Q => n18949, QN 
                           => n_3150);
   clk_r_REG5804_S1 : DFF_X1 port map( D => n14239, CK => CLK, Q => n18948, QN 
                           => n_3151);
   clk_r_REG5936_S1 : DFF_X1 port map( D => n14232, CK => CLK, Q => n18947, QN 
                           => n_3152);
   clk_r_REG6279_S1 : DFF_X1 port map( D => n14231, CK => CLK, Q => n18946, QN 
                           => n_3153);
   clk_r_REG6223_S1 : DFF_X1 port map( D => n14230, CK => CLK, Q => n18945, QN 
                           => n_3154);
   clk_r_REG6165_S1 : DFF_X1 port map( D => n14354, CK => CLK, Q => n18944, QN 
                           => n_3155);
   clk_r_REG5611_S1 : DFF_X1 port map( D => n14521, CK => CLK, Q => n18943, QN 
                           => n_3156);
   clk_r_REG4955_S1 : DFF_X1 port map( D => n14529, CK => CLK, Q => n18942, QN 
                           => n_3157);
   clk_r_REG4811_S1 : DFF_X1 port map( D => n14525, CK => CLK, Q => n18941, QN 
                           => n_3158);
   clk_r_REG4527_S1 : DFF_X1 port map( D => n14518, CK => CLK, Q => n18940, QN 
                           => n_3159);
   clk_r_REG4723_S1 : DFF_X1 port map( D => n14551, CK => CLK, Q => n18939, QN 
                           => n_3160);
   clk_r_REG6593_S1 : DFF_X1 port map( D => n14576, CK => CLK, Q => n18938, QN 
                           => n_3161);
   clk_r_REG4186_S1 : DFF_X1 port map( D => n14584, CK => CLK, Q => n18937, QN 
                           => n_3162);
   clk_r_REG3531_S1 : DFF_X1 port map( D => n14221, CK => CLK, Q => n18936, QN 
                           => n_3163);
   clk_r_REG4061_S1 : DFF_X1 port map( D => n14219, CK => CLK, Q => n18935, QN 
                           => n_3164);
   clk_r_REG5870_S1 : DFF_X1 port map( D => n14208, CK => CLK, Q => n18934, QN 
                           => n_3165);
   clk_r_REG5068_S1 : DFF_X1 port map( D => n14207, CK => CLK, Q => n18933, QN 
                           => n_3166);
   clk_r_REG5197_S1 : DFF_X1 port map( D => n14206, CK => CLK, Q => n18932, QN 
                           => n_3167);
   clk_r_REG4859_S1 : DFF_X1 port map( D => n14205, CK => CLK, Q => n18931, QN 
                           => n_3168);
   clk_r_REG5004_S1 : DFF_X1 port map( D => n14203, CK => CLK, Q => n18930, QN 
                           => n_3169);
   clk_r_REG5141_S1 : DFF_X1 port map( D => n14202, CK => CLK, Q => n18929, QN 
                           => n_3170);
   clk_r_REG6082_S1 : DFF_X1 port map( D => n14252, CK => CLK, Q => n18928, QN 
                           => n_3171);
   clk_r_REG6013_S1 : DFF_X1 port map( D => n14228, CK => CLK, Q => n18927, QN 
                           => n_3172);
   clk_r_REG5515_S1 : DFF_X1 port map( D => n14201, CK => CLK, Q => n18926, QN 
                           => n_3173);
   clk_r_REG5450_S1 : DFF_X1 port map( D => n14192, CK => CLK, Q => n18925, QN 
                           => n_3174);
   clk_r_REG5414_S1 : DFF_X1 port map( D => n14191, CK => CLK, Q => n18924, QN 
                           => n_3175);
   clk_r_REG5324_S1 : DFF_X1 port map( D => n14199, CK => CLK, Q => n18923, QN 
                           => n_3176);
   clk_r_REG5744_S1 : DFF_X1 port map( D => n14190, CK => CLK, Q => n18922, QN 
                           => n_3177);
   clk_r_REG5680_S1 : DFF_X1 port map( D => n14189, CK => CLK, Q => n18921, QN 
                           => n_3178);
   clk_r_REG6455_S1 : DFF_X1 port map( D => n14259, CK => CLK, Q => n18920, QN 
                           => n_3179);
   clk_r_REG5288_S1 : DFF_X1 port map( D => n14180, CK => CLK, Q => n18919, QN 
                           => n_3180);
   clk_r_REG6396_S1 : DFF_X1 port map( D => n14060, CK => CLK, Q => n18918, QN 
                           => n_3181);
   clk_r_REG6360_S1 : DFF_X1 port map( D => n14087, CK => CLK, Q => n18917, QN 
                           => n_3182);
   clk_r_REG5818_S1 : DFF_X1 port map( D => n14078, CK => CLK, Q => n18916, QN 
                           => n_3183);
   clk_r_REG5946_S1 : DFF_X1 port map( D => n14113, CK => CLK, Q => n18915, QN 
                           => n_3184);
   clk_r_REG6289_S1 : DFF_X1 port map( D => n14101, CK => CLK, Q => n18914, QN 
                           => n_3185);
   clk_r_REG6197_S1 : DFF_X1 port map( D => n14157, CK => CLK, Q => n18913, QN 
                           => n_3186);
   clk_r_REG6141_S1 : DFF_X1 port map( D => n14469, CK => CLK, Q => n18912, QN 
                           => n_3187);
   clk_r_REG5613_S1 : DFF_X1 port map( D => n14520, CK => CLK, Q => n18911, QN 
                           => n_3188);
   clk_r_REG4957_S1 : DFF_X1 port map( D => n14526, CK => CLK, Q => n18910, QN 
                           => n_3189);
   clk_r_REG3979_S1 : DFF_X1 port map( D => n14600, CK => CLK, Q => n18909, QN 
                           => n_3190);
   clk_r_REG4048_S1 : DFF_X1 port map( D => n14605, CK => CLK, Q => n18908, QN 
                           => n_3191);
   clk_r_REG3993_S1 : DFF_X1 port map( D => n14574, CK => CLK, Q => n18907, QN 
                           => n_3192);
   clk_r_REG6591_S1 : DFF_X1 port map( D => n14579, CK => CLK, Q => n18906, QN 
                           => n_3193);
   clk_r_REG4188_S1 : DFF_X1 port map( D => n14572, CK => CLK, Q => n18905, QN 
                           => n_3194);
   clk_r_REG6523_S1 : DFF_X1 port map( D => n14042, CK => CLK, Q => n18904, QN 
                           => n_3195);
   clk_r_REG4262_S1 : DFF_X1 port map( D => n14043, CK => CLK, Q => n18903, QN 
                           => n_3196);
   clk_r_REG5876_S1 : DFF_X1 port map( D => n14044, CK => CLK, Q => n18902, QN 
                           => n_3197);
   clk_r_REG5074_S1 : DFF_X1 port map( D => n14045, CK => CLK, Q => n18901, QN 
                           => n_3198);
   clk_r_REG5203_S1 : DFF_X1 port map( D => n14046, CK => CLK, Q => n18900, QN 
                           => n_3199);
   clk_r_REG4865_S1 : DFF_X1 port map( D => n14047, CK => CLK, Q => n18899, QN 
                           => n_3200);
   clk_r_REG5010_S1 : DFF_X1 port map( D => n14048, CK => CLK, Q => n18898, QN 
                           => n_3201);
   clk_r_REG5147_S1 : DFF_X1 port map( D => n14050, CK => CLK, Q => n18897, QN 
                           => n_3202);
   clk_r_REG6084_S1 : DFF_X1 port map( D => n14251, CK => CLK, Q => n18896, QN 
                           => n_3203);
   clk_r_REG6015_S1 : DFF_X1 port map( D => n14227, CK => CLK, Q => n18895, QN 
                           => n_3204);
   clk_r_REG5521_S1 : DFF_X1 port map( D => n14051, CK => CLK, Q => n18894, QN 
                           => n_3205);
   clk_r_REG5456_S1 : DFF_X1 port map( D => n14061, CK => CLK, Q => n18893, QN 
                           => n_3206);
   clk_r_REG5420_S1 : DFF_X1 port map( D => n14062, CK => CLK, Q => n18892, QN 
                           => n_3207);
   clk_r_REG5326_S1 : DFF_X1 port map( D => n14198, CK => CLK, Q => n18891, QN 
                           => n_3208);
   clk_r_REG5750_S1 : DFF_X1 port map( D => n14063, CK => CLK, Q => n18890, QN 
                           => n_3209);
   clk_r_REG5684_S1 : DFF_X1 port map( D => n14064, CK => CLK, Q => n18889, QN 
                           => n_3210);
   clk_r_REG6457_S1 : DFF_X1 port map( D => n14258, CK => CLK, Q => n18888, QN 
                           => n_3211);
   clk_r_REG5286_S1 : DFF_X1 port map( D => n14181, CK => CLK, Q => n18887, QN 
                           => n_3212);
   clk_r_REG6394_S1 : DFF_X1 port map( D => n14068, CK => CLK, Q => n18886, QN 
                           => n_3213);
   clk_r_REG6358_S1 : DFF_X1 port map( D => n14088, CK => CLK, Q => n18885, QN 
                           => n_3214);
   clk_r_REG5810_S1 : DFF_X1 port map( D => n14102, CK => CLK, Q => n18884, QN 
                           => n_3215);
   clk_r_REG5944_S1 : DFF_X1 port map( D => n14115, CK => CLK, Q => n18883, QN 
                           => n_3216);
   clk_r_REG6285_S1 : DFF_X1 port map( D => n14104, CK => CLK, Q => n18882, QN 
                           => n_3217);
   clk_r_REG6225_S1 : DFF_X1 port map( D => n14158, CK => CLK, Q => n18881, QN 
                           => n_3218);
   clk_r_REG6163_S1 : DFF_X1 port map( D => n14362, CK => CLK, Q => n18880, QN 
                           => n_3219);
   clk_r_REG5599_S1 : DFF_X1 port map( D => n14545, CK => CLK, Q => n18879, QN 
                           => n_3220);
   clk_r_REG4953_S1 : DFF_X1 port map( D => n14544, CK => CLK, Q => n18878, QN 
                           => n_3221);
   clk_r_REG4797_S1 : DFF_X1 port map( D => n14543, CK => CLK, Q => n18877, QN 
                           => n_3222);
   clk_r_REG4521_S1 : DFF_X1 port map( D => n14534, CK => CLK, Q => n18876, QN 
                           => n_3223);
   clk_r_REG4719_S1 : DFF_X1 port map( D => n14556, CK => CLK, Q => n18875, QN 
                           => n_3224);
   clk_r_REG6589_S1 : DFF_X1 port map( D => n14581, CK => CLK, Q => n18874, QN 
                           => n_3225);
   clk_r_REG4190_S1 : DFF_X1 port map( D => n14533, CK => CLK, Q => n18873, QN 
                           => n_3226);
   clk_r_REG6551_S1 : DFF_X1 port map( D => n14119, CK => CLK, Q => n18872, QN 
                           => n_3227);
   clk_r_REG4288_S1 : DFF_X1 port map( D => n14120, CK => CLK, Q => n18871, QN 
                           => n_3228);
   clk_r_REG5860_S1 : DFF_X1 port map( D => n14300, CK => CLK, Q => n18870, QN 
                           => n_3229);
   clk_r_REG5098_S1 : DFF_X1 port map( D => n14130, CK => CLK, Q => n18869, QN 
                           => n_3230);
   clk_r_REG5227_S1 : DFF_X1 port map( D => n14132, CK => CLK, Q => n18868, QN 
                           => n_3231);
   clk_r_REG4861_S1 : DFF_X1 port map( D => n14133, CK => CLK, Q => n18867, QN 
                           => n_3232);
   clk_r_REG5006_S1 : DFF_X1 port map( D => n14139, CK => CLK, Q => n18866, QN 
                           => n_3233);
   clk_r_REG5143_S1 : DFF_X1 port map( D => n14140, CK => CLK, Q => n18865, QN 
                           => n_3234);
   clk_r_REG6088_S1 : DFF_X1 port map( D => n14249, CK => CLK, Q => n18864, QN 
                           => n_3235);
   clk_r_REG6017_S1 : DFF_X1 port map( D => n14226, CK => CLK, Q => n18863, QN 
                           => n_3236);
   clk_r_REG5517_S1 : DFF_X1 port map( D => n14141, CK => CLK, Q => n18862, QN 
                           => n_3237);
   clk_r_REG5452_S1 : DFF_X1 port map( D => n14142, CK => CLK, Q => n18861, QN 
                           => n_3238);
   clk_r_REG5416_S1 : DFF_X1 port map( D => n14143, CK => CLK, Q => n18860, QN 
                           => n_3239);
   clk_r_REG5328_S1 : DFF_X1 port map( D => n14197, CK => CLK, Q => n18859, QN 
                           => n_3240);
   clk_r_REG5746_S1 : DFF_X1 port map( D => n14144, CK => CLK, Q => n18858, QN 
                           => n_3241);
   clk_r_REG5682_S1 : DFF_X1 port map( D => n14148, CK => CLK, Q => n18857, QN 
                           => n_3242);
   clk_r_REG6459_S1 : DFF_X1 port map( D => n14256, CK => CLK, Q => n18856, QN 
                           => n_3243);
   clk_r_REG5282_S1 : DFF_X1 port map( D => n14204, CK => CLK, Q => n18855, QN 
                           => n_3244);
   clk_r_REG6390_S1 : DFF_X1 port map( D => n14149, CK => CLK, Q => n18854, QN 
                           => n_3245);
   clk_r_REG6346_S1 : DFF_X1 port map( D => n14159, CK => CLK, Q => n18853, QN 
                           => n_3246);
   clk_r_REG5806_S1 : DFF_X1 port map( D => n14160, CK => CLK, Q => n18852, QN 
                           => n_3247);
   clk_r_REG5938_S1 : DFF_X1 port map( D => n14161, CK => CLK, Q => n18851, QN 
                           => n_3248);
   clk_r_REG6281_S1 : DFF_X1 port map( D => n14162, CK => CLK, Q => n18850, QN 
                           => n_3249);
   clk_r_REG3580_S1 : DFF_X1 port map( D => n14164, CK => CLK, Q => n18849, QN 
                           => n_3250);
   clk_r_REG6137_S1 : DFF_X1 port map( D => n14473, CK => CLK, Q => n18848, QN 
                           => n_3251);
   clk_r_REG5637_S1 : DFF_X1 port map( D => n14504, CK => CLK, Q => n18847, QN 
                           => n_3252);
   clk_r_REG4979_S1 : DFF_X1 port map( D => n14506, CK => CLK, Q => n18846, QN 
                           => n_3253);
   clk_r_REG4833_S1 : DFF_X1 port map( D => n14512, CK => CLK, Q => n18845, QN 
                           => n_3254);
   clk_r_REG4551_S1 : DFF_X1 port map( D => n14498, CK => CLK, Q => n18844, QN 
                           => n_3255);
   clk_r_REG4753_S1 : DFF_X1 port map( D => n14501, CK => CLK, Q => n18843, QN 
                           => n_3256);
   clk_r_REG6627_S1 : DFF_X1 port map( D => n14495, CK => CLK, Q => n18842, QN 
                           => n_3257);
   clk_r_REG4202_S1 : DFF_X1 port map( D => n14496, CK => CLK, Q => n18841, QN 
                           => n_3258);
   clk_r_REG6519_S1 : DFF_X1 port map( D => n14177, CK => CLK, Q => n18840, QN 
                           => n_3259);
   clk_r_REG4258_S1 : DFF_X1 port map( D => n14178, CK => CLK, Q => n18839, QN 
                           => n_3260);
   clk_r_REG5872_S1 : DFF_X1 port map( D => n14179, CK => CLK, Q => n18838, QN 
                           => n_3261);
   clk_r_REG5070_S1 : DFF_X1 port map( D => n14176, CK => CLK, Q => n18837, QN 
                           => n_3262);
   clk_r_REG5199_S1 : DFF_X1 port map( D => n14175, CK => CLK, Q => n18836, QN 
                           => n_3263);
   clk_r_REG4889_S1 : DFF_X1 port map( D => n14174, CK => CLK, Q => n18835, QN 
                           => n_3264);
   clk_r_REG5034_S1 : DFF_X1 port map( D => n14172, CK => CLK, Q => n18834, QN 
                           => n_3265);
   clk_r_REG5163_S1 : DFF_X1 port map( D => n14170, CK => CLK, Q => n18833, QN 
                           => n_3266);
   clk_r_REG6100_S1 : DFF_X1 port map( D => n14248, CK => CLK, Q => n18832, QN 
                           => n_3267);
   clk_r_REG6035_S1 : DFF_X1 port map( D => n14225, CK => CLK, Q => n18831, QN 
                           => n_3268);
   clk_r_REG5545_S1 : DFF_X1 port map( D => n14168, CK => CLK, Q => n18830, QN 
                           => n_3269);
   clk_r_REG5480_S1 : DFF_X1 port map( D => n14166, CK => CLK, Q => n18829, QN 
                           => n_3270);
   clk_r_REG5392_S1 : DFF_X1 port map( D => n14413, CK => CLK, Q => n18828, QN 
                           => n_3271);
   clk_r_REG5352_S1 : DFF_X1 port map( D => n14196, CK => CLK, Q => n18827, QN 
                           => n_3272);
   clk_r_REG5724_S1 : DFF_X1 port map( D => n14352, CK => CLK, Q => n18826, QN 
                           => n_3273);
   clk_r_REG5666_S1 : DFF_X1 port map( D => n14347, CK => CLK, Q => n18825, QN 
                           => n_3274);
   clk_r_REG6461_S1 : DFF_X1 port map( D => n14255, CK => CLK, Q => n18824, QN 
                           => n_3275);
   clk_r_REG5278_S1 : DFF_X1 port map( D => n14265, CK => CLK, Q => n18823, QN 
                           => n_3276);
   clk_r_REG6392_S1 : DFF_X1 port map( D => n14138, CK => CLK, Q => n18822, QN 
                           => n_3277);
   clk_r_REG6348_S1 : DFF_X1 port map( D => n14137, CK => CLK, Q => n18821, QN 
                           => n_3278);
   clk_r_REG5808_S1 : DFF_X1 port map( D => n14136, CK => CLK, Q => n18820, QN 
                           => n_3279);
   clk_r_REG5940_S1 : DFF_X1 port map( D => n14135, CK => CLK, Q => n18819, QN 
                           => n_3280);
   clk_r_REG6283_S1 : DFF_X1 port map( D => n14134, CK => CLK, Q => n18818, QN 
                           => n_3281);
   clk_r_REG6213_S1 : DFF_X1 port map( D => n14145, CK => CLK, Q => n18817, QN 
                           => n_3282);
   clk_r_REG6147_S1 : DFF_X1 port map( D => n14463, CK => CLK, Q => n18816, QN 
                           => n_3283);
   clk_r_REG5635_S1 : DFF_X1 port map( D => n14514, CK => CLK, Q => n18815, QN 
                           => n_3284);
   clk_r_REG4981_S1 : DFF_X1 port map( D => n14497, CK => CLK, Q => n18814, QN 
                           => n_3285);
   clk_r_REG4835_S1 : DFF_X1 port map( D => n14507, CK => CLK, Q => n18813, QN 
                           => n_3286);
   clk_r_REG4549_S1 : DFF_X1 port map( D => n14517, CK => CLK, Q => n18812, QN 
                           => n_3287);
   clk_r_REG4751_S1 : DFF_X1 port map( D => n14503, CK => CLK, Q => n18811, QN 
                           => n_3288);
   clk_r_REG6625_S1 : DFF_X1 port map( D => n14509, CK => CLK, Q => n18810, QN 
                           => n_3289);
   clk_r_REG4200_S1 : DFF_X1 port map( D => n14500, CK => CLK, Q => n18809, QN 
                           => n_3290);
   clk_r_REG6549_S1 : DFF_X1 port map( D => n14128, CK => CLK, Q => n18808, QN 
                           => n_3291);
   clk_r_REG4286_S1 : DFF_X1 port map( D => n14126, CK => CLK, Q => n18807, QN 
                           => n_3292);
   clk_r_REG5866_S1 : DFF_X1 port map( D => n14297, CK => CLK, Q => n18806, QN 
                           => n_3293);
   clk_r_REG5100_S1 : DFF_X1 port map( D => n14124, CK => CLK, Q => n18805, QN 
                           => n_3294);
   clk_r_REG5229_S1 : DFF_X1 port map( D => n14118, CK => CLK, Q => n18804, QN 
                           => n_3295);
   clk_r_REG4891_S1 : DFF_X1 port map( D => n14117, CK => CLK, Q => n18803, QN 
                           => n_3296);
   clk_r_REG5036_S1 : DFF_X1 port map( D => n14114, CK => CLK, Q => n18802, QN 
                           => n_3297);
   clk_r_REG5165_S1 : DFF_X1 port map( D => n14107, CK => CLK, Q => n18801, QN 
                           => n_3298);
   clk_r_REG6102_S1 : DFF_X1 port map( D => n14246, CK => CLK, Q => n18800, QN 
                           => n_3299);
   clk_r_REG6037_S1 : DFF_X1 port map( D => n14223, CK => CLK, Q => n18799, QN 
                           => n_3300);
   clk_r_REG5547_S1 : DFF_X1 port map( D => n14106, CK => CLK, Q => n18798, QN 
                           => n_3301);
   clk_r_REG5482_S1 : DFF_X1 port map( D => n14105, CK => CLK, Q => n18797, QN 
                           => n_3302);
   clk_r_REG5394_S1 : DFF_X1 port map( D => n14360, CK => CLK, Q => n18796, QN 
                           => n_3303);
   clk_r_REG5354_S1 : DFF_X1 port map( D => n14194, CK => CLK, Q => n18795, QN 
                           => n_3304);
   clk_r_REG3694_S1 : DFF_X1 port map( D => n14356, CK => CLK, Q => n18794, QN 
                           => n_3305);
   clk_r_REG5674_S1 : DFF_X1 port map( D => n14336, CK => CLK, Q => n18793, QN 
                           => n_3306);
   clk_r_REG6481_S1 : DFF_X1 port map( D => n14254, CK => CLK, Q => n18792, QN 
                           => n_3307);
   clk_r_REG5272_S1 : DFF_X1 port map( D => n14386, CK => CLK, Q => n18791, QN 
                           => n_3308);
   clk_r_REG6418_S1 : DFF_X1 port map( D => n14094, CK => CLK, Q => n18790, QN 
                           => n_3309);
   clk_r_REG6334_S1 : DFF_X1 port map( D => n14398, CK => CLK, Q => n18789, QN 
                           => n_3310);
   clk_r_REG5788_S1 : DFF_X1 port map( D => n14393, CK => CLK, Q => n18788, QN 
                           => n_3311);
   clk_r_REG5966_S1 : DFF_X1 port map( D => n14116, CK => CLK, Q => n18787, QN 
                           => n_3312);
   clk_r_REG6261_S1 : DFF_X1 port map( D => n14389, CK => CLK, Q => n18786, QN 
                           => n_3313);
   clk_r_REG6211_S1 : DFF_X1 port map( D => n14146, CK => CLK, Q => n18785, QN 
                           => n_3314);
   clk_r_REG6145_S1 : DFF_X1 port map( D => n14465, CK => CLK, Q => n18784, QN 
                           => n_3315);
   clk_r_REG5597_S1 : DFF_X1 port map( D => n14547, CK => CLK, Q => n18783, QN 
                           => n_3316);
   clk_r_REG4951_S1 : DFF_X1 port map( D => n14549, CK => CLK, Q => n18782, QN 
                           => n_3317);
   clk_r_REG4795_S1 : DFF_X1 port map( D => n14552, CK => CLK, Q => n18781, QN 
                           => n_3318);
   clk_r_REG4511_S1 : DFF_X1 port map( D => n14553, CK => CLK, Q => n18780, QN 
                           => n_3319);
   clk_r_REG4721_S1 : DFF_X1 port map( D => n14554, CK => CLK, Q => n18779, QN 
                           => n_3320);
   clk_r_REG6587_S1 : DFF_X1 port map( D => n14582, CK => CLK, Q => n18778, QN 
                           => n_3321);
   clk_r_REG4174_S1 : DFF_X1 port map( D => n14613, CK => CLK, Q => n18777, QN 
                           => n_3322);
   clk_r_REG6521_S1 : DFF_X1 port map( D => n14083, CK => CLK, Q => n18776, QN 
                           => n_3323);
   clk_r_REG4260_S1 : DFF_X1 port map( D => n14081, CK => CLK, Q => n18775, QN 
                           => n_3324);
   clk_r_REG5874_S1 : DFF_X1 port map( D => n14079, CK => CLK, Q => n18774, QN 
                           => n_3325);
   clk_r_REG5072_S1 : DFF_X1 port map( D => n14076, CK => CLK, Q => n18773, QN 
                           => n_3326);
   clk_r_REG5201_S1 : DFF_X1 port map( D => n14075, CK => CLK, Q => n18772, QN 
                           => n_3327);
   clk_r_REG4863_S1 : DFF_X1 port map( D => n14074, CK => CLK, Q => n18771, QN 
                           => n_3328);
   clk_r_REG5008_S1 : DFF_X1 port map( D => n14073, CK => CLK, Q => n18770, QN 
                           => n_3329);
   clk_r_REG5145_S1 : DFF_X1 port map( D => n14070, CK => CLK, Q => n18769, QN 
                           => n_3330);
   clk_r_REG6090_S1 : DFF_X1 port map( D => n14245, CK => CLK, Q => n18768, QN 
                           => n_3331);
   clk_r_REG6019_S1 : DFF_X1 port map( D => n14222, CK => CLK, Q => n18767, QN 
                           => n_3332);
   clk_r_REG5519_S1 : DFF_X1 port map( D => n14069, CK => CLK, Q => n18766, QN 
                           => n_3333);
   clk_r_REG5454_S1 : DFF_X1 port map( D => n14067, CK => CLK, Q => n18765, QN 
                           => n_3334);
   clk_r_REG5418_S1 : DFF_X1 port map( D => n14066, CK => CLK, Q => n18764, QN 
                           => n_3335);
   clk_r_REG5330_S1 : DFF_X1 port map( D => n14193, CK => CLK, Q => n18763, QN 
                           => n_3336);
   clk_r_REG5748_S1 : DFF_X1 port map( D => n14065, CK => CLK, Q => n18762, QN 
                           => n_3337);
   clk_r_REG5686_S1 : DFF_X1 port map( D => n14059, CK => CLK, Q => n18761, QN 
                           => n_3338);
   clk_r_REG6463_S1 : DFF_X1 port map( D => n14244, CK => CLK, Q => n18760, QN 
                           => n_3339);
   clk_r_REG5290_S1 : DFF_X1 port map( D => n14097, CK => CLK, Q => n18759, QN 
                           => n_3340);
   clk_r_REG6408_S1 : DFF_X1 port map( D => n14049, CK => CLK, Q => n18758, QN 
                           => n_3341);
   clk_r_REG6356_S1 : DFF_X1 port map( D => n14089, CK => CLK, Q => n18757, QN 
                           => n_3342);
   clk_r_REG5816_S1 : DFF_X1 port map( D => n14080, CK => CLK, Q => n18756, QN 
                           => n_3343);
   clk_r_REG3628_S1 : DFF_X1 port map( D => n14262, CK => CLK, Q => n18755, QN 
                           => n_3344);
   clk_r_REG6299_S1 : DFF_X1 port map( D => n14095, CK => CLK, Q => n18754, QN 
                           => n_3345);
   clk_r_REG6209_S1 : DFF_X1 port map( D => n14147, CK => CLK, Q => n18753, QN 
                           => n_3346);
   clk_r_REG6153_S1 : DFF_X1 port map( D => n14309, CK => CLK, Q => n18752, QN 
                           => n_3347);
   clk_r_REG5615_S1 : DFF_X1 port map( D => n14494, CK => CLK, Q => n18751, QN 
                           => n_3348);
   clk_r_REG4959_S1 : DFF_X1 port map( D => n14483, CK => CLK, Q => n18750, QN 
                           => n_3349);
   clk_r_REG4813_S1 : DFF_X1 port map( D => n14481, CK => CLK, Q => n18749, QN 
                           => n_3350);
   clk_r_REG4529_S1 : DFF_X1 port map( D => n14492, CK => CLK, Q => n18748, QN 
                           => n_3351);
   clk_r_REG4731_S1 : DFF_X1 port map( D => n14486, CK => CLK, Q => n18747, QN 
                           => n_3352);
   clk_r_REG6605_S1 : DFF_X1 port map( D => n14487, CK => CLK, Q => n18746, QN 
                           => n_3353);
   clk_r_REG4192_S1 : DFF_X1 port map( D => n14482, CK => CLK, Q => n18745, QN 
                           => n_3354);
   clk_r_REG6541_S1 : DFF_X1 port map( D => n13939, CK => CLK, Q => n18744, QN 
                           => n_3355);
   clk_r_REG4278_S1 : DFF_X1 port map( D => n13941, CK => CLK, Q => n18743, QN 
                           => n_3356);
   clk_r_REG5892_S1 : DFF_X1 port map( D => n13931, CK => CLK, Q => n18742, QN 
                           => n_3357);
   clk_r_REG5090_S1 : DFF_X1 port map( D => n13929, CK => CLK, Q => n18741, QN 
                           => n_3358);
   clk_r_REG5219_S1 : DFF_X1 port map( D => n13928, CK => CLK, Q => n18740, QN 
                           => n_3359);
   clk_r_REG4881_S1 : DFF_X1 port map( D => n13936, CK => CLK, Q => n18739, QN 
                           => n_3360);
   clk_r_REG5026_S1 : DFF_X1 port map( D => n13943, CK => CLK, Q => n18738, QN 
                           => n_3361);
   clk_r_REG3830_S1 : DFF_X1 port map( D => n14485, CK => CLK, Q => n18737, QN 
                           => n_3362);
   clk_r_REG6092_S1 : DFF_X1 port map( D => n13935, CK => CLK, Q => n18736, QN 
                           => n_3363);
   clk_r_REG3616_S1 : DFF_X1 port map( D => n14491, CK => CLK, Q => n18735, QN 
                           => n_3364);
   clk_r_REG5537_S1 : DFF_X1 port map( D => n13937, CK => CLK, Q => n18734, QN 
                           => n_3365);
   clk_r_REG5472_S1 : DFF_X1 port map( D => n13925, CK => CLK, Q => n18733, QN 
                           => n_3366);
   clk_r_REG3746_S1 : DFF_X1 port map( D => n14489, CK => CLK, Q => n18732, QN 
                           => n_3367);
   clk_r_REG5344_S1 : DFF_X1 port map( D => n13930, CK => CLK, Q => n18731, QN 
                           => n_3368);
   clk_r_REG5766_S1 : DFF_X1 port map( D => n13932, CK => CLK, Q => n18730, QN 
                           => n_3369);
   clk_r_REG5702_S1 : DFF_X1 port map( D => n13940, CK => CLK, Q => n18729, QN 
                           => n_3370);
   clk_r_REG6473_S1 : DFF_X1 port map( D => n13933, CK => CLK, Q => n18728, QN 
                           => n_3371);
   clk_r_REG5300_S1 : DFF_X1 port map( D => n13927, CK => CLK, Q => n18727, QN 
                           => n_3372);
   clk_r_REG6410_S1 : DFF_X1 port map( D => n13934, CK => CLK, Q => n18726, QN 
                           => n_3373);
   clk_r_REG6366_S1 : DFF_X1 port map( D => n13924, CK => CLK, Q => n18725, QN 
                           => n_3374);
   clk_r_REG5826_S1 : DFF_X1 port map( D => n13938, CK => CLK, Q => n18724, QN 
                           => n_3375);
   clk_r_REG5956_S1 : DFF_X1 port map( D => n13926, CK => CLK, Q => n18723, QN 
                           => n_3376);
   clk_r_REG6301_S1 : DFF_X1 port map( D => n13923, CK => CLK, Q => n18722, QN 
                           => n_3377);
   clk_r_REG6215_S1 : DFF_X1 port map( D => n13942, CK => CLK, Q => n18721, QN 
                           => n_3378);
   clk_r_REG6157_S1 : DFF_X1 port map( D => n14292, CK => CLK, Q => n18720, QN 
                           => n_3379);
   clk_r_REG5617_S1 : DFF_X1 port map( D => n14453, CK => CLK, Q => n18719, QN 
                           => n_3380);
   clk_r_REG4965_S1 : DFF_X1 port map( D => n14425, CK => CLK, Q => n18718, QN 
                           => n_3381);
   clk_r_REG4815_S1 : DFF_X1 port map( D => n14444, CK => CLK, Q => n18717, QN 
                           => n_3382);
   clk_r_REG4533_S1 : DFF_X1 port map( D => n14447, CK => CLK, Q => n18716, QN 
                           => n_3383);
   clk_r_REG4733_S1 : DFF_X1 port map( D => n14457, CK => CLK, Q => n18715, QN 
                           => n_3384);
   clk_r_REG6607_S1 : DFF_X1 port map( D => n14452, CK => CLK, Q => n18714, QN 
                           => n_3385);
   clk_r_REG4194_S1 : DFF_X1 port map( D => n14441, CK => CLK, Q => n18713, QN 
                           => n_3386);
   clk_r_REG6547_S1 : DFF_X1 port map( D => n13805, CK => CLK, Q => n18712, QN 
                           => n_3387);
   clk_r_REG4282_S1 : DFF_X1 port map( D => n13808, CK => CLK, Q => n18711, QN 
                           => n_3388);
   clk_r_REG5898_S1 : DFF_X1 port map( D => n13800, CK => CLK, Q => n18710, QN 
                           => n_3389);
   clk_r_REG5094_S1 : DFF_X1 port map( D => n13810, CK => CLK, Q => n18709, QN 
                           => n_3390);
   clk_r_REG5225_S1 : DFF_X1 port map( D => n13811, CK => CLK, Q => n18708, QN 
                           => n_3391);
   clk_r_REG4887_S1 : DFF_X1 port map( D => n13802, CK => CLK, Q => n18707, QN 
                           => n_3392);
   clk_r_REG5032_S1 : DFF_X1 port map( D => n13815, CK => CLK, Q => n18706, QN 
                           => n_3393);
   clk_r_REG5133_S1 : DFF_X1 port map( D => n14445, CK => CLK, Q => n18705, QN 
                           => n_3394);
   clk_r_REG6096_S1 : DFF_X1 port map( D => n13817, CK => CLK, Q => n18704, QN 
                           => n_3395);
   clk_r_REG6007_S1 : DFF_X1 port map( D => n14431, CK => CLK, Q => n18703, QN 
                           => n_3396);
   clk_r_REG5541_S1 : DFF_X1 port map( D => n13821, CK => CLK, Q => n18702, QN 
                           => n_3397);
   clk_r_REG5476_S1 : DFF_X1 port map( D => n13822, CK => CLK, Q => n18701, QN 
                           => n_3398);
   clk_r_REG5388_S1 : DFF_X1 port map( D => n14430, CK => CLK, Q => n18700, QN 
                           => n_3399);
   clk_r_REG5348_S1 : DFF_X1 port map( D => n13823, CK => CLK, Q => n18699, QN 
                           => n_3400);
   clk_r_REG5778_S1 : DFF_X1 port map( D => n13873, CK => CLK, Q => n18698, QN 
                           => n_3401);
   clk_r_REG5712_S1 : DFF_X1 port map( D => n13872, CK => CLK, Q => n18697, QN 
                           => n_3402);
   clk_r_REG6475_S1 : DFF_X1 port map( D => n13826, CK => CLK, Q => n18696, QN 
                           => n_3403);
   clk_r_REG5316_S1 : DFF_X1 port map( D => n13871, CK => CLK, Q => n18695, QN 
                           => n_3404);
   clk_r_REG6414_S1 : DFF_X1 port map( D => n13828, CK => CLK, Q => n18694, QN 
                           => n_3405);
   clk_r_REG6382_S1 : DFF_X1 port map( D => n13870, CK => CLK, Q => n18693, QN 
                           => n_3406);
   clk_r_REG5844_S1 : DFF_X1 port map( D => n13869, CK => CLK, Q => n18692, QN 
                           => n_3407);
   clk_r_REG5960_S1 : DFF_X1 port map( D => n13804, CK => CLK, Q => n18691, QN 
                           => n_3408);
   clk_r_REG6317_S1 : DFF_X1 port map( D => n13868, CK => CLK, Q => n18690, QN 
                           => n_3409);
   clk_r_REG6217_S1 : DFF_X1 port map( D => n13835, CK => CLK, Q => n18689, QN 
                           => n_3410);
   clk_r_REG6159_S1 : DFF_X1 port map( D => n14290, CK => CLK, Q => n18688, QN 
                           => n_3411);
   clk_r_REG5619_S1 : DFF_X1 port map( D => n14448, CK => CLK, Q => n18687, QN 
                           => n_3412);
   clk_r_REG4963_S1 : DFF_X1 port map( D => n14426, CK => CLK, Q => n18686, QN 
                           => n_3413);
   clk_r_REG4819_S1 : DFF_X1 port map( D => n14433, CK => CLK, Q => n18685, QN 
                           => n_3414);
   clk_r_REG4535_S1 : DFF_X1 port map( D => n14438, CK => CLK, Q => n18684, QN 
                           => n_3415);
   clk_r_REG4737_S1 : DFF_X1 port map( D => n14440, CK => CLK, Q => n18683, QN 
                           => n_3416);
   clk_r_REG6609_S1 : DFF_X1 port map( D => n14451, CK => CLK, Q => n18682, QN 
                           => n_3417);
   clk_r_REG4196_S1 : DFF_X1 port map( D => n14439, CK => CLK, Q => n18681, QN 
                           => n_3418);
   clk_r_REG6543_S1 : DFF_X1 port map( D => n13837, CK => CLK, Q => n18680, QN 
                           => n_3419);
   clk_r_REG4280_S1 : DFF_X1 port map( D => n13833, CK => CLK, Q => n18679, QN 
                           => n_3420);
   clk_r_REG5894_S1 : DFF_X1 port map( D => n13834, CK => CLK, Q => n18678, QN 
                           => n_3421);
   clk_r_REG5096_S1 : DFF_X1 port map( D => n13807, CK => CLK, Q => n18677, QN 
                           => n_3422);
   clk_r_REG5221_S1 : DFF_X1 port map( D => n13841, CK => CLK, Q => n18676, QN 
                           => n_3423);
   clk_r_REG4885_S1 : DFF_X1 port map( D => n13809, CK => CLK, Q => n18675, QN 
                           => n_3424);
   clk_r_REG5028_S1 : DFF_X1 port map( D => n13838, CK => CLK, Q => n18674, QN 
                           => n_3425);
   clk_r_REG5137_S1 : DFF_X1 port map( D => n14429, CK => CLK, Q => n18673, QN 
                           => n_3426);
   clk_r_REG6094_S1 : DFF_X1 port map( D => n13830, CK => CLK, Q => n18672, QN 
                           => n_3427);
   clk_r_REG6009_S1 : DFF_X1 port map( D => n14428, CK => CLK, Q => n18671, QN 
                           => n_3428);
   clk_r_REG5539_S1 : DFF_X1 port map( D => n13831, CK => CLK, Q => n18670, QN 
                           => n_3429);
   clk_r_REG5474_S1 : DFF_X1 port map( D => n13825, CK => CLK, Q => n18669, QN 
                           => n_3430);
   clk_r_REG5390_S1 : DFF_X1 port map( D => n14427, CK => CLK, Q => n18668, QN 
                           => n_3431);
   clk_r_REG5346_S1 : DFF_X1 port map( D => n13839, CK => CLK, Q => n18667, QN 
                           => n_3432);
   clk_r_REG5780_S1 : DFF_X1 port map( D => n13866, CK => CLK, Q => n18666, QN 
                           => n_3433);
   clk_r_REG5716_S1 : DFF_X1 port map( D => n13865, CK => CLK, Q => n18665, QN 
                           => n_3434);
   clk_r_REG6479_S1 : DFF_X1 port map( D => n13798, CK => CLK, Q => n18664, QN 
                           => n_3435);
   clk_r_REG5318_S1 : DFF_X1 port map( D => n13864, CK => CLK, Q => n18663, QN 
                           => n_3436);
   clk_r_REG6412_S1 : DFF_X1 port map( D => n13829, CK => CLK, Q => n18662, QN 
                           => n_3437);
   clk_r_REG6384_S1 : DFF_X1 port map( D => n13863, CK => CLK, Q => n18661, QN 
                           => n_3438);
   clk_r_REG5846_S1 : DFF_X1 port map( D => n13862, CK => CLK, Q => n18660, QN 
                           => n_3439);
   clk_r_REG5958_S1 : DFF_X1 port map( D => n13814, CK => CLK, Q => n18659, QN 
                           => n_3440);
   clk_r_REG6319_S1 : DFF_X1 port map( D => n13861, CK => CLK, Q => n18658, QN 
                           => n_3441);
   clk_r_REG6219_S1 : DFF_X1 port map( D => n13816, CK => CLK, Q => n18657, QN 
                           => n_3442);
   clk_r_REG6155_S1 : DFF_X1 port map( D => n14294, CK => CLK, Q => n18656, QN 
                           => n_3443);
   clk_r_REG5621_S1 : DFF_X1 port map( D => n14442, CK => CLK, Q => n18655, QN 
                           => n_3444);
   clk_r_REG4961_S1 : DFF_X1 port map( D => n14432, CK => CLK, Q => n18654, QN 
                           => n_3445);
   clk_r_REG4817_S1 : DFF_X1 port map( D => n14437, CK => CLK, Q => n18653, QN 
                           => n_3446);
   clk_r_REG4531_S1 : DFF_X1 port map( D => n14449, CK => CLK, Q => n18652, QN 
                           => n_3447);
   clk_r_REG4735_S1 : DFF_X1 port map( D => n14455, CK => CLK, Q => n18651, QN 
                           => n_3448);
   clk_r_REG6611_S1 : DFF_X1 port map( D => n14435, CK => CLK, Q => n18650, QN 
                           => n_3449);
   clk_r_REG4198_S1 : DFF_X1 port map( D => n14436, CK => CLK, Q => n18649, QN 
                           => n_3450);
   clk_r_REG6545_S1 : DFF_X1 port map( D => n13832, CK => CLK, Q => n18648, QN 
                           => n_3451);
   clk_r_REG4284_S1 : DFF_X1 port map( D => n13799, CK => CLK, Q => n18647, QN 
                           => n_3452);
   clk_r_REG5896_S1 : DFF_X1 port map( D => n13824, CK => CLK, Q => n18646, QN 
                           => n_3453);
   clk_r_REG5092_S1 : DFF_X1 port map( D => n13827, CK => CLK, Q => n18645, QN 
                           => n_3454);
   clk_r_REG5223_S1 : DFF_X1 port map( D => n13840, CK => CLK, Q => n18644, QN 
                           => n_3455);
   clk_r_REG4883_S1 : DFF_X1 port map( D => n13819, CK => CLK, Q => n18643, QN 
                           => n_3456);
   clk_r_REG5030_S1 : DFF_X1 port map( D => n13836, CK => CLK, Q => n18642, QN 
                           => n_3457);
   clk_r_REG5135_S1 : DFF_X1 port map( D => n14443, CK => CLK, Q => n18641, QN 
                           => n_3458);
   clk_r_REG6098_S1 : DFF_X1 port map( D => n13813, CK => CLK, Q => n18640, QN 
                           => n_3459);
   clk_r_REG6005_S1 : DFF_X1 port map( D => n14446, CK => CLK, Q => n18639, QN 
                           => n_3460);
   clk_r_REG5543_S1 : DFF_X1 port map( D => n13801, CK => CLK, Q => n18638, QN 
                           => n_3461);
   clk_r_REG5478_S1 : DFF_X1 port map( D => n13820, CK => CLK, Q => n18637, QN 
                           => n_3462);
   clk_r_REG5386_S1 : DFF_X1 port map( D => n14434, CK => CLK, Q => n18636, QN 
                           => n_3463);
   clk_r_REG5350_S1 : DFF_X1 port map( D => n13812, CK => CLK, Q => n18635, QN 
                           => n_3464);
   clk_r_REG5782_S1 : DFF_X1 port map( D => n13860, CK => CLK, Q => n18634, QN 
                           => n_3465);
   clk_r_REG5718_S1 : DFF_X1 port map( D => n13859, CK => CLK, Q => n18633, QN 
                           => n_3466);
   clk_r_REG6477_S1 : DFF_X1 port map( D => n13818, CK => CLK, Q => n18632, QN 
                           => n_3467);
   clk_r_REG5320_S1 : DFF_X1 port map( D => n13857, CK => CLK, Q => n18631, QN 
                           => n_3468);
   clk_r_REG6416_S1 : DFF_X1 port map( D => n13806, CK => CLK, Q => n18630, QN 
                           => n_3469);
   clk_r_REG6386_S1 : DFF_X1 port map( D => n13855, CK => CLK, Q => n18629, QN 
                           => n_3470);
   clk_r_REG5838_S1 : DFF_X1 port map( D => n13884, CK => CLK, Q => n18628, QN 
                           => n_3471);
   clk_r_REG5962_S1 : DFF_X1 port map( D => n13803, CK => CLK, Q => n18627, QN 
                           => n_3472);
   clk_r_REG6321_S1 : DFF_X1 port map( D => n13854, CK => CLK, Q => n18626, QN 
                           => n_3473);
   clk_r_REG6221_S1 : DFF_X1 port map( D => n13797, CK => CLK, Q => n18625, QN 
                           => n_3474);
   clk_r_REG6167_S1 : DFF_X1 port map( D => n13754, CK => CLK, Q => n18624, QN 
                           => n_3475);
   clk_r_REG5641_S1 : DFF_X1 port map( D => n13737, CK => CLK, Q => n18623, QN 
                           => n_3476);
   clk_r_REG4995_S1 : DFF_X1 port map( D => n13710, CK => CLK, Q => n18622, QN 
                           => n_3477);
   clk_r_REG4845_S1 : DFF_X1 port map( D => n13714, CK => CLK, Q => n18621, QN 
                           => n_3478);
   clk_r_REG4555_S1 : DFF_X1 port map( D => n13735, CK => CLK, Q => n18620, QN 
                           => n_3479);
   clk_r_REG4761_S1 : DFF_X1 port map( D => n13693, CK => CLK, Q => n18619, QN 
                           => n_3480);
   clk_r_REG6635_S1 : DFF_X1 port map( D => n13692, CK => CLK, Q => n18618, QN 
                           => n_3481);
   clk_r_REG4214_S1 : DFF_X1 port map( D => n14312, CK => CLK, Q => n18617, QN 
                           => n_3482);
   clk_r_REG6567_S1 : DFF_X1 port map( D => n13585, CK => CLK, Q => n18616, QN 
                           => n_3483);
   clk_r_REG4294_S1 : DFF_X1 port map( D => n13576, CK => CLK, Q => n18615, QN 
                           => n_3484);
   clk_r_REG5864_S1 : DFF_X1 port map( D => n14298, CK => CLK, Q => n18614, QN 
                           => n_3485);
   clk_r_REG5116_S1 : DFF_X1 port map( D => n13639, CK => CLK, Q => n18613, QN 
                           => n_3486);
   clk_r_REG5243_S1 : DFF_X1 port map( D => n13628, CK => CLK, Q => n18612, QN 
                           => n_3487);
   clk_r_REG4903_S1 : DFF_X1 port map( D => n13618, CK => CLK, Q => n18611, QN 
                           => n_3488);
   clk_r_REG5048_S1 : DFF_X1 port map( D => n13604, CK => CLK, Q => n18610, QN 
                           => n_3489);
   clk_r_REG5177_S1 : DFF_X1 port map( D => n13694, CK => CLK, Q => n18609, QN 
                           => n_3490);
   clk_r_REG6106_S1 : DFF_X1 port map( D => n13654, CK => CLK, Q => n18608, QN 
                           => n_3491);
   clk_r_REG5549_S1 : DFF_X1 port map( D => n13671, CK => CLK, Q => n18607, QN 
                           => n_3492);
   clk_r_REG5488_S1 : DFF_X1 port map( D => n13674, CK => CLK, Q => n18606, QN 
                           => n_3493);
   clk_r_REG5406_S1 : DFF_X1 port map( D => n14319, CK => CLK, Q => n18605, QN 
                           => n_3494);
   clk_r_REG5356_S1 : DFF_X1 port map( D => n13664, CK => CLK, Q => n18604, QN 
                           => n_3495);
   clk_r_REG5740_S1 : DFF_X1 port map( D => n14338, CK => CLK, Q => n18603, QN 
                           => n_3496);
   clk_r_REG5676_S1 : DFF_X1 port map( D => n14335, CK => CLK, Q => n18602, QN 
                           => n_3497);
   clk_r_REG6491_S1 : DFF_X1 port map( D => n13583, CK => CLK, Q => n18601, QN 
                           => n_3498);
   clk_r_REG5266_S1 : DFF_X1 port map( D => n14411, CK => CLK, Q => n18600, QN 
                           => n_3499);
   clk_r_REG6434_S1 : DFF_X1 port map( D => n13601, CK => CLK, Q => n18599, QN 
                           => n_3500);
   clk_r_REG6336_S1 : DFF_X1 port map( D => n14397, CK => CLK, Q => n18598, QN 
                           => n_3501);
   clk_r_REG5802_S1 : DFF_X1 port map( D => n14376, CK => CLK, Q => n18597, QN 
                           => n_3502);
   clk_r_REG5982_S1 : DFF_X1 port map( D => n13593, CK => CLK, Q => n18596, QN 
                           => n_3503);
   clk_r_REG6265_S1 : DFF_X1 port map( D => n14377, CK => CLK, Q => n18595, QN 
                           => n_3504);
   clk_r_REG6253_S1 : DFF_X1 port map( D => n13471, CK => CLK, Q => n18594, QN 
                           => n_3505);
   clk_r_REG6179_S1 : DFF_X1 port map( D => n13748, CK => CLK, Q => n18593, QN 
                           => n_3506);
   clk_r_REG5653_S1 : DFF_X1 port map( D => n13720, CK => CLK, Q => n18592, QN 
                           => n_3507);
   clk_r_REG4997_S1 : DFF_X1 port map( D => n13709, CK => CLK, Q => n18591, QN 
                           => n_3508);
   clk_r_REG4843_S1 : DFF_X1 port map( D => n13715, CK => CLK, Q => n18590, QN 
                           => n_3509);
   clk_r_REG4567_S1 : DFF_X1 port map( D => n13707, CK => CLK, Q => n18589, QN 
                           => n_3510);
   clk_r_REG4765_S1 : DFF_X1 port map( D => n13685, CK => CLK, Q => n18588, QN 
                           => n_3511);
   clk_r_REG6637_S1 : DFF_X1 port map( D => n13691, CK => CLK, Q => n18587, QN 
                           => n_3512);
   clk_r_REG4216_S1 : DFF_X1 port map( D => n14311, CK => CLK, Q => n18586, QN 
                           => n_3513);
   clk_r_REG6553_S1 : DFF_X1 port map( D => n13592, CK => CLK, Q => n18585, QN 
                           => n_3514);
   clk_r_REG4292_S1 : DFF_X1 port map( D => n13577, CK => CLK, Q => n18584, QN 
                           => n_3515);
   clk_r_REG5858_S1 : DFF_X1 port map( D => n14301, CK => CLK, Q => n18583, QN 
                           => n_3516);
   clk_r_REG5102_S1 : DFF_X1 port map( D => n13653, CK => CLK, Q => n18582, QN 
                           => n_3517);
   clk_r_REG5245_S1 : DFF_X1 port map( D => n13627, CK => CLK, Q => n18581, QN 
                           => n_3518);
   clk_r_REG4905_S1 : DFF_X1 port map( D => n13617, CK => CLK, Q => n18580, QN 
                           => n_3519);
   clk_r_REG5046_S1 : DFF_X1 port map( D => n13605, CK => CLK, Q => n18579, QN 
                           => n_3520);
   clk_r_REG5175_S1 : DFF_X1 port map( D => n13695, CK => CLK, Q => n18578, QN 
                           => n_3521);
   clk_r_REG6108_S1 : DFF_X1 port map( D => n13652, CK => CLK, Q => n18577, QN 
                           => n_3522);
   clk_r_REG6047_S1 : DFF_X1 port map( D => n13740, CK => CLK, Q => n18576, QN 
                           => n_3523);
   clk_r_REG5551_S1 : DFF_X1 port map( D => n13670, CK => CLK, Q => n18575, QN 
                           => n_3524);
   clk_r_REG5484_S1 : DFF_X1 port map( D => n13676, CK => CLK, Q => n18574, QN 
                           => n_3525);
   clk_r_REG5408_S1 : DFF_X1 port map( D => n14317, CK => CLK, Q => n18573, QN 
                           => n_3526);
   clk_r_REG5358_S1 : DFF_X1 port map( D => n13663, CK => CLK, Q => n18572, QN 
                           => n_3527);
   clk_r_REG5738_S1 : DFF_X1 port map( D => n14340, CK => CLK, Q => n18571, QN 
                           => n_3528);
   clk_r_REG5672_S1 : DFF_X1 port map( D => n14339, CK => CLK, Q => n18570, QN 
                           => n_3529);
   clk_r_REG6501_S1 : DFF_X1 port map( D => n13578, CK => CLK, Q => n18569, QN 
                           => n_3530);
   clk_r_REG3768_S1 : DFF_X1 port map( D => n14421, CK => CLK, Q => n18568, QN 
                           => n_3531);
   clk_r_REG6436_S1 : DFF_X1 port map( D => n13600, CK => CLK, Q => n18567, QN 
                           => n_3532);
   clk_r_REG6332_S1 : DFF_X1 port map( D => n14399, CK => CLK, Q => n18566, QN 
                           => n_3533);
   clk_r_REG5800_S1 : DFF_X1 port map( D => n14378, CK => CLK, Q => n18565, QN 
                           => n_3534);
   clk_r_REG5980_S1 : DFF_X1 port map( D => n13594, CK => CLK, Q => n18564, QN 
                           => n_3535);
   clk_r_REG6267_S1 : DFF_X1 port map( D => n14372, CK => CLK, Q => n18563, QN 
                           => n_3536);
   clk_r_REG6247_S1 : DFF_X1 port map( D => n13478, CK => CLK, Q => n18562, QN 
                           => n_3537);
   clk_r_REG6171_S1 : DFF_X1 port map( D => n13752, CK => CLK, Q => n18561, QN 
                           => n_3538);
   clk_r_REG5651_S1 : DFF_X1 port map( D => n13724, CK => CLK, Q => n18560, QN 
                           => n_3539);
   clk_r_REG4983_S1 : DFF_X1 port map( D => n13734, CK => CLK, Q => n18559, QN 
                           => n_3540);
   clk_r_REG4841_S1 : DFF_X1 port map( D => n13716, CK => CLK, Q => n18558, QN 
                           => n_3541);
   clk_r_REG4565_S1 : DFF_X1 port map( D => n13708, CK => CLK, Q => n18557, QN 
                           => n_3542);
   clk_r_REG4769_S1 : DFF_X1 port map( D => n13683, CK => CLK, Q => n18556, QN 
                           => n_3543);
   clk_r_REG6639_S1 : DFF_X1 port map( D => n13690, CK => CLK, Q => n18555, QN 
                           => n_3544);
   clk_r_REG4210_S1 : DFF_X1 port map( D => n14322, CK => CLK, Q => n18554, QN 
                           => n_3545);
   clk_r_REG6555_S1 : DFF_X1 port map( D => n13591, CK => CLK, Q => n18553, QN 
                           => n_3546);
   clk_r_REG4296_S1 : DFF_X1 port map( D => n13575, CK => CLK, Q => n18552, QN 
                           => n_3547);
   clk_r_REG5868_S1 : DFF_X1 port map( D => n14296, CK => CLK, Q => n18551, QN 
                           => n_3548);
   clk_r_REG5104_S1 : DFF_X1 port map( D => n13646, CK => CLK, Q => n18550, QN 
                           => n_3549);
   clk_r_REG5231_S1 : DFF_X1 port map( D => n13636, CK => CLK, Q => n18549, QN 
                           => n_3550);
   clk_r_REG4907_S1 : DFF_X1 port map( D => n13616, CK => CLK, Q => n18548, QN 
                           => n_3551);
   clk_r_REG5044_S1 : DFF_X1 port map( D => n13607, CK => CLK, Q => n18547, QN 
                           => n_3552);
   clk_r_REG5173_S1 : DFF_X1 port map( D => n13698, CK => CLK, Q => n18546, QN 
                           => n_3553);
   clk_r_REG6110_S1 : DFF_X1 port map( D => n13651, CK => CLK, Q => n18545, QN 
                           => n_3554);
   clk_r_REG6039_S1 : DFF_X1 port map( D => n13746, CK => CLK, Q => n18544, QN 
                           => n_3555);
   clk_r_REG5553_S1 : DFF_X1 port map( D => n13669, CK => CLK, Q => n18543, QN 
                           => n_3556);
   clk_r_REG5486_S1 : DFF_X1 port map( D => n13675, CK => CLK, Q => n18542, QN 
                           => n_3557);
   clk_r_REG5402_S1 : DFF_X1 port map( D => n14324, CK => CLK, Q => n18541, QN 
                           => n_3558);
   clk_r_REG5360_S1 : DFF_X1 port map( D => n13662, CK => CLK, Q => n18540, QN 
                           => n_3559);
   clk_r_REG5736_S1 : DFF_X1 port map( D => n14343, CK => CLK, Q => n18539, QN 
                           => n_3560);
   clk_r_REG5670_S1 : DFF_X1 port map( D => n14341, CK => CLK, Q => n18538, QN 
                           => n_3561);
   clk_r_REG6499_S1 : DFF_X1 port map( D => n13579, CK => CLK, Q => n18537, QN 
                           => n_3562);
   clk_r_REG5268_S1 : DFF_X1 port map( D => n14409, CK => CLK, Q => n18536, QN 
                           => n_3563);
   clk_r_REG6426_S1 : DFF_X1 port map( D => n13614, CK => CLK, Q => n18535, QN 
                           => n_3564);
   clk_r_REG6330_S1 : DFF_X1 port map( D => n14402, CK => CLK, Q => n18534, QN 
                           => n_3565);
   clk_r_REG5798_S1 : DFF_X1 port map( D => n14379, CK => CLK, Q => n18533, QN 
                           => n_3566);
   clk_r_REG5978_S1 : DFF_X1 port map( D => n13595, CK => CLK, Q => n18532, QN 
                           => n_3567);
   clk_r_REG6269_S1 : DFF_X1 port map( D => n14371, CK => CLK, Q => n18531, QN 
                           => n_3568);
   clk_r_REG6257_S1 : DFF_X1 port map( D => n13469, CK => CLK, Q => n18530, QN 
                           => n_3569);
   clk_r_REG6169_S1 : DFF_X1 port map( D => n13753, CK => CLK, Q => n18529, QN 
                           => n_3570);
   clk_r_REG5649_S1 : DFF_X1 port map( D => n13727, CK => CLK, Q => n18528, QN 
                           => n_3571);
   clk_r_REG4985_S1 : DFF_X1 port map( D => n13733, CK => CLK, Q => n18527, QN 
                           => n_3572);
   clk_r_REG4839_S1 : DFF_X1 port map( D => n13717, CK => CLK, Q => n18526, QN 
                           => n_3573);
   clk_r_REG4557_S1 : DFF_X1 port map( D => n13725, CK => CLK, Q => n18525, QN 
                           => n_3574);
   clk_r_REG4767_S1 : DFF_X1 port map( D => n13684, CK => CLK, Q => n18524, QN 
                           => n_3575);
   clk_r_REG6641_S1 : DFF_X1 port map( D => n13688, CK => CLK, Q => n18523, QN 
                           => n_3576);
   clk_r_REG4218_S1 : DFF_X1 port map( D => n14310, CK => CLK, Q => n18522, QN 
                           => n_3577);
   clk_r_REG6565_S1 : DFF_X1 port map( D => n13586, CK => CLK, Q => n18521, QN 
                           => n_3578);
   clk_r_REG4300_S1 : DFF_X1 port map( D => n13573, CK => CLK, Q => n18520, QN 
                           => n_3579);
   clk_r_REG5856_S1 : DFF_X1 port map( D => n14302, CK => CLK, Q => n18519, QN 
                           => n_3580);
   clk_r_REG5106_S1 : DFF_X1 port map( D => n13645, CK => CLK, Q => n18518, QN 
                           => n_3581);
   clk_r_REG5233_S1 : DFF_X1 port map( D => n13635, CK => CLK, Q => n18517, QN 
                           => n_3582);
   clk_r_REG4893_S1 : DFF_X1 port map( D => n13626, CK => CLK, Q => n18516, QN 
                           => n_3583);
   clk_r_REG5042_S1 : DFF_X1 port map( D => n13608, CK => CLK, Q => n18515, QN 
                           => n_3584);
   clk_r_REG5171_S1 : DFF_X1 port map( D => n13699, CK => CLK, Q => n18514, QN 
                           => n_3585);
   clk_r_REG6112_S1 : DFF_X1 port map( D => n13650, CK => CLK, Q => n18513, QN 
                           => n_3586);
   clk_r_REG6049_S1 : DFF_X1 port map( D => n13738, CK => CLK, Q => n18512, QN 
                           => n_3587);
   clk_r_REG5555_S1 : DFF_X1 port map( D => n13668, CK => CLK, Q => n18511, QN 
                           => n_3588);
   clk_r_REG5494_S1 : DFF_X1 port map( D => n13659, CK => CLK, Q => n18510, QN 
                           => n_3589);
   clk_r_REG5410_S1 : DFF_X1 port map( D => n14315, CK => CLK, Q => n18509, QN 
                           => n_3590);
   clk_r_REG5362_S1 : DFF_X1 port map( D => n13661, CK => CLK, Q => n18508, QN 
                           => n_3591);
   clk_r_REG5734_S1 : DFF_X1 port map( D => n14346, CK => CLK, Q => n18507, QN 
                           => n_3592);
   clk_r_REG5668_S1 : DFF_X1 port map( D => n14342, CK => CLK, Q => n18506, QN 
                           => n_3593);
   clk_r_REG6489_S1 : DFF_X1 port map( D => n13584, CK => CLK, Q => n18505, QN 
                           => n_3594);
   clk_r_REG5270_S1 : DFF_X1 port map( D => n14405, CK => CLK, Q => n18504, QN 
                           => n_3595);
   clk_r_REG6428_S1 : DFF_X1 port map( D => n13613, CK => CLK, Q => n18503, QN 
                           => n_3596);
   clk_r_REG6328_S1 : DFF_X1 port map( D => n14403, CK => CLK, Q => n18502, QN 
                           => n_3597);
   clk_r_REG5796_S1 : DFF_X1 port map( D => n14380, CK => CLK, Q => n18501, QN 
                           => n_3598);
   clk_r_REG5976_S1 : DFF_X1 port map( D => n13597, CK => CLK, Q => n18500, QN 
                           => n_3599);
   clk_r_REG6271_S1 : DFF_X1 port map( D => n14370, CK => CLK, Q => n18499, QN 
                           => n_3600);
   clk_r_REG6255_S1 : DFF_X1 port map( D => n13470, CK => CLK, Q => n18498, QN 
                           => n_3601);
   clk_r_REG6173_S1 : DFF_X1 port map( D => n13751, CK => CLK, Q => n18497, QN 
                           => n_3602);
   clk_r_REG5647_S1 : DFF_X1 port map( D => n13728, CK => CLK, Q => n18496, QN 
                           => n_3603);
   clk_r_REG4987_S1 : DFF_X1 port map( D => n13731, CK => CLK, Q => n18495, QN 
                           => n_3604);
   clk_r_REG4851_S1 : DFF_X1 port map( D => n13702, CK => CLK, Q => n18494, QN 
                           => n_3605);
   clk_r_REG4553_S1 : DFF_X1 port map( D => n13739, CK => CLK, Q => n18493, QN 
                           => n_3606);
   clk_r_REG4763_S1 : DFF_X1 port map( D => n13686, CK => CLK, Q => n18492, QN 
                           => n_3607);
   clk_r_REG6643_S1 : DFF_X1 port map( D => n13687, CK => CLK, Q => n18491, QN 
                           => n_3608);
   clk_r_REG4206_S1 : DFF_X1 port map( D => n14326, CK => CLK, Q => n18490, QN 
                           => n_3609);
   clk_r_REG6557_S1 : DFF_X1 port map( D => n13590, CK => CLK, Q => n18489, QN 
                           => n_3610);
   clk_r_REG4304_S1 : DFF_X1 port map( D => n13571, CK => CLK, Q => n18488, QN 
                           => n_3611);
   clk_r_REG5862_S1 : DFF_X1 port map( D => n14299, CK => CLK, Q => n18487, QN 
                           => n_3612);
   clk_r_REG5108_S1 : DFF_X1 port map( D => n13643, CK => CLK, Q => n18486, QN 
                           => n_3613);
   clk_r_REG5235_S1 : DFF_X1 port map( D => n13634, CK => CLK, Q => n18485, QN 
                           => n_3614);
   clk_r_REG4895_S1 : DFF_X1 port map( D => n13625, CK => CLK, Q => n18484, QN 
                           => n_3615);
   clk_r_REG5040_S1 : DFF_X1 port map( D => n13609, CK => CLK, Q => n18483, QN 
                           => n_3616);
   clk_r_REG5179_S1 : DFF_X1 port map( D => n13689, CK => CLK, Q => n18482, QN 
                           => n_3617);
   clk_r_REG6114_S1 : DFF_X1 port map( D => n13649, CK => CLK, Q => n18481, QN 
                           => n_3618);
   clk_r_REG6051_S1 : DFF_X1 port map( D => n13736, CK => CLK, Q => n18480, QN 
                           => n_3619);
   clk_r_REG5557_S1 : DFF_X1 port map( D => n13667, CK => CLK, Q => n18479, QN 
                           => n_3620);
   clk_r_REG5490_S1 : DFF_X1 port map( D => n13673, CK => CLK, Q => n18478, QN 
                           => n_3621);
   clk_r_REG5400_S1 : DFF_X1 port map( D => n14328, CK => CLK, Q => n18477, QN 
                           => n_3622);
   clk_r_REG5364_S1 : DFF_X1 port map( D => n13660, CK => CLK, Q => n18476, QN 
                           => n_3623);
   clk_r_REG5732_S1 : DFF_X1 port map( D => n14348, CK => CLK, Q => n18475, QN 
                           => n_3624);
   clk_r_REG3701_S1 : DFF_X1 port map( D => n14382, CK => CLK, Q => n18474, QN 
                           => n_3625);
   clk_r_REG6495_S1 : DFF_X1 port map( D => n13581, CK => CLK, Q => n18473, QN 
                           => n_3626);
   clk_r_REG5274_S1 : DFF_X1 port map( D => n14357, CK => CLK, Q => n18472, QN 
                           => n_3627);
   clk_r_REG6430_S1 : DFF_X1 port map( D => n13612, CK => CLK, Q => n18471, QN 
                           => n_3628);
   clk_r_REG3562_S1 : DFF_X1 port map( D => n14424, CK => CLK, Q => n18470, QN 
                           => n_3629);
   clk_r_REG5794_S1 : DFF_X1 port map( D => n14387, CK => CLK, Q => n18469, QN 
                           => n_3630);
   clk_r_REG5974_S1 : DFF_X1 port map( D => n13598, CK => CLK, Q => n18468, QN 
                           => n_3631);
   clk_r_REG6273_S1 : DFF_X1 port map( D => n14369, CK => CLK, Q => n18467, QN 
                           => n_3632);
   clk_r_REG6245_S1 : DFF_X1 port map( D => n13479, CK => CLK, Q => n18466, QN 
                           => n_3633);
   clk_r_REG6181_S1 : DFF_X1 port map( D => n13747, CK => CLK, Q => n18465, QN 
                           => n_3634);
   clk_r_REG5645_S1 : DFF_X1 port map( D => n13729, CK => CLK, Q => n18464, QN 
                           => n_3635);
   clk_r_REG4991_S1 : DFF_X1 port map( D => n13721, CK => CLK, Q => n18463, QN 
                           => n_3636);
   clk_r_REG4849_S1 : DFF_X1 port map( D => n13703, CK => CLK, Q => n18462, QN 
                           => n_3637);
   clk_r_REG4561_S1 : DFF_X1 port map( D => n13718, CK => CLK, Q => n18461, QN 
                           => n_3638);
   clk_r_REG4759_S1 : DFF_X1 port map( D => n13696, CK => CLK, Q => n18460, QN 
                           => n_3639);
   clk_r_REG6633_S1 : DFF_X1 port map( D => n13697, CK => CLK, Q => n18459, QN 
                           => n_3640);
   clk_r_REG4208_S1 : DFF_X1 port map( D => n14325, CK => CLK, Q => n18458, QN 
                           => n_3641);
   clk_r_REG6563_S1 : DFF_X1 port map( D => n13587, CK => CLK, Q => n18457, QN 
                           => n_3642);
   clk_r_REG4302_S1 : DFF_X1 port map( D => n13572, CK => CLK, Q => n18456, QN 
                           => n_3643);
   clk_r_REG5854_S1 : DFF_X1 port map( D => n14303, CK => CLK, Q => n18455, QN 
                           => n_3644);
   clk_r_REG5110_S1 : DFF_X1 port map( D => n13642, CK => CLK, Q => n18454, QN 
                           => n_3645);
   clk_r_REG5237_S1 : DFF_X1 port map( D => n13633, CK => CLK, Q => n18453, QN 
                           => n_3646);
   clk_r_REG4897_S1 : DFF_X1 port map( D => n13624, CK => CLK, Q => n18452, QN 
                           => n_3647);
   clk_r_REG5052_S1 : DFF_X1 port map( D => n13602, CK => CLK, Q => n18451, QN 
                           => n_3648);
   clk_r_REG5169_S1 : DFF_X1 port map( D => n13700, CK => CLK, Q => n18450, QN 
                           => n_3649);
   clk_r_REG6116_S1 : DFF_X1 port map( D => n13648, CK => CLK, Q => n18449, QN 
                           => n_3650);
   clk_r_REG6041_S1 : DFF_X1 port map( D => n13745, CK => CLK, Q => n18448, QN 
                           => n_3651);
   clk_r_REG5559_S1 : DFF_X1 port map( D => n13666, CK => CLK, Q => n18447, QN 
                           => n_3652);
   clk_r_REG5492_S1 : DFF_X1 port map( D => n13672, CK => CLK, Q => n18446, QN 
                           => n_3653);
   clk_r_REG5396_S1 : DFF_X1 port map( D => n14333, CK => CLK, Q => n18445, QN 
                           => n_3654);
   clk_r_REG5366_S1 : DFF_X1 port map( D => n13658, CK => CLK, Q => n18444, QN 
                           => n_3655);
   clk_r_REG5730_S1 : DFF_X1 port map( D => n14349, CK => CLK, Q => n18443, QN 
                           => n_3656);
   clk_r_REG5660_S1 : DFF_X1 port map( D => n14367, CK => CLK, Q => n18442, QN 
                           => n_3657);
   clk_r_REG6493_S1 : DFF_X1 port map( D => n13582, CK => CLK, Q => n18441, QN 
                           => n_3658);
   clk_r_REG5276_S1 : DFF_X1 port map( D => n14345, CK => CLK, Q => n18440, QN 
                           => n_3659);
   clk_r_REG6432_S1 : DFF_X1 port map( D => n13611, CK => CLK, Q => n18439, QN 
                           => n_3660);
   clk_r_REG6326_S1 : DFF_X1 port map( D => n14407, CK => CLK, Q => n18438, QN 
                           => n_3661);
   clk_r_REG5792_S1 : DFF_X1 port map( D => n14388, CK => CLK, Q => n18437, QN 
                           => n_3662);
   clk_r_REG5972_S1 : DFF_X1 port map( D => n13599, CK => CLK, Q => n18436, QN 
                           => n_3663);
   clk_r_REG3572_S1 : DFF_X1 port map( D => n14401, CK => CLK, Q => n18435, QN 
                           => n_3664);
   clk_r_REG6251_S1 : DFF_X1 port map( D => n13476, CK => CLK, Q => n18434, QN 
                           => n_3665);
   clk_r_REG6175_S1 : DFF_X1 port map( D => n13750, CK => CLK, Q => n18433, QN 
                           => n_3666);
   clk_r_REG5643_S1 : DFF_X1 port map( D => n13730, CK => CLK, Q => n18432, QN 
                           => n_3667);
   clk_r_REG4993_S1 : DFF_X1 port map( D => n13713, CK => CLK, Q => n18431, QN 
                           => n_3668);
   clk_r_REG4847_S1 : DFF_X1 port map( D => n13706, CK => CLK, Q => n18430, QN 
                           => n_3669);
   clk_r_REG4559_S1 : DFF_X1 port map( D => n13719, CK => CLK, Q => n18429, QN 
                           => n_3670);
   clk_r_REG4755_S1 : DFF_X1 port map( D => n13704, CK => CLK, Q => n18428, QN 
                           => n_3671);
   clk_r_REG6631_S1 : DFF_X1 port map( D => n13705, CK => CLK, Q => n18427, QN 
                           => n_3672);
   clk_r_REG4212_S1 : DFF_X1 port map( D => n14313, CK => CLK, Q => n18426, QN 
                           => n_3673);
   clk_r_REG6559_S1 : DFF_X1 port map( D => n13589, CK => CLK, Q => n18425, QN 
                           => n_3674);
   clk_r_REG4298_S1 : DFF_X1 port map( D => n13574, CK => CLK, Q => n18424, QN 
                           => n_3675);
   clk_r_REG3658_S1 : DFF_X1 port map( D => n14307, CK => CLK, Q => n18423, QN 
                           => n_3676);
   clk_r_REG5112_S1 : DFF_X1 port map( D => n13641, CK => CLK, Q => n18422, QN 
                           => n_3677);
   clk_r_REG5239_S1 : DFF_X1 port map( D => n13632, CK => CLK, Q => n18421, QN 
                           => n_3678);
   clk_r_REG4899_S1 : DFF_X1 port map( D => n13623, CK => CLK, Q => n18420, QN 
                           => n_3679);
   clk_r_REG5050_S1 : DFF_X1 port map( D => n13603, CK => CLK, Q => n18419, QN 
                           => n_3680);
   clk_r_REG5167_S1 : DFF_X1 port map( D => n13711, CK => CLK, Q => n18418, QN 
                           => n_3681);
   clk_r_REG6118_S1 : DFF_X1 port map( D => n13647, CK => CLK, Q => n18417, QN 
                           => n_3682);
   clk_r_REG6043_S1 : DFF_X1 port map( D => n13744, CK => CLK, Q => n18416, QN 
                           => n_3683);
   clk_r_REG5561_S1 : DFF_X1 port map( D => n13665, CK => CLK, Q => n18415, QN 
                           => n_3684);
   clk_r_REG5496_S1 : DFF_X1 port map( D => n13656, CK => CLK, Q => n18414, QN 
                           => n_3685);
   clk_r_REG5404_S1 : DFF_X1 port map( D => n14321, CK => CLK, Q => n18413, QN 
                           => n_3686);
   clk_r_REG5368_S1 : DFF_X1 port map( D => n13657, CK => CLK, Q => n18412, QN 
                           => n_3687);
   clk_r_REG5728_S1 : DFF_X1 port map( D => n14350, CK => CLK, Q => n18411, QN 
                           => n_3688);
   clk_r_REG5662_S1 : DFF_X1 port map( D => n14366, CK => CLK, Q => n18410, QN 
                           => n_3689);
   clk_r_REG6515_S1 : DFF_X1 port map( D => n13472, CK => CLK, Q => n18409, QN 
                           => n_3690);
   clk_r_REG5306_S1 : DFF_X1 port map( D => n13905, CK => CLK, Q => n18408, QN 
                           => n_3691);
   clk_r_REG6448_S1 : DFF_X1 port map( D => n13481, CK => CLK, Q => n18407, QN 
                           => n_3692);
   clk_r_REG6376_S1 : DFF_X1 port map( D => n13885, CK => CLK, Q => n18406, QN 
                           => n_3693);
   clk_r_REG5830_S1 : DFF_X1 port map( D => n13903, CK => CLK, Q => n18405, QN 
                           => n_3694);
   clk_r_REG5996_S1 : DFF_X1 port map( D => n13474, CK => CLK, Q => n18404, QN 
                           => n_3695);
   clk_r_REG6309_S1 : DFF_X1 port map( D => n13902, CK => CLK, Q => n18403, QN 
                           => n_3696);
   clk_r_REG6249_S1 : DFF_X1 port map( D => n13477, CK => CLK, Q => n18402, QN 
                           => n_3697);
   clk_r_REG6177_S1 : DFF_X1 port map( D => n13749, CK => CLK, Q => n18401, QN 
                           => n_3698);
   clk_r_REG5639_S1 : DFF_X1 port map( D => n13743, CK => CLK, Q => n18400, QN 
                           => n_3699);
   clk_r_REG4989_S1 : DFF_X1 port map( D => n13722, CK => CLK, Q => n18399, QN 
                           => n_3700);
   clk_r_REG4837_S1 : DFF_X1 port map( D => n13723, CK => CLK, Q => n18398, QN 
                           => n_3701);
   clk_r_REG4563_S1 : DFF_X1 port map( D => n13712, CK => CLK, Q => n18397, QN 
                           => n_3702);
   clk_r_REG4757_S1 : DFF_X1 port map( D => n13701, CK => CLK, Q => n18396, QN 
                           => n_3703);
   clk_r_REG6629_S1 : DFF_X1 port map( D => n13726, CK => CLK, Q => n18395, QN 
                           => n_3704);
   clk_r_REG4204_S1 : DFF_X1 port map( D => n14331, CK => CLK, Q => n18394, QN 
                           => n_3705);
   clk_r_REG6561_S1 : DFF_X1 port map( D => n13588, CK => CLK, Q => n18393, QN 
                           => n_3706);
   clk_r_REG4306_S1 : DFF_X1 port map( D => n13570, CK => CLK, Q => n18392, QN 
                           => n_3707);
   clk_r_REG5850_S1 : DFF_X1 port map( D => n14305, CK => CLK, Q => n18391, QN 
                           => n_3708);
   clk_r_REG5114_S1 : DFF_X1 port map( D => n13640, CK => CLK, Q => n18390, QN 
                           => n_3709);
   clk_r_REG5241_S1 : DFF_X1 port map( D => n13631, CK => CLK, Q => n18389, QN 
                           => n_3710);
   clk_r_REG4901_S1 : DFF_X1 port map( D => n13622, CK => CLK, Q => n18388, QN 
                           => n_3711);
   clk_r_REG5038_S1 : DFF_X1 port map( D => n13732, CK => CLK, Q => n18387, QN 
                           => n_3712);
   clk_r_REG5181_S1 : DFF_X1 port map( D => n13606, CK => CLK, Q => n18386, QN 
                           => n_3713);
   clk_r_REG6104_S1 : DFF_X1 port map( D => n13741, CK => CLK, Q => n18385, QN 
                           => n_3714);
   clk_r_REG6053_S1 : DFF_X1 port map( D => n13637, CK => CLK, Q => n18384, QN 
                           => n_3715);
   clk_r_REG5563_S1 : DFF_X1 port map( D => n13629, CK => CLK, Q => n18383, QN 
                           => n_3716);
   clk_r_REG5498_S1 : DFF_X1 port map( D => n13644, CK => CLK, Q => n18382, QN 
                           => n_3717);
   clk_r_REG5398_S1 : DFF_X1 port map( D => n14329, CK => CLK, Q => n18381, QN 
                           => n_3718);
   clk_r_REG5370_S1 : DFF_X1 port map( D => n13655, CK => CLK, Q => n18380, QN 
                           => n_3719);
   clk_r_REG5726_S1 : DFF_X1 port map( D => n14351, CK => CLK, Q => n18379, QN 
                           => n_3720);
   clk_r_REG5664_S1 : DFF_X1 port map( D => n14359, CK => CLK, Q => n18378, QN 
                           => n_3721);
   clk_r_REG5312_S1 : DFF_X1 port map( D => n13883, CK => CLK, Q => n18377, QN 
                           => n_3722);
   clk_r_REG6450_S1 : DFF_X1 port map( D => n13473, CK => CLK, Q => n18376, QN 
                           => n_3723);
   clk_r_REG6378_S1 : DFF_X1 port map( D => n13882, CK => CLK, Q => n18375, QN 
                           => n_3724);
   clk_r_REG5840_S1 : DFF_X1 port map( D => n13881, CK => CLK, Q => n18374, QN 
                           => n_3725);
   clk_r_REG5994_S1 : DFF_X1 port map( D => n13475, CK => CLK, Q => n18373, QN 
                           => n_3726);
   clk_r_REG6313_S1 : DFF_X1 port map( D => n13880, CK => CLK, Q => n18372, QN 
                           => n_3727);
   clk_r_REG6243_S1 : DFF_X1 port map( D => n13482, CK => CLK, Q => n18371, QN 
                           => n_3728);
   clk_r_REG6879_S6 : DFFR_X1 port map( D => ADD_RD2(3), CK => CLK, RN => 
                           RESET_BAR, Q => n18370, QN => n_3729);
   clk_r_REG6849_S6 : DFFR_X1 port map( D => ADD_RD1(3), CK => CLK, RN => 
                           RESET_BAR, Q => n18369, QN => n_3730);
   clk_r_REG6808_S6 : DFFS_X1 port map( D => n25146, CK => CLK, SN => RESET_BAR
                           , Q => n25155, QN => n26756);
   clk_r_REG6805_S6 : DFFS_X1 port map( D => n25147, CK => CLK, SN => RESET_BAR
                           , Q => n_3731, QN => n26755);
   clk_r_REG6789_S6 : DFFS_X1 port map( D => n25143, CK => CLK, SN => RESET_BAR
                           , Q => n25150, QN => n26758);
   clk_r_REG6802_S6 : DFFS_X1 port map( D => n25148, CK => CLK, SN => RESET_BAR
                           , Q => n25154, QN => n26757);
   clk_r_REG6722_S5 : DFFR_X1 port map( D => n14634, CK => CLK, RN => RESET_BAR
                           , Q => n18358, QN => n_3732);
   clk_r_REG6721_S5 : DFFR_X1 port map( D => n14635, CK => CLK, RN => RESET_BAR
                           , Q => n18356, QN => n_3733);
   clk_r_REG6718_S5 : DFFR_X1 port map( D => n14638, CK => CLK, RN => RESET_BAR
                           , Q => n18352, QN => n_3734);
   clk_r_REG6717_S5 : DFFR_X1 port map( D => n14640, CK => CLK, RN => RESET_BAR
                           , Q => n18350, QN => n_3735);
   clk_r_REG6893_S6 : DFFS_X1 port map( D => n25158, CK => CLK, SN => RESET_BAR
                           , Q => n25153, QN => n26760);
   clk_r_REG6888_S6 : DFFS_X1 port map( D => n25157, CK => CLK, SN => RESET_BAR
                           , Q => n25152, QN => n26761);
   clk_r_REG6799_S6 : DFFS_X1 port map( D => n25145, CK => CLK, SN => RESET_BAR
                           , Q => n_3736, QN => n26754);
   clk_r_REG6796_S6 : DFFS_X1 port map( D => n25144, CK => CLK, SN => RESET_BAR
                           , Q => n25151, QN => n26759);
   clk_r_REG6724_S5 : DFFS_X1 port map( D => n14632, CK => CLK, SN => RESET_BAR
                           , Q => n18284, QN => n_3737);
   clk_r_REG6723_S5 : DFFR_X1 port map( D => n14633, CK => CLK, RN => RESET_BAR
                           , Q => n18283, QN => n_3738);
   clk_r_REG6720_S5 : DFFR_X1 port map( D => n14636, CK => CLK, RN => RESET_BAR
                           , Q => n18282, QN => n_3739);
   clk_r_REG6719_S5 : DFFR_X1 port map( D => n14637, CK => CLK, RN => RESET_BAR
                           , Q => n18281, QN => n_3740);
   clk_r_REG6810_S6 : DFFR_X1 port map( D => n11172, CK => CLK, RN => RESET_BAR
                           , Q => n18319, QN => n_3741);
   clk_r_REG6801_S6 : DFFR_X1 port map( D => n11174, CK => CLK, RN => RESET_BAR
                           , Q => n18323, QN => n_3742);
   clk_r_REG6804_S6 : DFFR_X1 port map( D => n11189, CK => CLK, RN => RESET_BAR
                           , Q => n18313, QN => n_3743);
   clk_r_REG6795_S6 : DFFR_X1 port map( D => n11173, CK => CLK, RN => RESET_BAR
                           , Q => n18322, QN => n_3744);
   clk_r_REG6800_S6 : DFFR_X1 port map( D => n11186, CK => CLK, RN => RESET_BAR
                           , Q => n18310, QN => n_3745);
   clk_r_REG6844_S6 : DFFR_X1 port map( D => n11137, CK => CLK, RN => RESET_BAR
                           , Q => n18300, QN => n_3746);
   clk_r_REG6835_S6 : DFFR_X1 port map( D => n11152, CK => CLK, RN => RESET_BAR
                           , Q => n18303, QN => n_3747);
   clk_r_REG6841_S6 : DFFR_X1 port map( D => n11140, CK => CLK, RN => RESET_BAR
                           , Q => n18295, QN => n_3748);
   clk_r_REG6840_S6 : DFFR_X1 port map( D => n11142, CK => CLK, RN => RESET_BAR
                           , Q => n18294, QN => n_3749);
   clk_r_REG6833_S6 : DFFR_X1 port map( D => n11151, CK => CLK, RN => RESET_BAR
                           , Q => n18301, QN => n_3750);
   clk_r_REG6845_S6 : DFFR_X1 port map( D => n11153, CK => CLK, RN => RESET_BAR
                           , Q => n18305, QN => n_3751);
   clk_r_REG6797_S6 : DFFR_X1 port map( D => n11190, CK => CLK, RN => RESET_BAR
                           , Q => n18315, QN => n_3752);
   clk_r_REG6898_S6 : DFFS_X1 port map( D => n1517, CK => CLK, SN => RESET_BAR,
                           Q => n_3753, QN => n18367);
   clk_r_REG6794_S6 : DFFR_X1 port map( D => n11168, CK => CLK, RN => RESET_BAR
                           , Q => n18320, QN => n_3754);
   clk_r_REG6807_S6 : DFFR_X1 port map( D => n11191, CK => CLK, RN => RESET_BAR
                           , Q => n18321, QN => n_3755);
   clk_r_REG6806_S6 : DFFR_X1 port map( D => n11165, CK => CLK, RN => RESET_BAR
                           , Q => n18317, QN => n_3756);
   clk_r_REG6813_S6 : DFFR_X1 port map( D => n11157, CK => CLK, RN => RESET_BAR
                           , Q => n18314, QN => n_3757);
   clk_r_REG6837_S6 : DFFR_X1 port map( D => n11136, CK => CLK, RN => RESET_BAR
                           , Q => n18306, QN => n_3758);
   clk_r_REG6834_S6 : DFFR_X1 port map( D => n11141, CK => CLK, RN => RESET_BAR
                           , Q => n18302, QN => n_3759);
   clk_r_REG6842_S6 : DFFR_X1 port map( D => n11149, CK => CLK, RN => RESET_BAR
                           , Q => n18297, QN => n_3760);
   clk_r_REG6838_S6 : DFFR_X1 port map( D => n11154, CK => CLK, RN => RESET_BAR
                           , Q => n18307, QN => n_3761);
   clk_r_REG6846_S6 : DFFR_X1 port map( D => n11132, CK => CLK, RN => RESET_BAR
                           , Q => n18308, QN => n_3762);
   clk_r_REG6843_S6 : DFFR_X1 port map( D => n11150, CK => CLK, RN => RESET_BAR
                           , Q => n18299, QN => n_3763);
   clk_r_REG6814_S6 : DFFR_X1 port map( D => n11167, CK => CLK, RN => RESET_BAR
                           , Q => n18316, QN => n_3764);
   clk_r_REG6811_S6 : DFFR_X1 port map( D => n1520, CK => CLK, RN => RESET_BAR,
                           Q => n_3765, QN => n18291);
   clk_r_REG6896_S6 : DFFR_X1 port map( D => n1518, CK => CLK, RN => RESET_BAR,
                           Q => n_3766, QN => n18292);
   clk_r_REG6889_S6 : DFFS_X1 port map( D => n1515, CK => CLK, SN => RESET_BAR,
                           Q => n_3767, QN => n18363);
   clk_r_REG6809_S6 : DFFR_X1 port map( D => n11187, CK => CLK, RN => RESET_BAR
                           , Q => n18311, QN => n_3768);
   clk_r_REG6798_S6 : DFFR_X1 port map( D => n11175, CK => CLK, RN => RESET_BAR
                           , Q => n18324, QN => n_3769);
   clk_r_REG6836_S6 : DFFR_X1 port map( D => n11139, CK => CLK, RN => RESET_BAR
                           , Q => n18304, QN => n_3770);
   clk_r_REG6832_S6 : DFFR_X1 port map( D => n11138, CK => CLK, RN => RESET_BAR
                           , Q => n18298, QN => n_3771);
   clk_r_REG6831_S6 : DFFR_X1 port map( D => n11133, CK => CLK, RN => RESET_BAR
                           , Q => n18296, QN => n_3772);
   clk_r_REG6839_S6 : DFFR_X1 port map( D => n11143, CK => CLK, RN => RESET_BAR
                           , Q => n18293, QN => n_3773);
   clk_r_REG6791_S6 : DFFR_X1 port map( D => n11166, CK => CLK, RN => RESET_BAR
                           , Q => n18318, QN => n_3774);
   clk_r_REG6790_S6 : DFFR_X1 port map( D => n11162, CK => CLK, RN => RESET_BAR
                           , Q => n18309, QN => n_3775);
   clk_r_REG6792_S6 : DFFS_X1 port map( D => n1521, CK => CLK, SN => RESET_BAR,
                           Q => n_3776, QN => n18288);
   clk_r_REG6900_S6 : DFFS_X1 port map( D => n1516, CK => CLK, SN => RESET_BAR,
                           Q => n_3777, QN => n18368);
   clk_r_REG6894_S6 : DFFS_X1 port map( D => n1519, CK => CLK, SN => RESET_BAR,
                           Q => n_3778, QN => n18290);
   clk_r_REG6891_S6 : DFFS_X1 port map( D => n1514, CK => CLK, SN => RESET_BAR,
                           Q => n_3779, QN => n18364);
   clk_r_REG6803_S6 : DFFR_X1 port map( D => n11188, CK => CLK, RN => RESET_BAR
                           , Q => n18312, QN => n_3780);
   clk_r_REG6897_S6 : DFFS_X1 port map( D => n11231, CK => CLK, SN => RESET_BAR
                           , Q => n19400, QN => n_3781);
   clk_r_REG6901_S6 : DFFR_X1 port map( D => n11225, CK => CLK, RN => RESET_BAR
                           , Q => n19398, QN => n_3782);
   clk_r_REG6895_S6 : DFFR_X1 port map( D => n11230, CK => CLK, RN => RESET_BAR
                           , Q => n19399, QN => n_3783);
   clk_r_REG6892_S6 : DFFR_X1 port map( D => n11232, CK => CLK, RN => RESET_BAR
                           , Q => n19397, QN => n_3784);
   clk_r_REG6890_S6 : DFFR_X1 port map( D => n11228, CK => CLK, RN => RESET_BAR
                           , Q => n19396, QN => n_3785);
   clk_r_REG6696_S6 : DFFS_X2 port map( D => n10100, CK => CLK, SN => RESET_BAR
                           , Q => n18357, QN => n_3786);
   clk_r_REG6697_S6 : DFFS_X2 port map( D => n10101, CK => CLK, SN => RESET_BAR
                           , Q => n18359, QN => n_3787);
   clk_r_REG6698_S6 : DFFS_X2 port map( D => n10102, CK => CLK, SN => RESET_BAR
                           , Q => n18360, QN => n_3788);
   clk_r_REG6694_S6 : DFFS_X2 port map( D => n10098, CK => CLK, SN => RESET_BAR
                           , Q => n18354, QN => n_3789);
   clk_r_REG6695_S6 : DFFS_X2 port map( D => n10099, CK => CLK, SN => RESET_BAR
                           , Q => n18355, QN => n_3790);
   clk_r_REG6692_S6 : DFFS_X2 port map( D => n10096, CK => CLK, SN => RESET_BAR
                           , Q => n18351, QN => n_3791);
   clk_r_REG6693_S6 : DFFS_X2 port map( D => n10097, CK => CLK, SN => RESET_BAR
                           , Q => n18353, QN => n_3792);
   clk_r_REG6682_S6 : DFFS_X2 port map( D => n10094, CK => CLK, SN => RESET_BAR
                           , Q => n18348, QN => n_3793);
   clk_r_REG6691_S6 : DFFS_X2 port map( D => n10095, CK => CLK, SN => RESET_BAR
                           , Q => n18349, QN => n_3794);
   clk_r_REG6680_S6 : DFFS_X2 port map( D => n10092, CK => CLK, SN => RESET_BAR
                           , Q => n18346, QN => n_3795);
   clk_r_REG6681_S6 : DFFS_X2 port map( D => n10093, CK => CLK, SN => RESET_BAR
                           , Q => n18347, QN => n_3796);
   clk_r_REG6678_S6 : DFFS_X2 port map( D => n10090, CK => CLK, SN => RESET_BAR
                           , Q => n18344, QN => n_3797);
   clk_r_REG6679_S6 : DFFS_X2 port map( D => n10091, CK => CLK, SN => RESET_BAR
                           , Q => n18345, QN => n_3798);
   clk_r_REG6676_S6 : DFFS_X2 port map( D => n10088, CK => CLK, SN => RESET_BAR
                           , Q => n18342, QN => n_3799);
   clk_r_REG6677_S6 : DFFS_X2 port map( D => n10089, CK => CLK, SN => RESET_BAR
                           , Q => n18343, QN => n_3800);
   clk_r_REG6690_S6 : DFFS_X2 port map( D => n10086, CK => CLK, SN => RESET_BAR
                           , Q => n18340, QN => n_3801);
   clk_r_REG6688_S6 : DFFS_X2 port map( D => n10084, CK => CLK, SN => RESET_BAR
                           , Q => n18338, QN => n_3802);
   clk_r_REG6689_S6 : DFFS_X2 port map( D => n10085, CK => CLK, SN => RESET_BAR
                           , Q => n18339, QN => n_3803);
   clk_r_REG6686_S6 : DFFS_X2 port map( D => n10082, CK => CLK, SN => RESET_BAR
                           , Q => n18336, QN => n_3804);
   clk_r_REG6684_S6 : DFFS_X2 port map( D => n10080, CK => CLK, SN => RESET_BAR
                           , Q => n18334, QN => n_3805);
   clk_r_REG6685_S6 : DFFS_X2 port map( D => n10081, CK => CLK, SN => RESET_BAR
                           , Q => n18335, QN => n_3806);
   clk_r_REG6674_S6 : DFFS_X2 port map( D => n10078, CK => CLK, SN => RESET_BAR
                           , Q => n18332, QN => n_3807);
   clk_r_REG6683_S6 : DFFS_X2 port map( D => n10079, CK => CLK, SN => RESET_BAR
                           , Q => n18333, QN => n_3808);
   clk_r_REG6672_S6 : DFFS_X2 port map( D => n10076, CK => CLK, SN => RESET_BAR
                           , Q => n18330, QN => n_3809);
   clk_r_REG6673_S6 : DFFS_X2 port map( D => n10077, CK => CLK, SN => RESET_BAR
                           , Q => n18331, QN => n_3810);
   clk_r_REG6670_S6 : DFFS_X2 port map( D => n10074, CK => CLK, SN => RESET_BAR
                           , Q => n18328, QN => n_3811);
   clk_r_REG6671_S6 : DFFS_X2 port map( D => n10075, CK => CLK, SN => RESET_BAR
                           , Q => n18329, QN => n_3812);
   clk_r_REG6668_S6 : DFFS_X2 port map( D => n10072, CK => CLK, SN => RESET_BAR
                           , Q => n18326, QN => n_3813);
   clk_r_REG6669_S6 : DFFS_X2 port map( D => n10073, CK => CLK, SN => RESET_BAR
                           , Q => n18327, QN => n_3814);
   clk_r_REG6667_S6 : DFFS_X2 port map( D => n10071, CK => CLK, SN => RESET_BAR
                           , Q => n18325, QN => n_3815);
   clk_r_REG6675_S6 : DFFS_X2 port map( D => n10087, CK => CLK, SN => RESET_BAR
                           , Q => n18341, QN => n_3816);
   clk_r_REG6687_S6 : DFFS_X2 port map( D => n10083, CK => CLK, SN => RESET_BAR
                           , Q => n18337, QN => n_3817);
   U3 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18342, ZN => n25241);
   U4 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18343, ZN => n25236);
   U5 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18339, ZN => n25225);
   U6 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18344, ZN => n25238);
   U7 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18340, ZN => n25240);
   U8 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18334, ZN => n25244);
   U9 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18333, ZN => n25213);
   U10 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18338, ZN => n25214);
   U11 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18332, ZN => n25243);
   U12 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18331, ZN => n25242);
   U13 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18335, ZN => n25239);
   U14 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18336, ZN => n25231);
   U15 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18345, ZN => n25245);
   U16 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18346, ZN => n25233);
   U17 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18347, ZN => n25232);
   U18 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18348, ZN => n25234);
   U19 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18328, ZN => n25187);
   U20 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18326, ZN => n25189);
   U21 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18327, ZN => n25191);
   U22 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18330, ZN => n25188);
   U23 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18329, ZN => n25192);
   U24 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18325, ZN => n25190);
   U25 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18355, ZN => n25221);
   U26 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18351, ZN => n25218);
   U27 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18357, ZN => n25220);
   U28 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18360, ZN => n25193);
   U29 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18359, ZN => n25194);
   U30 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18349, ZN => n25219);
   U31 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18354, ZN => n25217);
   U32 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n18353, ZN => n25215);
   U33 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n18341, ZN => n25227);
   U34 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n18337, ZN => n25235);
   U35 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n20442, ZN => n25201);
   U36 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n20460, ZN => n25205);
   U37 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n20470, A3 => n20467, ZN => 
                           n26012);
   U38 : CLKBUF_X1 port map( A => n26012, Z => n25828);
   U39 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n20470, A3 => n20468, ZN => 
                           n26753);
   U40 : CLKBUF_X1 port map( A => n26753, Z => n26689);
   U41 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n25268);
   U42 : INV_X1 port map( A => ADD_RD2(0), ZN => n25266);
   U43 : NAND2_X1 port map( A1 => n25268, A2 => n25266, ZN => n1520);
   U44 : INV_X1 port map( A => n1520, ZN => n11227);
   U45 : INV_X1 port map( A => ADD_RD1(1), ZN => n25184);
   U46 : INV_X1 port map( A => ADD_RD1(2), ZN => n25186);
   U47 : OR3_X1 port map( A1 => n25184, A2 => n25186, A3 => ADD_RD1(0), ZN => 
                           n25157);
   U48 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), A3 => n25184, ZN
                           => n11230);
   U49 : INV_X1 port map( A => n11230, ZN => n1519);
   U50 : NAND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n25183);
   U51 : NOR2_X1 port map( A1 => n25186, A2 => n25183, ZN => n11225);
   U52 : INV_X1 port map( A => n11225, ZN => n1516);
   U53 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => n25183, ZN => n11232);
   U54 : INV_X1 port map( A => n11232, ZN => n1514);
   U55 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(1), A3 => ADD_RD1(0)
                           , ZN => n11231);
   U56 : INV_X1 port map( A => n11231, ZN => n1518);
   U57 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n25184, ZN => n25185);
   U58 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => n25185, ZN => n11228);
   U59 : INV_X1 port map( A => n11228, ZN => n1515);
   U60 : NOR2_X1 port map( A1 => n25186, A2 => n25185, ZN => n11229);
   U61 : INV_X1 port map( A => n11229, ZN => n1517);
   U62 : INV_X1 port map( A => ADD_RD2(1), ZN => n25269);
   U63 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n25269, ZN
                           => n11226);
   U64 : INV_X1 port map( A => n11226, ZN => n1521);
   U65 : INV_X1 port map( A => ADD_WR(3), ZN => n1513);
   U66 : INV_X1 port map( A => ADD_WR(4), ZN => n1512);
   U67 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20462, ZN => n25206);
   U68 : OAI22_X1 port map( A1 => n18353, A2 => n25206, B1 => n20428, B2 => 
                           n25215, ZN => n13469);
   U69 : OAI22_X1 port map( A1 => n18354, A2 => n25206, B1 => n20427, B2 => 
                           n25217, ZN => n13470);
   U70 : OAI22_X1 port map( A1 => n18349, A2 => n25206, B1 => n20426, B2 => 
                           n25219, ZN => n13471);
   U71 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20455, ZN => n25210);
   U72 : OAI22_X1 port map( A1 => n18359, A2 => n25210, B1 => n20425, B2 => 
                           n25194, ZN => n13472);
   U73 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20457, ZN => n25203);
   U74 : OAI22_X1 port map( A1 => n18360, A2 => n25203, B1 => n20424, B2 => 
                           n25193, ZN => n13473);
   U75 : OAI22_X1 port map( A1 => n18359, A2 => n25205, B1 => n20423, B2 => 
                           n25194, ZN => n13474);
   U76 : OAI22_X1 port map( A1 => n18360, A2 => n25205, B1 => n20422, B2 => 
                           n25193, ZN => n13475);
   U77 : OAI22_X1 port map( A1 => n18357, A2 => n25206, B1 => n20421, B2 => 
                           n25220, ZN => n13476);
   U78 : OAI22_X1 port map( A1 => n18359, A2 => n25206, B1 => n20420, B2 => 
                           n25194, ZN => n13477);
   U79 : OAI22_X1 port map( A1 => n18351, A2 => n25206, B1 => n20419, B2 => 
                           n25218, ZN => n13478);
   U80 : OAI22_X1 port map( A1 => n18355, A2 => n25206, B1 => n20418, B2 => 
                           n25221, ZN => n13479);
   U81 : OAI22_X1 port map( A1 => n18360, A2 => n25210, B1 => n20417, B2 => 
                           n25193, ZN => n13480);
   U82 : OAI22_X1 port map( A1 => n18359, A2 => n25203, B1 => n20416, B2 => 
                           n25194, ZN => n13481);
   U83 : OAI22_X1 port map( A1 => n18360, A2 => n25206, B1 => n20415, B2 => 
                           n25193, ZN => n13482);
   U84 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20446, ZN => n25204);
   U85 : OAI22_X1 port map( A1 => n18325, A2 => n25204, B1 => n20414, B2 => 
                           n25190, ZN => n13483);
   U86 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20448, ZN => n25209);
   U87 : OAI22_X1 port map( A1 => n18325, A2 => n25209, B1 => n20413, B2 => 
                           n25190, ZN => n13484);
   U88 : OAI22_X1 port map( A1 => n18329, A2 => n25210, B1 => n20412, B2 => 
                           n25192, ZN => n13485);
   U89 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20449, ZN => n25196);
   U90 : OAI22_X1 port map( A1 => n18325, A2 => n25196, B1 => n20411, B2 => 
                           n25190, ZN => n13486);
   U91 : OAI22_X1 port map( A1 => n18329, A2 => n25203, B1 => n20410, B2 => 
                           n25192, ZN => n13487);
   U92 : OAI22_X1 port map( A1 => n18329, A2 => n25205, B1 => n20409, B2 => 
                           n25192, ZN => n13488);
   U93 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20450, ZN => n25197);
   U94 : OAI22_X1 port map( A1 => n18325, A2 => n25197, B1 => n20408, B2 => 
                           n25190, ZN => n13489);
   U95 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20445, ZN => n25198);
   U96 : OAI22_X1 port map( A1 => n18325, A2 => n25198, B1 => n20407, B2 => 
                           n25190, ZN => n13490);
   U97 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20452, ZN => n25207);
   U98 : OAI22_X1 port map( A1 => n18325, A2 => n25207, B1 => n20406, B2 => 
                           n25190, ZN => n13491);
   U99 : OAI22_X1 port map( A1 => n18325, A2 => n25210, B1 => n20405, B2 => 
                           n25190, ZN => n13492);
   U100 : OAI22_X1 port map( A1 => n18325, A2 => n25203, B1 => n20404, B2 => 
                           n25190, ZN => n13493);
   U101 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20439, ZN => n25195);
   U102 : OAI22_X1 port map( A1 => n18330, A2 => n25195, B1 => n20403, B2 => 
                           n25188, ZN => n13494);
   U103 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20440, ZN => n25202);
   U104 : OAI22_X1 port map( A1 => n18330, A2 => n25202, B1 => n20402, B2 => 
                           n25188, ZN => n13495);
   U105 : OAI22_X1 port map( A1 => n18330, A2 => n25201, B1 => n20401, B2 => 
                           n25188, ZN => n13496);
   U106 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20443, ZN => n25200);
   U107 : OAI22_X1 port map( A1 => n18330, A2 => n25200, B1 => n20400, B2 => 
                           n25188, ZN => n13497);
   U108 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20444, ZN => n25199);
   U109 : OAI22_X1 port map( A1 => n18330, A2 => n25199, B1 => n20399, B2 => 
                           n25188, ZN => n13498);
   U110 : OAI22_X1 port map( A1 => n18330, A2 => n25198, B1 => n20398, B2 => 
                           n25188, ZN => n13499);
   U111 : OAI22_X1 port map( A1 => n18325, A2 => n25205, B1 => n20397, B2 => 
                           n25190, ZN => n13500);
   U112 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20447, ZN => n25211);
   U113 : OAI22_X1 port map( A1 => n18329, A2 => n25211, B1 => n20396, B2 => 
                           n25192, ZN => n13501);
   U114 : OAI22_X1 port map( A1 => n18327, A2 => n25209, B1 => n20395, B2 => 
                           n25191, ZN => n13502);
   U115 : OAI22_X1 port map( A1 => n18330, A2 => n25204, B1 => n20394, B2 => 
                           n25188, ZN => n13503);
   U116 : OAI22_X1 port map( A1 => n18330, A2 => n25211, B1 => n20393, B2 => 
                           n25188, ZN => n13504);
   U117 : OAI22_X1 port map( A1 => n18330, A2 => n25209, B1 => n20392, B2 => 
                           n25188, ZN => n13505);
   U118 : OAI22_X1 port map( A1 => n18330, A2 => n25196, B1 => n20391, B2 => 
                           n25188, ZN => n13506);
   U119 : OAI22_X1 port map( A1 => n18330, A2 => n25197, B1 => n20390, B2 => 
                           n25188, ZN => n13507);
   U120 : OAI22_X1 port map( A1 => n18329, A2 => n25204, B1 => n20389, B2 => 
                           n25192, ZN => n13508);
   U121 : OAI22_X1 port map( A1 => n18329, A2 => n25209, B1 => n20388, B2 => 
                           n25192, ZN => n13509);
   U122 : OAI22_X1 port map( A1 => n18329, A2 => n25198, B1 => n20387, B2 => 
                           n25192, ZN => n13510);
   U123 : OAI22_X1 port map( A1 => n18330, A2 => n25207, B1 => n20386, B2 => 
                           n25188, ZN => n13511);
   U124 : OAI22_X1 port map( A1 => n18329, A2 => n25199, B1 => n20385, B2 => 
                           n25192, ZN => n13512);
   U125 : OAI22_X1 port map( A1 => n18329, A2 => n25200, B1 => n20384, B2 => 
                           n25192, ZN => n13513);
   U126 : OAI22_X1 port map( A1 => n18329, A2 => n25201, B1 => n20383, B2 => 
                           n25192, ZN => n13514);
   U127 : OAI22_X1 port map( A1 => n18329, A2 => n25196, B1 => n20382, B2 => 
                           n25192, ZN => n13515);
   U128 : OAI22_X1 port map( A1 => n18329, A2 => n25202, B1 => n20381, B2 => 
                           n25192, ZN => n13516);
   U129 : OAI22_X1 port map( A1 => n18326, A2 => n25195, B1 => n20380, B2 => 
                           n25189, ZN => n13517);
   U130 : OAI22_X1 port map( A1 => n18326, A2 => n25202, B1 => n20379, B2 => 
                           n25189, ZN => n13518);
   U131 : OAI22_X1 port map( A1 => n18329, A2 => n25197, B1 => n20378, B2 => 
                           n25192, ZN => n13519);
   U132 : OAI22_X1 port map( A1 => n18326, A2 => n25201, B1 => n20377, B2 => 
                           n25189, ZN => n13520);
   U133 : OAI22_X1 port map( A1 => n18326, A2 => n25200, B1 => n20376, B2 => 
                           n25189, ZN => n13521);
   U134 : OAI22_X1 port map( A1 => n18329, A2 => n25207, B1 => n20375, B2 => 
                           n25192, ZN => n13522);
   U135 : OAI22_X1 port map( A1 => n18326, A2 => n25199, B1 => n20374, B2 => 
                           n25189, ZN => n13523);
   U136 : OAI22_X1 port map( A1 => n18326, A2 => n25198, B1 => n20373, B2 => 
                           n25189, ZN => n13524);
   U137 : OAI22_X1 port map( A1 => n18329, A2 => n25195, B1 => n20372, B2 => 
                           n25192, ZN => n13525);
   U138 : OAI22_X1 port map( A1 => n18328, A2 => n25205, B1 => n20371, B2 => 
                           n25187, ZN => n13526);
   U139 : OAI22_X1 port map( A1 => n18328, A2 => n25203, B1 => n20370, B2 => 
                           n25187, ZN => n13527);
   U140 : OAI22_X1 port map( A1 => n18328, A2 => n25210, B1 => n20369, B2 => 
                           n25187, ZN => n13528);
   U141 : OAI22_X1 port map( A1 => n18328, A2 => n25207, B1 => n20368, B2 => 
                           n25187, ZN => n13529);
   U142 : OAI22_X1 port map( A1 => n18328, A2 => n25197, B1 => n20367, B2 => 
                           n25187, ZN => n13530);
   U143 : OAI22_X1 port map( A1 => n18328, A2 => n25196, B1 => n20366, B2 => 
                           n25187, ZN => n13531);
   U144 : OAI22_X1 port map( A1 => n18326, A2 => n25204, B1 => n20365, B2 => 
                           n25189, ZN => n13532);
   U145 : OAI22_X1 port map( A1 => n18326, A2 => n25211, B1 => n20364, B2 => 
                           n25189, ZN => n13533);
   U146 : OAI22_X1 port map( A1 => n18326, A2 => n25209, B1 => n20363, B2 => 
                           n25189, ZN => n13534);
   U147 : OAI22_X1 port map( A1 => n18325, A2 => n25211, B1 => n20362, B2 => 
                           n25190, ZN => n13535);
   U148 : OAI22_X1 port map( A1 => n18326, A2 => n25196, B1 => n20361, B2 => 
                           n25189, ZN => n13536);
   U149 : OAI22_X1 port map( A1 => n18327, A2 => n25195, B1 => n20360, B2 => 
                           n25191, ZN => n13537);
   U150 : OAI22_X1 port map( A1 => n18326, A2 => n25197, B1 => n20359, B2 => 
                           n25189, ZN => n13538);
   U151 : OAI22_X1 port map( A1 => n18328, A2 => n25201, B1 => n20358, B2 => 
                           n25187, ZN => n13539);
   U152 : OAI22_X1 port map( A1 => n18328, A2 => n25202, B1 => n20357, B2 => 
                           n25187, ZN => n13540);
   U153 : OAI22_X1 port map( A1 => n18328, A2 => n25209, B1 => n20356, B2 => 
                           n25187, ZN => n13541);
   U154 : OAI22_X1 port map( A1 => n18328, A2 => n25195, B1 => n20355, B2 => 
                           n25187, ZN => n13542);
   U155 : OAI22_X1 port map( A1 => n18328, A2 => n25211, B1 => n20354, B2 => 
                           n25187, ZN => n13543);
   U156 : OAI22_X1 port map( A1 => n18326, A2 => n25207, B1 => n20353, B2 => 
                           n25189, ZN => n13544);
   U157 : OAI22_X1 port map( A1 => n18328, A2 => n25204, B1 => n20352, B2 => 
                           n25187, ZN => n13545);
   U158 : OAI22_X1 port map( A1 => n18327, A2 => n25203, B1 => n20351, B2 => 
                           n25191, ZN => n13546);
   U159 : OAI22_X1 port map( A1 => n18328, A2 => n25198, B1 => n20350, B2 => 
                           n25187, ZN => n13547);
   U160 : OAI22_X1 port map( A1 => n18327, A2 => n25202, B1 => n20349, B2 => 
                           n25191, ZN => n13548);
   U161 : OAI22_X1 port map( A1 => n18328, A2 => n25199, B1 => n20348, B2 => 
                           n25187, ZN => n13549);
   U162 : OAI22_X1 port map( A1 => n18326, A2 => n25210, B1 => n20347, B2 => 
                           n25189, ZN => n13550);
   U163 : OAI22_X1 port map( A1 => n18327, A2 => n25200, B1 => n20346, B2 => 
                           n25191, ZN => n13551);
   U164 : OAI22_X1 port map( A1 => n18325, A2 => n25199, B1 => n20345, B2 => 
                           n25190, ZN => n13552);
   U165 : OAI22_X1 port map( A1 => n18326, A2 => n25205, B1 => n20344, B2 => 
                           n25189, ZN => n13553);
   U166 : OAI22_X1 port map( A1 => n18327, A2 => n25196, B1 => n20343, B2 => 
                           n25191, ZN => n13554);
   U167 : OAI22_X1 port map( A1 => n18325, A2 => n25200, B1 => n20342, B2 => 
                           n25190, ZN => n13555);
   U168 : OAI22_X1 port map( A1 => n18327, A2 => n25204, B1 => n20341, B2 => 
                           n25191, ZN => n13556);
   U169 : OAI22_X1 port map( A1 => n18327, A2 => n25197, B1 => n20340, B2 => 
                           n25191, ZN => n13557);
   U170 : OAI22_X1 port map( A1 => n18327, A2 => n25210, B1 => n20339, B2 => 
                           n25191, ZN => n13558);
   U171 : OAI22_X1 port map( A1 => n18325, A2 => n25201, B1 => n20338, B2 => 
                           n25190, ZN => n13559);
   U172 : OAI22_X1 port map( A1 => n18325, A2 => n25202, B1 => n20337, B2 => 
                           n25190, ZN => n13560);
   U173 : OAI22_X1 port map( A1 => n18327, A2 => n25211, B1 => n20336, B2 => 
                           n25191, ZN => n13561);
   U174 : OAI22_X1 port map( A1 => n18325, A2 => n25195, B1 => n20335, B2 => 
                           n25190, ZN => n13562);
   U175 : OAI22_X1 port map( A1 => n18328, A2 => n25200, B1 => n20334, B2 => 
                           n25187, ZN => n13563);
   U176 : OAI22_X1 port map( A1 => n18327, A2 => n25207, B1 => n20333, B2 => 
                           n25191, ZN => n13564);
   U177 : OAI22_X1 port map( A1 => n18326, A2 => n25203, B1 => n20332, B2 => 
                           n25189, ZN => n13565);
   U178 : OAI22_X1 port map( A1 => n18327, A2 => n25205, B1 => n20331, B2 => 
                           n25191, ZN => n13566);
   U179 : OAI22_X1 port map( A1 => n18327, A2 => n25201, B1 => n20330, B2 => 
                           n25191, ZN => n13567);
   U180 : OAI22_X1 port map( A1 => n18327, A2 => n25198, B1 => n20329, B2 => 
                           n25191, ZN => n13568);
   U181 : OAI22_X1 port map( A1 => n18327, A2 => n25199, B1 => n20328, B2 => 
                           n25191, ZN => n13569);
   U182 : OAI22_X1 port map( A1 => n18360, A2 => n25202, B1 => n20327, B2 => 
                           n25193, ZN => n13570);
   U183 : OAI22_X1 port map( A1 => n18355, A2 => n25202, B1 => n20326, B2 => 
                           n25221, ZN => n13571);
   U184 : OAI22_X1 port map( A1 => n18357, A2 => n25202, B1 => n20325, B2 => 
                           n25220, ZN => n13572);
   U185 : OAI22_X1 port map( A1 => n18354, A2 => n25202, B1 => n20324, B2 => 
                           n25217, ZN => n13573);
   U186 : OAI22_X1 port map( A1 => n18359, A2 => n25202, B1 => n20323, B2 => 
                           n25194, ZN => n13574);
   U187 : OAI22_X1 port map( A1 => n18353, A2 => n25202, B1 => n20322, B2 => 
                           n25215, ZN => n13575);
   U188 : OAI22_X1 port map( A1 => n18349, A2 => n25202, B1 => n20321, B2 => 
                           n25219, ZN => n13576);
   U189 : OAI22_X1 port map( A1 => n18351, A2 => n25202, B1 => n20320, B2 => 
                           n25218, ZN => n13577);
   U190 : OAI22_X1 port map( A1 => n18351, A2 => n25210, B1 => n20319, B2 => 
                           n25218, ZN => n13578);
   U191 : OAI22_X1 port map( A1 => n18353, A2 => n25210, B1 => n20318, B2 => 
                           n25215, ZN => n13579);
   U192 : OAI22_X1 port map( A1 => n18330, A2 => n25210, B1 => n20317, B2 => 
                           n25188, ZN => n13580);
   U193 : OAI22_X1 port map( A1 => n18355, A2 => n25210, B1 => n20316, B2 => 
                           n25221, ZN => n13581);
   U194 : OAI22_X1 port map( A1 => n18357, A2 => n25210, B1 => n20315, B2 => 
                           n25220, ZN => n13582);
   U195 : OAI22_X1 port map( A1 => n18349, A2 => n25210, B1 => n20314, B2 => 
                           n25219, ZN => n13583);
   U196 : OAI22_X1 port map( A1 => n18354, A2 => n25210, B1 => n20313, B2 => 
                           n25217, ZN => n13584);
   U197 : OAI22_X1 port map( A1 => n18349, A2 => n25195, B1 => n20312, B2 => 
                           n25219, ZN => n13585);
   U198 : OAI22_X1 port map( A1 => n18354, A2 => n25195, B1 => n20311, B2 => 
                           n25217, ZN => n13586);
   U199 : OAI22_X1 port map( A1 => n18357, A2 => n25195, B1 => n20310, B2 => 
                           n25220, ZN => n13587);
   U200 : OAI22_X1 port map( A1 => n18360, A2 => n25195, B1 => n20309, B2 => 
                           n25193, ZN => n13588);
   U201 : OAI22_X1 port map( A1 => n18359, A2 => n25195, B1 => n20308, B2 => 
                           n25194, ZN => n13589);
   U202 : OAI22_X1 port map( A1 => n18355, A2 => n25195, B1 => n20307, B2 => 
                           n25221, ZN => n13590);
   U203 : OAI22_X1 port map( A1 => n18353, A2 => n25195, B1 => n20306, B2 => 
                           n25215, ZN => n13591);
   U204 : OAI22_X1 port map( A1 => n18351, A2 => n25195, B1 => n20305, B2 => 
                           n25218, ZN => n13592);
   U205 : OAI22_X1 port map( A1 => n18349, A2 => n25205, B1 => n20304, B2 => 
                           n25219, ZN => n13593);
   U206 : OAI22_X1 port map( A1 => n18351, A2 => n25205, B1 => n20303, B2 => 
                           n25218, ZN => n13594);
   U207 : OAI22_X1 port map( A1 => n18353, A2 => n25205, B1 => n20302, B2 => 
                           n25215, ZN => n13595);
   U208 : OAI22_X1 port map( A1 => n18326, A2 => n25206, B1 => n20301, B2 => 
                           n25189, ZN => n13596);
   U209 : OAI22_X1 port map( A1 => n18354, A2 => n25205, B1 => n20300, B2 => 
                           n25217, ZN => n13597);
   U210 : CLKBUF_X1 port map( A => n25205, Z => n25212);
   U211 : OAI22_X1 port map( A1 => n18355, A2 => n25212, B1 => n20299, B2 => 
                           n25221, ZN => n13598);
   U212 : OAI22_X1 port map( A1 => n18357, A2 => n25205, B1 => n20298, B2 => 
                           n25220, ZN => n13599);
   U213 : OAI22_X1 port map( A1 => n18351, A2 => n25203, B1 => n20297, B2 => 
                           n25218, ZN => n13600);
   U214 : OAI22_X1 port map( A1 => n18349, A2 => n25203, B1 => n20296, B2 => 
                           n25219, ZN => n13601);
   U215 : OAI22_X1 port map( A1 => n18357, A2 => n25198, B1 => n20295, B2 => 
                           n25220, ZN => n13602);
   U216 : OAI22_X1 port map( A1 => n18359, A2 => n25198, B1 => n20294, B2 => 
                           n25194, ZN => n13603);
   U217 : OAI22_X1 port map( A1 => n18349, A2 => n25198, B1 => n20293, B2 => 
                           n25219, ZN => n13604);
   U218 : OAI22_X1 port map( A1 => n18351, A2 => n25198, B1 => n20292, B2 => 
                           n25218, ZN => n13605);
   U219 : OAI22_X1 port map( A1 => n18360, A2 => n25204, B1 => n20291, B2 => 
                           n25193, ZN => n13606);
   U220 : OAI22_X1 port map( A1 => n18353, A2 => n25198, B1 => n20290, B2 => 
                           n25215, ZN => n13607);
   U221 : OAI22_X1 port map( A1 => n18354, A2 => n25198, B1 => n20289, B2 => 
                           n25217, ZN => n13608);
   U222 : OAI22_X1 port map( A1 => n18355, A2 => n25198, B1 => n20288, B2 => 
                           n25221, ZN => n13609);
   U223 : OAI22_X1 port map( A1 => n18328, A2 => n25206, B1 => n20287, B2 => 
                           n25187, ZN => n13610);
   U224 : OAI22_X1 port map( A1 => n18357, A2 => n25203, B1 => n20286, B2 => 
                           n25220, ZN => n13611);
   U225 : OAI22_X1 port map( A1 => n18355, A2 => n25203, B1 => n20285, B2 => 
                           n25221, ZN => n13612);
   U226 : OAI22_X1 port map( A1 => n18354, A2 => n25203, B1 => n20284, B2 => 
                           n25217, ZN => n13613);
   U227 : OAI22_X1 port map( A1 => n18353, A2 => n25203, B1 => n20283, B2 => 
                           n25215, ZN => n13614);
   U228 : OAI22_X1 port map( A1 => n18329, A2 => n25206, B1 => n20282, B2 => 
                           n25192, ZN => n13615);
   U229 : OAI22_X1 port map( A1 => n18353, A2 => n25199, B1 => n20281, B2 => 
                           n25215, ZN => n13616);
   U230 : OAI22_X1 port map( A1 => n18351, A2 => n25199, B1 => n20280, B2 => 
                           n25218, ZN => n13617);
   U231 : OAI22_X1 port map( A1 => n18349, A2 => n25199, B1 => n20279, B2 => 
                           n25219, ZN => n13618);
   U232 : OAI22_X1 port map( A1 => n18327, A2 => n25206, B1 => n20278, B2 => 
                           n25191, ZN => n13619);
   U233 : OAI22_X1 port map( A1 => n18330, A2 => n25203, B1 => n20277, B2 => 
                           n25188, ZN => n13620);
   U234 : OAI22_X1 port map( A1 => n18330, A2 => n25205, B1 => n20276, B2 => 
                           n25188, ZN => n13621);
   U235 : OAI22_X1 port map( A1 => n18360, A2 => n25199, B1 => n20275, B2 => 
                           n25193, ZN => n13622);
   U236 : OAI22_X1 port map( A1 => n18359, A2 => n25199, B1 => n20274, B2 => 
                           n25194, ZN => n13623);
   U237 : OAI22_X1 port map( A1 => n18357, A2 => n25199, B1 => n20273, B2 => 
                           n25220, ZN => n13624);
   U238 : OAI22_X1 port map( A1 => n18355, A2 => n25199, B1 => n20272, B2 => 
                           n25221, ZN => n13625);
   U239 : OAI22_X1 port map( A1 => n18354, A2 => n25199, B1 => n20271, B2 => 
                           n25217, ZN => n13626);
   U240 : OAI22_X1 port map( A1 => n18351, A2 => n25200, B1 => n20270, B2 => 
                           n25218, ZN => n13627);
   U241 : OAI22_X1 port map( A1 => n18349, A2 => n25200, B1 => n20269, B2 => 
                           n25219, ZN => n13628);
   U242 : OAI22_X1 port map( A1 => n18360, A2 => n25196, B1 => n20268, B2 => 
                           n25193, ZN => n13629);
   U243 : OAI22_X1 port map( A1 => n18325, A2 => n25206, B1 => n20267, B2 => 
                           n25190, ZN => n13630);
   U244 : OAI22_X1 port map( A1 => n18360, A2 => n25200, B1 => n20266, B2 => 
                           n25193, ZN => n13631);
   U245 : OAI22_X1 port map( A1 => n18359, A2 => n25200, B1 => n20265, B2 => 
                           n25194, ZN => n13632);
   U246 : OAI22_X1 port map( A1 => n18357, A2 => n25200, B1 => n20264, B2 => 
                           n25220, ZN => n13633);
   U247 : OAI22_X1 port map( A1 => n18355, A2 => n25200, B1 => n20263, B2 => 
                           n25221, ZN => n13634);
   U248 : OAI22_X1 port map( A1 => n18354, A2 => n25200, B1 => n20262, B2 => 
                           n25217, ZN => n13635);
   U249 : OAI22_X1 port map( A1 => n18353, A2 => n25200, B1 => n20261, B2 => 
                           n25215, ZN => n13636);
   U250 : OAI22_X1 port map( A1 => n18360, A2 => n25209, B1 => n20260, B2 => 
                           n25193, ZN => n13637);
   U251 : OAI22_X1 port map( A1 => n18330, A2 => n25206, B1 => n20259, B2 => 
                           n25188, ZN => n13638);
   U252 : OAI22_X1 port map( A1 => n18349, A2 => n25201, B1 => n20258, B2 => 
                           n25219, ZN => n13639);
   U253 : OAI22_X1 port map( A1 => n18360, A2 => n25201, B1 => n20257, B2 => 
                           n25193, ZN => n13640);
   U254 : OAI22_X1 port map( A1 => n18359, A2 => n25201, B1 => n20256, B2 => 
                           n25194, ZN => n13641);
   U255 : OAI22_X1 port map( A1 => n18357, A2 => n25201, B1 => n20255, B2 => 
                           n25220, ZN => n13642);
   U256 : OAI22_X1 port map( A1 => n18355, A2 => n25201, B1 => n20254, B2 => 
                           n25221, ZN => n13643);
   U257 : OAI22_X1 port map( A1 => n18360, A2 => n25197, B1 => n20253, B2 => 
                           n25193, ZN => n13644);
   U258 : OAI22_X1 port map( A1 => n18354, A2 => n25201, B1 => n20252, B2 => 
                           n25217, ZN => n13645);
   U259 : OAI22_X1 port map( A1 => n18353, A2 => n25201, B1 => n20251, B2 => 
                           n25215, ZN => n13646);
   U260 : OAI22_X1 port map( A1 => n18359, A2 => n25211, B1 => n20250, B2 => 
                           n25194, ZN => n13647);
   U261 : OAI22_X1 port map( A1 => n18357, A2 => n25211, B1 => n20249, B2 => 
                           n25220, ZN => n13648);
   U262 : OAI22_X1 port map( A1 => n18355, A2 => n25211, B1 => n20248, B2 => 
                           n25221, ZN => n13649);
   U263 : OAI22_X1 port map( A1 => n18354, A2 => n25211, B1 => n20247, B2 => 
                           n25217, ZN => n13650);
   U264 : OAI22_X1 port map( A1 => n18353, A2 => n25211, B1 => n20246, B2 => 
                           n25215, ZN => n13651);
   U265 : OAI22_X1 port map( A1 => n18351, A2 => n25211, B1 => n20245, B2 => 
                           n25218, ZN => n13652);
   U266 : OAI22_X1 port map( A1 => n18351, A2 => n25201, B1 => n20244, B2 => 
                           n25218, ZN => n13653);
   U267 : OAI22_X1 port map( A1 => n18349, A2 => n25211, B1 => n20243, B2 => 
                           n25219, ZN => n13654);
   U268 : OAI22_X1 port map( A1 => n18360, A2 => n25207, B1 => n20242, B2 => 
                           n25193, ZN => n13655);
   U269 : OAI22_X1 port map( A1 => n18359, A2 => n25197, B1 => n20241, B2 => 
                           n25194, ZN => n13656);
   U270 : OAI22_X1 port map( A1 => n18359, A2 => n25207, B1 => n20240, B2 => 
                           n25194, ZN => n13657);
   U271 : OAI22_X1 port map( A1 => n18357, A2 => n25207, B1 => n20239, B2 => 
                           n25220, ZN => n13658);
   U272 : OAI22_X1 port map( A1 => n18354, A2 => n25197, B1 => n20238, B2 => 
                           n25217, ZN => n13659);
   U273 : OAI22_X1 port map( A1 => n18355, A2 => n25207, B1 => n20237, B2 => 
                           n25221, ZN => n13660);
   U274 : OAI22_X1 port map( A1 => n18354, A2 => n25207, B1 => n20236, B2 => 
                           n25217, ZN => n13661);
   U275 : OAI22_X1 port map( A1 => n18353, A2 => n25207, B1 => n20235, B2 => 
                           n25215, ZN => n13662);
   U276 : OAI22_X1 port map( A1 => n18351, A2 => n25207, B1 => n20234, B2 => 
                           n25218, ZN => n13663);
   U277 : OAI22_X1 port map( A1 => n18349, A2 => n25207, B1 => n20233, B2 => 
                           n25219, ZN => n13664);
   U278 : OAI22_X1 port map( A1 => n18359, A2 => n25196, B1 => n20232, B2 => 
                           n25194, ZN => n13665);
   U279 : OAI22_X1 port map( A1 => n18357, A2 => n25196, B1 => n20231, B2 => 
                           n25220, ZN => n13666);
   U280 : OAI22_X1 port map( A1 => n18355, A2 => n25196, B1 => n20230, B2 => 
                           n25221, ZN => n13667);
   U281 : OAI22_X1 port map( A1 => n18354, A2 => n25196, B1 => n20229, B2 => 
                           n25217, ZN => n13668);
   U282 : OAI22_X1 port map( A1 => n18353, A2 => n25196, B1 => n20228, B2 => 
                           n25215, ZN => n13669);
   U283 : OAI22_X1 port map( A1 => n18351, A2 => n25196, B1 => n20227, B2 => 
                           n25218, ZN => n13670);
   U284 : OAI22_X1 port map( A1 => n18349, A2 => n25196, B1 => n20226, B2 => 
                           n25219, ZN => n13671);
   U285 : OAI22_X1 port map( A1 => n18357, A2 => n25197, B1 => n20225, B2 => 
                           n25220, ZN => n13672);
   U286 : OAI22_X1 port map( A1 => n18355, A2 => n25197, B1 => n20224, B2 => 
                           n25221, ZN => n13673);
   U287 : OAI22_X1 port map( A1 => n18349, A2 => n25197, B1 => n20223, B2 => 
                           n25219, ZN => n13674);
   U288 : OAI22_X1 port map( A1 => n18353, A2 => n25197, B1 => n20222, B2 => 
                           n25215, ZN => n13675);
   U289 : OAI22_X1 port map( A1 => n18351, A2 => n25197, B1 => n20221, B2 => 
                           n25218, ZN => n13676);
   U290 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20431, ZN => n25237);
   U291 : OAI22_X1 port map( A1 => n18330, A2 => n25237, B1 => n20220, B2 => 
                           n25188, ZN => n13677);
   U292 : OAI22_X1 port map( A1 => n18326, A2 => n25237, B1 => n20219, B2 => 
                           n25189, ZN => n13678);
   U293 : OAI22_X1 port map( A1 => n18327, A2 => n25237, B1 => n20218, B2 => 
                           n25191, ZN => n13679);
   U294 : OAI22_X1 port map( A1 => n18329, A2 => n25237, B1 => n20217, B2 => 
                           n25192, ZN => n13680);
   U295 : OAI22_X1 port map( A1 => n18325, A2 => n25237, B1 => n20216, B2 => 
                           n25190, ZN => n13681);
   U296 : OAI22_X1 port map( A1 => n18328, A2 => n25237, B1 => n20215, B2 => 
                           n25187, ZN => n13682);
   U297 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20436, ZN => n25250);
   U298 : OAI22_X1 port map( A1 => n18353, A2 => n25250, B1 => n20214, B2 => 
                           n25215, ZN => n13683);
   U299 : OAI22_X1 port map( A1 => n18354, A2 => n25250, B1 => n20213, B2 => 
                           n25217, ZN => n13684);
   U300 : OAI22_X1 port map( A1 => n18351, A2 => n25250, B1 => n20212, B2 => 
                           n25218, ZN => n13685);
   U301 : OAI22_X1 port map( A1 => n18355, A2 => n25250, B1 => n20211, B2 => 
                           n25221, ZN => n13686);
   U302 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20437, ZN => n25251);
   U303 : OAI22_X1 port map( A1 => n18355, A2 => n25251, B1 => n20210, B2 => 
                           n25221, ZN => n13687);
   U304 : OAI22_X1 port map( A1 => n18354, A2 => n25251, B1 => n20209, B2 => 
                           n25217, ZN => n13688);
   U305 : OAI22_X1 port map( A1 => n18355, A2 => n25204, B1 => n20208, B2 => 
                           n25221, ZN => n13689);
   U306 : OAI22_X1 port map( A1 => n18353, A2 => n25251, B1 => n20207, B2 => 
                           n25215, ZN => n13690);
   U307 : OAI22_X1 port map( A1 => n18351, A2 => n25251, B1 => n20206, B2 => 
                           n25218, ZN => n13691);
   U308 : OAI22_X1 port map( A1 => n18349, A2 => n25251, B1 => n20205, B2 => 
                           n25219, ZN => n13692);
   U309 : OAI22_X1 port map( A1 => n18349, A2 => n25250, B1 => n20204, B2 => 
                           n25219, ZN => n13693);
   U310 : OAI22_X1 port map( A1 => n18349, A2 => n25204, B1 => n20203, B2 => 
                           n25219, ZN => n13694);
   U311 : OAI22_X1 port map( A1 => n18351, A2 => n25204, B1 => n20202, B2 => 
                           n25218, ZN => n13695);
   U312 : OAI22_X1 port map( A1 => n18357, A2 => n25250, B1 => n20201, B2 => 
                           n25220, ZN => n13696);
   U313 : OAI22_X1 port map( A1 => n18357, A2 => n25251, B1 => n20200, B2 => 
                           n25220, ZN => n13697);
   U314 : OAI22_X1 port map( A1 => n18353, A2 => n25204, B1 => n20199, B2 => 
                           n25215, ZN => n13698);
   U315 : OAI22_X1 port map( A1 => n18354, A2 => n25204, B1 => n20198, B2 => 
                           n25217, ZN => n13699);
   U316 : OAI22_X1 port map( A1 => n18357, A2 => n25204, B1 => n20197, B2 => 
                           n25220, ZN => n13700);
   U317 : OAI22_X1 port map( A1 => n18360, A2 => n25250, B1 => n20196, B2 => 
                           n25193, ZN => n13701);
   U318 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20434, ZN => n25247);
   U319 : OAI22_X1 port map( A1 => n18355, A2 => n25247, B1 => n20195, B2 => 
                           n25221, ZN => n13702);
   U320 : OAI22_X1 port map( A1 => n18357, A2 => n25247, B1 => n20194, B2 => 
                           n25220, ZN => n13703);
   U321 : OAI22_X1 port map( A1 => n18359, A2 => n25250, B1 => n20193, B2 => 
                           n25194, ZN => n13704);
   U322 : OAI22_X1 port map( A1 => n18359, A2 => n25251, B1 => n20192, B2 => 
                           n25194, ZN => n13705);
   U323 : OAI22_X1 port map( A1 => n18359, A2 => n25247, B1 => n20191, B2 => 
                           n25194, ZN => n13706);
   U324 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20435, ZN => n25248);
   U325 : OAI22_X1 port map( A1 => n18351, A2 => n25248, B1 => n20190, B2 => 
                           n25218, ZN => n13707);
   U326 : OAI22_X1 port map( A1 => n18353, A2 => n25248, B1 => n20189, B2 => 
                           n25215, ZN => n13708);
   U327 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20433, ZN => n25249);
   U328 : OAI22_X1 port map( A1 => n18351, A2 => n25249, B1 => n20188, B2 => 
                           n25218, ZN => n13709);
   U329 : OAI22_X1 port map( A1 => n18349, A2 => n25249, B1 => n20187, B2 => 
                           n25219, ZN => n13710);
   U330 : OAI22_X1 port map( A1 => n18359, A2 => n25204, B1 => n20186, B2 => 
                           n25194, ZN => n13711);
   U331 : OAI22_X1 port map( A1 => n18360, A2 => n25248, B1 => n20185, B2 => 
                           n25193, ZN => n13712);
   U332 : OAI22_X1 port map( A1 => n18359, A2 => n25249, B1 => n20184, B2 => 
                           n25194, ZN => n13713);
   U333 : OAI22_X1 port map( A1 => n18349, A2 => n25247, B1 => n20183, B2 => 
                           n25219, ZN => n13714);
   U334 : OAI22_X1 port map( A1 => n18351, A2 => n25247, B1 => n20182, B2 => 
                           n25218, ZN => n13715);
   U335 : OAI22_X1 port map( A1 => n18353, A2 => n25247, B1 => n20181, B2 => 
                           n25215, ZN => n13716);
   U336 : OAI22_X1 port map( A1 => n18354, A2 => n25247, B1 => n20180, B2 => 
                           n25217, ZN => n13717);
   U337 : OAI22_X1 port map( A1 => n18357, A2 => n25248, B1 => n20179, B2 => 
                           n25220, ZN => n13718);
   U338 : OAI22_X1 port map( A1 => n18359, A2 => n25248, B1 => n20178, B2 => 
                           n25194, ZN => n13719);
   U339 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20432, ZN => n25246);
   U340 : OAI22_X1 port map( A1 => n18351, A2 => n25246, B1 => n20177, B2 => 
                           n25218, ZN => n13720);
   U341 : OAI22_X1 port map( A1 => n18357, A2 => n25249, B1 => n20176, B2 => 
                           n25220, ZN => n13721);
   U342 : OAI22_X1 port map( A1 => n18360, A2 => n25249, B1 => n20175, B2 => 
                           n25193, ZN => n13722);
   U343 : OAI22_X1 port map( A1 => n18360, A2 => n25247, B1 => n20174, B2 => 
                           n25193, ZN => n13723);
   U344 : OAI22_X1 port map( A1 => n18353, A2 => n25246, B1 => n20173, B2 => 
                           n25215, ZN => n13724);
   U345 : OAI22_X1 port map( A1 => n18354, A2 => n25248, B1 => n20172, B2 => 
                           n25217, ZN => n13725);
   U346 : OAI22_X1 port map( A1 => n18360, A2 => n25251, B1 => n20171, B2 => 
                           n25193, ZN => n13726);
   U347 : OAI22_X1 port map( A1 => n18354, A2 => n25246, B1 => n20170, B2 => 
                           n25217, ZN => n13727);
   U348 : OAI22_X1 port map( A1 => n18355, A2 => n25246, B1 => n20169, B2 => 
                           n25221, ZN => n13728);
   U349 : OAI22_X1 port map( A1 => n18357, A2 => n25246, B1 => n20168, B2 => 
                           n25220, ZN => n13729);
   U350 : OAI22_X1 port map( A1 => n18359, A2 => n25246, B1 => n20167, B2 => 
                           n25194, ZN => n13730);
   U351 : OAI22_X1 port map( A1 => n18355, A2 => n25249, B1 => n20166, B2 => 
                           n25221, ZN => n13731);
   U352 : OAI22_X1 port map( A1 => n18360, A2 => n25198, B1 => n20165, B2 => 
                           n25193, ZN => n13732);
   U353 : OAI22_X1 port map( A1 => n18354, A2 => n25249, B1 => n20164, B2 => 
                           n25217, ZN => n13733);
   U354 : OAI22_X1 port map( A1 => n18353, A2 => n25249, B1 => n20163, B2 => 
                           n25215, ZN => n13734);
   U355 : OAI22_X1 port map( A1 => n18349, A2 => n25248, B1 => n20162, B2 => 
                           n25219, ZN => n13735);
   U356 : OAI22_X1 port map( A1 => n18355, A2 => n25209, B1 => n20161, B2 => 
                           n25221, ZN => n13736);
   U357 : OAI22_X1 port map( A1 => n18349, A2 => n25246, B1 => n20160, B2 => 
                           n25219, ZN => n13737);
   U358 : OAI22_X1 port map( A1 => n18354, A2 => n25209, B1 => n20159, B2 => 
                           n25217, ZN => n13738);
   U359 : OAI22_X1 port map( A1 => n18355, A2 => n25248, B1 => n20158, B2 => 
                           n25221, ZN => n13739);
   U360 : OAI22_X1 port map( A1 => n18351, A2 => n25209, B1 => n20157, B2 => 
                           n25218, ZN => n13740);
   U361 : OAI22_X1 port map( A1 => n18360, A2 => n25211, B1 => n20156, B2 => 
                           n25193, ZN => n13741);
   U362 : OAI22_X1 port map( A1 => n18349, A2 => n25209, B1 => n20155, B2 => 
                           n25219, ZN => n13742);
   U363 : OAI22_X1 port map( A1 => n18360, A2 => n25246, B1 => n20154, B2 => 
                           n25193, ZN => n13743);
   U364 : OAI22_X1 port map( A1 => n18359, A2 => n25209, B1 => n20153, B2 => 
                           n25194, ZN => n13744);
   U365 : OAI22_X1 port map( A1 => n18357, A2 => n25209, B1 => n20152, B2 => 
                           n25220, ZN => n13745);
   U366 : OAI22_X1 port map( A1 => n18353, A2 => n25209, B1 => n20151, B2 => 
                           n25215, ZN => n13746);
   U367 : OAI22_X1 port map( A1 => n18357, A2 => n25237, B1 => n20150, B2 => 
                           n25220, ZN => n13747);
   U368 : OAI22_X1 port map( A1 => n18351, A2 => n25237, B1 => n20149, B2 => 
                           n25218, ZN => n13748);
   U369 : OAI22_X1 port map( A1 => n18360, A2 => n25237, B1 => n20148, B2 => 
                           n25193, ZN => n13749);
   U370 : OAI22_X1 port map( A1 => n18359, A2 => n25237, B1 => n20147, B2 => 
                           n25194, ZN => n13750);
   U371 : OAI22_X1 port map( A1 => n18355, A2 => n25237, B1 => n20146, B2 => 
                           n25221, ZN => n13751);
   U372 : OAI22_X1 port map( A1 => n18353, A2 => n25237, B1 => n20145, B2 => 
                           n25215, ZN => n13752);
   U373 : OAI22_X1 port map( A1 => n18354, A2 => n25237, B1 => n20144, B2 => 
                           n25217, ZN => n13753);
   U374 : OAI22_X1 port map( A1 => n18349, A2 => n25237, B1 => n20143, B2 => 
                           n25219, ZN => n13754);
   U375 : OAI22_X1 port map( A1 => n18327, A2 => n25247, B1 => n20142, B2 => 
                           n25191, ZN => n13755);
   U376 : OAI22_X1 port map( A1 => n18325, A2 => n25251, B1 => n20141, B2 => 
                           n25190, ZN => n13756);
   U377 : OAI22_X1 port map( A1 => n18326, A2 => n25246, B1 => n20140, B2 => 
                           n25189, ZN => n13757);
   U378 : OAI22_X1 port map( A1 => n18330, A2 => n25250, B1 => n20139, B2 => 
                           n25188, ZN => n13758);
   U379 : OAI22_X1 port map( A1 => n18325, A2 => n25250, B1 => n20138, B2 => 
                           n25190, ZN => n13759);
   U380 : OAI22_X1 port map( A1 => n18325, A2 => n25248, B1 => n20137, B2 => 
                           n25190, ZN => n13760);
   U381 : OAI22_X1 port map( A1 => n18325, A2 => n25247, B1 => n20136, B2 => 
                           n25190, ZN => n13761);
   U382 : OAI22_X1 port map( A1 => n18325, A2 => n25249, B1 => n20135, B2 => 
                           n25190, ZN => n13762);
   U383 : OAI22_X1 port map( A1 => n18330, A2 => n25246, B1 => n20134, B2 => 
                           n25188, ZN => n13763);
   U384 : OAI22_X1 port map( A1 => n18325, A2 => n25246, B1 => n20133, B2 => 
                           n25190, ZN => n13764);
   U385 : OAI22_X1 port map( A1 => n18327, A2 => n25251, B1 => n20132, B2 => 
                           n25191, ZN => n13765);
   U386 : OAI22_X1 port map( A1 => n18328, A2 => n25251, B1 => n20131, B2 => 
                           n25187, ZN => n13766);
   U387 : OAI22_X1 port map( A1 => n18326, A2 => n25249, B1 => n20130, B2 => 
                           n25189, ZN => n13767);
   U388 : OAI22_X1 port map( A1 => n18327, A2 => n25246, B1 => n20129, B2 => 
                           n25191, ZN => n13768);
   U389 : OAI22_X1 port map( A1 => n18327, A2 => n25249, B1 => n20128, B2 => 
                           n25191, ZN => n13769);
   U390 : OAI22_X1 port map( A1 => n18326, A2 => n25247, B1 => n20127, B2 => 
                           n25189, ZN => n13770);
   U391 : OAI22_X1 port map( A1 => n18328, A2 => n25246, B1 => n20126, B2 => 
                           n25187, ZN => n13771);
   U392 : OAI22_X1 port map( A1 => n18326, A2 => n25248, B1 => n20125, B2 => 
                           n25189, ZN => n13772);
   U393 : OAI22_X1 port map( A1 => n18326, A2 => n25250, B1 => n20124, B2 => 
                           n25189, ZN => n13773);
   U394 : OAI22_X1 port map( A1 => n18326, A2 => n25251, B1 => n20123, B2 => 
                           n25189, ZN => n13774);
   U395 : OAI22_X1 port map( A1 => n18328, A2 => n25248, B1 => n20122, B2 => 
                           n25187, ZN => n13775);
   U396 : OAI22_X1 port map( A1 => n18328, A2 => n25250, B1 => n20121, B2 => 
                           n25187, ZN => n13776);
   U397 : OAI22_X1 port map( A1 => n18329, A2 => n25248, B1 => n20120, B2 => 
                           n25192, ZN => n13777);
   U398 : OAI22_X1 port map( A1 => n18327, A2 => n25250, B1 => n20119, B2 => 
                           n25191, ZN => n13778);
   U399 : OAI22_X1 port map( A1 => n18329, A2 => n25249, B1 => n20118, B2 => 
                           n25192, ZN => n13779);
   U400 : OAI22_X1 port map( A1 => n18330, A2 => n25248, B1 => n20117, B2 => 
                           n25188, ZN => n13780);
   U401 : OAI22_X1 port map( A1 => n18327, A2 => n25248, B1 => n20116, B2 => 
                           n25191, ZN => n13781);
   U402 : OAI22_X1 port map( A1 => n18330, A2 => n25251, B1 => n20115, B2 => 
                           n25188, ZN => n13782);
   U403 : OAI22_X1 port map( A1 => n18329, A2 => n25247, B1 => n20114, B2 => 
                           n25192, ZN => n13783);
   U404 : OAI22_X1 port map( A1 => n18329, A2 => n25251, B1 => n20113, B2 => 
                           n25192, ZN => n13784);
   U405 : OAI22_X1 port map( A1 => n18330, A2 => n25249, B1 => n20112, B2 => 
                           n25188, ZN => n13785);
   U406 : OAI22_X1 port map( A1 => n18330, A2 => n25247, B1 => n20111, B2 => 
                           n25188, ZN => n13786);
   U407 : OAI22_X1 port map( A1 => n18329, A2 => n25250, B1 => n20110, B2 => 
                           n25192, ZN => n13787);
   U408 : OAI22_X1 port map( A1 => n18329, A2 => n25246, B1 => n20109, B2 => 
                           n25192, ZN => n13788);
   U409 : OAI22_X1 port map( A1 => n18328, A2 => n25247, B1 => n20108, B2 => 
                           n25187, ZN => n13789);
   U410 : OAI22_X1 port map( A1 => n18328, A2 => n25249, B1 => n20107, B2 => 
                           n25187, ZN => n13790);
   U411 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20441, ZN => n25216);
   U412 : OAI22_X1 port map( A1 => n18330, A2 => n25216, B1 => n20106, B2 => 
                           n25188, ZN => n13791);
   U413 : OAI22_X1 port map( A1 => n18326, A2 => n25216, B1 => n20105, B2 => 
                           n25189, ZN => n13792);
   U414 : OAI22_X1 port map( A1 => n18325, A2 => n25216, B1 => n20104, B2 => 
                           n25190, ZN => n13793);
   U415 : OAI22_X1 port map( A1 => n18329, A2 => n25216, B1 => n20103, B2 => 
                           n25192, ZN => n13794);
   U416 : OAI22_X1 port map( A1 => n18327, A2 => n25216, B1 => n20102, B2 => 
                           n25191, ZN => n13795);
   U417 : OAI22_X1 port map( A1 => n18328, A2 => n25216, B1 => n20101, B2 => 
                           n25187, ZN => n13796);
   U418 : OAI22_X1 port map( A1 => n18348, A2 => n25206, B1 => n20100, B2 => 
                           n25234, ZN => n13797);
   U419 : OAI22_X1 port map( A1 => n18347, A2 => n25210, B1 => n20099, B2 => 
                           n25232, ZN => n13798);
   U420 : OAI22_X1 port map( A1 => n18348, A2 => n25202, B1 => n20098, B2 => 
                           n25234, ZN => n13799);
   U421 : OAI22_X1 port map( A1 => n18346, A2 => n25216, B1 => n20097, B2 => 
                           n25233, ZN => n13800);
   U422 : OAI22_X1 port map( A1 => n18348, A2 => n25196, B1 => n20096, B2 => 
                           n25234, ZN => n13801);
   U423 : OAI22_X1 port map( A1 => n18346, A2 => n25199, B1 => n20095, B2 => 
                           n25233, ZN => n13802);
   U424 : OAI22_X1 port map( A1 => n18348, A2 => n25205, B1 => n20094, B2 => 
                           n25234, ZN => n13803);
   U425 : OAI22_X1 port map( A1 => n18346, A2 => n25205, B1 => n20093, B2 => 
                           n25233, ZN => n13804);
   U426 : OAI22_X1 port map( A1 => n18346, A2 => n25195, B1 => n20092, B2 => 
                           n25233, ZN => n13805);
   U427 : OAI22_X1 port map( A1 => n18348, A2 => n25203, B1 => n20091, B2 => 
                           n25234, ZN => n13806);
   U428 : OAI22_X1 port map( A1 => n18347, A2 => n25201, B1 => n20090, B2 => 
                           n25232, ZN => n13807);
   U429 : OAI22_X1 port map( A1 => n18346, A2 => n25202, B1 => n20089, B2 => 
                           n25233, ZN => n13808);
   U430 : OAI22_X1 port map( A1 => n18347, A2 => n25199, B1 => n20088, B2 => 
                           n25232, ZN => n13809);
   U431 : OAI22_X1 port map( A1 => n18346, A2 => n25201, B1 => n20087, B2 => 
                           n25233, ZN => n13810);
   U432 : OAI22_X1 port map( A1 => n18346, A2 => n25200, B1 => n20086, B2 => 
                           n25233, ZN => n13811);
   U433 : OAI22_X1 port map( A1 => n18348, A2 => n25207, B1 => n20085, B2 => 
                           n25234, ZN => n13812);
   U434 : OAI22_X1 port map( A1 => n18348, A2 => n25211, B1 => n20084, B2 => 
                           n25234, ZN => n13813);
   U435 : OAI22_X1 port map( A1 => n18347, A2 => n25205, B1 => n20083, B2 => 
                           n25232, ZN => n13814);
   U436 : OAI22_X1 port map( A1 => n18346, A2 => n25198, B1 => n20082, B2 => 
                           n25233, ZN => n13815);
   U437 : OAI22_X1 port map( A1 => n18347, A2 => n25206, B1 => n20081, B2 => 
                           n25232, ZN => n13816);
   U438 : OAI22_X1 port map( A1 => n18346, A2 => n25211, B1 => n20080, B2 => 
                           n25233, ZN => n13817);
   U439 : OAI22_X1 port map( A1 => n18348, A2 => n25210, B1 => n20079, B2 => 
                           n25234, ZN => n13818);
   U440 : OAI22_X1 port map( A1 => n18348, A2 => n25199, B1 => n20078, B2 => 
                           n25234, ZN => n13819);
   U441 : OAI22_X1 port map( A1 => n18348, A2 => n25197, B1 => n20077, B2 => 
                           n25234, ZN => n13820);
   U442 : OAI22_X1 port map( A1 => n18346, A2 => n25196, B1 => n20076, B2 => 
                           n25233, ZN => n13821);
   U443 : OAI22_X1 port map( A1 => n18346, A2 => n25197, B1 => n20075, B2 => 
                           n25233, ZN => n13822);
   U444 : OAI22_X1 port map( A1 => n18346, A2 => n25207, B1 => n20074, B2 => 
                           n25233, ZN => n13823);
   U445 : OAI22_X1 port map( A1 => n18348, A2 => n25216, B1 => n20073, B2 => 
                           n25234, ZN => n13824);
   U446 : OAI22_X1 port map( A1 => n18347, A2 => n25197, B1 => n20072, B2 => 
                           n25232, ZN => n13825);
   U447 : OAI22_X1 port map( A1 => n18346, A2 => n25210, B1 => n20071, B2 => 
                           n25233, ZN => n13826);
   U448 : OAI22_X1 port map( A1 => n18348, A2 => n25201, B1 => n20070, B2 => 
                           n25234, ZN => n13827);
   U449 : OAI22_X1 port map( A1 => n18346, A2 => n25203, B1 => n20069, B2 => 
                           n25233, ZN => n13828);
   U450 : OAI22_X1 port map( A1 => n18347, A2 => n25203, B1 => n20068, B2 => 
                           n25232, ZN => n13829);
   U451 : OAI22_X1 port map( A1 => n18347, A2 => n25211, B1 => n20067, B2 => 
                           n25232, ZN => n13830);
   U452 : OAI22_X1 port map( A1 => n18347, A2 => n25196, B1 => n20066, B2 => 
                           n25232, ZN => n13831);
   U453 : OAI22_X1 port map( A1 => n18348, A2 => n25195, B1 => n20065, B2 => 
                           n25234, ZN => n13832);
   U454 : OAI22_X1 port map( A1 => n18347, A2 => n25202, B1 => n20064, B2 => 
                           n25232, ZN => n13833);
   U455 : OAI22_X1 port map( A1 => n18347, A2 => n25216, B1 => n20063, B2 => 
                           n25232, ZN => n13834);
   U456 : OAI22_X1 port map( A1 => n18346, A2 => n25206, B1 => n20062, B2 => 
                           n25233, ZN => n13835);
   U457 : OAI22_X1 port map( A1 => n18348, A2 => n25198, B1 => n20061, B2 => 
                           n25234, ZN => n13836);
   U458 : OAI22_X1 port map( A1 => n18347, A2 => n25195, B1 => n20060, B2 => 
                           n25232, ZN => n13837);
   U459 : OAI22_X1 port map( A1 => n18347, A2 => n25198, B1 => n20059, B2 => 
                           n25232, ZN => n13838);
   U460 : OAI22_X1 port map( A1 => n18347, A2 => n25207, B1 => n20058, B2 => 
                           n25232, ZN => n13839);
   U461 : OAI22_X1 port map( A1 => n18348, A2 => n25200, B1 => n20057, B2 => 
                           n25234, ZN => n13840);
   U462 : OAI22_X1 port map( A1 => n18347, A2 => n25200, B1 => n20056, B2 => 
                           n25232, ZN => n13841);
   U463 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20438, ZN => n25253);
   U464 : OAI22_X1 port map( A1 => n18328, A2 => n25253, B1 => n20055, B2 => 
                           n25187, ZN => n13843);
   U465 : OAI22_X1 port map( A1 => n18330, A2 => n25253, B1 => n20054, B2 => 
                           n25188, ZN => n13845);
   U466 : OAI22_X1 port map( A1 => n18326, A2 => n25253, B1 => n20053, B2 => 
                           n25189, ZN => n13847);
   U467 : OAI22_X1 port map( A1 => n18325, A2 => n25253, B1 => n20052, B2 => 
                           n25190, ZN => n13849);
   U468 : OAI22_X1 port map( A1 => n18327, A2 => n25253, B1 => n20051, B2 => 
                           n25191, ZN => n13851);
   U469 : OAI22_X1 port map( A1 => n18329, A2 => n25253, B1 => n20050, B2 => 
                           n25192, ZN => n13853);
   U470 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20461, ZN => n25228);
   U471 : OAI22_X1 port map( A1 => n18348, A2 => n25228, B1 => n20049, B2 => 
                           n25234, ZN => n13854);
   U472 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20458, ZN => n25230);
   U473 : OAI22_X1 port map( A1 => n18348, A2 => n25230, B1 => n20048, B2 => 
                           n25234, ZN => n13855);
   U474 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20454, ZN => n25223);
   U475 : OAI22_X1 port map( A1 => n18329, A2 => n25223, B1 => n20047, B2 => 
                           n25192, ZN => n13856);
   U476 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20456, ZN => n25226);
   U477 : OAI22_X1 port map( A1 => n18348, A2 => n25226, B1 => n20046, B2 => 
                           n25234, ZN => n13857);
   U478 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20453, ZN => n25224);
   U479 : OAI22_X1 port map( A1 => n18329, A2 => n25224, B1 => n20045, B2 => 
                           n25192, ZN => n13858);
   U480 : OAI22_X1 port map( A1 => n18348, A2 => n25223, B1 => n20044, B2 => 
                           n25234, ZN => n13859);
   U481 : OAI22_X1 port map( A1 => n18348, A2 => n25224, B1 => n20043, B2 => 
                           n25234, ZN => n13860);
   U482 : OAI22_X1 port map( A1 => n18347, A2 => n25228, B1 => n20042, B2 => 
                           n25232, ZN => n13861);
   U483 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20459, ZN => n25229);
   U484 : OAI22_X1 port map( A1 => n18347, A2 => n25229, B1 => n20041, B2 => 
                           n25232, ZN => n13862);
   U485 : OAI22_X1 port map( A1 => n18347, A2 => n25230, B1 => n20040, B2 => 
                           n25232, ZN => n13863);
   U486 : OAI22_X1 port map( A1 => n18347, A2 => n25226, B1 => n20039, B2 => 
                           n25232, ZN => n13864);
   U487 : OAI22_X1 port map( A1 => n18347, A2 => n25223, B1 => n20038, B2 => 
                           n25232, ZN => n13865);
   U488 : OAI22_X1 port map( A1 => n18347, A2 => n25224, B1 => n20037, B2 => 
                           n25232, ZN => n13866);
   U489 : OAI22_X1 port map( A1 => n18330, A2 => n25223, B1 => n20036, B2 => 
                           n25188, ZN => n13867);
   U490 : OAI22_X1 port map( A1 => n18346, A2 => n25228, B1 => n20035, B2 => 
                           n25233, ZN => n13868);
   U491 : OAI22_X1 port map( A1 => n18346, A2 => n25229, B1 => n20034, B2 => 
                           n25233, ZN => n13869);
   U492 : OAI22_X1 port map( A1 => n18346, A2 => n25230, B1 => n20033, B2 => 
                           n25233, ZN => n13870);
   U493 : OAI22_X1 port map( A1 => n18346, A2 => n25226, B1 => n20032, B2 => 
                           n25233, ZN => n13871);
   U494 : OAI22_X1 port map( A1 => n18346, A2 => n25223, B1 => n20031, B2 => 
                           n25233, ZN => n13872);
   U495 : OAI22_X1 port map( A1 => n18346, A2 => n25224, B1 => n20030, B2 => 
                           n25233, ZN => n13873);
   U496 : OAI22_X1 port map( A1 => n18328, A2 => n25224, B1 => n20029, B2 => 
                           n25187, ZN => n13874);
   U497 : NAND2_X2 port map( A1 => RESET_BAR, A2 => n20451, ZN => n25222);
   U498 : OAI22_X1 port map( A1 => n18328, A2 => n25222, B1 => n20028, B2 => 
                           n25187, ZN => n13875);
   U499 : OAI22_X1 port map( A1 => n18327, A2 => n25228, B1 => n20027, B2 => 
                           n25191, ZN => n13876);
   U500 : OAI22_X1 port map( A1 => n18327, A2 => n25229, B1 => n20026, B2 => 
                           n25191, ZN => n13877);
   U501 : OAI22_X1 port map( A1 => n18327, A2 => n25230, B1 => n20025, B2 => 
                           n25191, ZN => n13878);
   U502 : OAI22_X1 port map( A1 => n18327, A2 => n25226, B1 => n20024, B2 => 
                           n25191, ZN => n13879);
   U503 : OAI22_X1 port map( A1 => n18360, A2 => n25228, B1 => n20023, B2 => 
                           n25193, ZN => n13880);
   U504 : OAI22_X1 port map( A1 => n18360, A2 => n25229, B1 => n20022, B2 => 
                           n25193, ZN => n13881);
   U505 : OAI22_X1 port map( A1 => n18360, A2 => n25230, B1 => n20021, B2 => 
                           n25193, ZN => n13882);
   U506 : OAI22_X1 port map( A1 => n18360, A2 => n25226, B1 => n20020, B2 => 
                           n25193, ZN => n13883);
   U507 : OAI22_X1 port map( A1 => n18348, A2 => n25229, B1 => n20019, B2 => 
                           n25234, ZN => n13884);
   U508 : OAI22_X1 port map( A1 => n18359, A2 => n25230, B1 => n20018, B2 => 
                           n25194, ZN => n13885);
   U509 : OAI22_X1 port map( A1 => n18330, A2 => n25224, B1 => n20017, B2 => 
                           n25188, ZN => n13886);
   U510 : OAI22_X1 port map( A1 => n18327, A2 => n25224, B1 => n20016, B2 => 
                           n25191, ZN => n13887);
   U511 : OAI22_X1 port map( A1 => n18330, A2 => n25222, B1 => n20015, B2 => 
                           n25188, ZN => n13888);
   U512 : OAI22_X1 port map( A1 => n18329, A2 => n25228, B1 => n20014, B2 => 
                           n25192, ZN => n13889);
   U513 : OAI22_X1 port map( A1 => n18329, A2 => n25229, B1 => n20013, B2 => 
                           n25192, ZN => n13890);
   U514 : OAI22_X1 port map( A1 => n18329, A2 => n25230, B1 => n20012, B2 => 
                           n25192, ZN => n13891);
   U515 : OAI22_X1 port map( A1 => n18329, A2 => n25226, B1 => n20011, B2 => 
                           n25192, ZN => n13892);
   U516 : OAI22_X1 port map( A1 => n18326, A2 => n25230, B1 => n20010, B2 => 
                           n25189, ZN => n13893);
   U517 : OAI22_X1 port map( A1 => n18326, A2 => n25226, B1 => n20009, B2 => 
                           n25189, ZN => n13894);
   U518 : OAI22_X1 port map( A1 => n18326, A2 => n25223, B1 => n20008, B2 => 
                           n25189, ZN => n13895);
   U519 : OAI22_X1 port map( A1 => n18326, A2 => n25224, B1 => n20007, B2 => 
                           n25189, ZN => n13896);
   U520 : OAI22_X1 port map( A1 => n18326, A2 => n25229, B1 => n20006, B2 => 
                           n25189, ZN => n13897);
   U521 : OAI22_X1 port map( A1 => n18328, A2 => n25229, B1 => n20005, B2 => 
                           n25187, ZN => n13898);
   U522 : OAI22_X1 port map( A1 => n18325, A2 => n25230, B1 => n20004, B2 => 
                           n25190, ZN => n13899);
   U523 : OAI22_X1 port map( A1 => n18329, A2 => n25222, B1 => n20003, B2 => 
                           n25192, ZN => n13901);
   U524 : OAI22_X1 port map( A1 => n18359, A2 => n25228, B1 => n20002, B2 => 
                           n25194, ZN => n13902);
   U525 : OAI22_X1 port map( A1 => n18359, A2 => n25229, B1 => n20001, B2 => 
                           n25194, ZN => n13903);
   U526 : OAI22_X1 port map( A1 => n18325, A2 => n25224, B1 => n20000, B2 => 
                           n25190, ZN => n13904);
   U527 : OAI22_X1 port map( A1 => n18359, A2 => n25226, B1 => n19999, B2 => 
                           n25194, ZN => n13905);
   U528 : OAI22_X1 port map( A1 => n18328, A2 => n25228, B1 => n19998, B2 => 
                           n25187, ZN => n13906);
   U529 : OAI22_X1 port map( A1 => n18328, A2 => n25223, B1 => n19997, B2 => 
                           n25187, ZN => n13907);
   U530 : OAI22_X1 port map( A1 => n18325, A2 => n25223, B1 => n19996, B2 => 
                           n25190, ZN => n13908);
   U531 : OAI22_X1 port map( A1 => n18325, A2 => n25229, B1 => n19995, B2 => 
                           n25190, ZN => n13909);
   U532 : OAI22_X1 port map( A1 => n18327, A2 => n25223, B1 => n19994, B2 => 
                           n25191, ZN => n13910);
   U533 : OAI22_X1 port map( A1 => n18328, A2 => n25230, B1 => n19993, B2 => 
                           n25187, ZN => n13911);
   U534 : OAI22_X1 port map( A1 => n18328, A2 => n25226, B1 => n19992, B2 => 
                           n25187, ZN => n13913);
   U535 : OAI22_X1 port map( A1 => n18326, A2 => n25228, B1 => n19991, B2 => 
                           n25189, ZN => n13914);
   U536 : OAI22_X1 port map( A1 => n18325, A2 => n25222, B1 => n19990, B2 => 
                           n25190, ZN => n13915);
   U537 : OAI22_X1 port map( A1 => n18326, A2 => n25222, B1 => n19989, B2 => 
                           n25189, ZN => n13917);
   U538 : OAI22_X1 port map( A1 => n18327, A2 => n25222, B1 => n19988, B2 => 
                           n25191, ZN => n13919);
   U539 : OAI22_X1 port map( A1 => n18325, A2 => n25226, B1 => n19987, B2 => 
                           n25190, ZN => n13920);
   U540 : OAI22_X1 port map( A1 => n18325, A2 => n25228, B1 => n19986, B2 => 
                           n25190, ZN => n13922);
   U541 : OAI22_X1 port map( A1 => n18345, A2 => n25228, B1 => n19985, B2 => 
                           n25245, ZN => n13923);
   U542 : OAI22_X1 port map( A1 => n18345, A2 => n25230, B1 => n19984, B2 => 
                           n25245, ZN => n13924);
   U543 : OAI22_X1 port map( A1 => n18345, A2 => n25197, B1 => n19983, B2 => 
                           n25245, ZN => n13925);
   U544 : OAI22_X1 port map( A1 => n18345, A2 => n25205, B1 => n19982, B2 => 
                           n25245, ZN => n13926);
   U545 : OAI22_X1 port map( A1 => n18345, A2 => n25226, B1 => n19981, B2 => 
                           n25245, ZN => n13927);
   U546 : OAI22_X1 port map( A1 => n18345, A2 => n25200, B1 => n19980, B2 => 
                           n25245, ZN => n13928);
   U547 : OAI22_X1 port map( A1 => n18345, A2 => n25201, B1 => n19979, B2 => 
                           n25245, ZN => n13929);
   U548 : OAI22_X1 port map( A1 => n18345, A2 => n25207, B1 => n19978, B2 => 
                           n25245, ZN => n13930);
   U549 : OAI22_X1 port map( A1 => n18345, A2 => n25216, B1 => n19977, B2 => 
                           n25245, ZN => n13931);
   U550 : OAI22_X1 port map( A1 => n18345, A2 => n25224, B1 => n19976, B2 => 
                           n25245, ZN => n13932);
   U551 : OAI22_X1 port map( A1 => n18345, A2 => n25210, B1 => n19975, B2 => 
                           n25245, ZN => n13933);
   U552 : OAI22_X1 port map( A1 => n18345, A2 => n25203, B1 => n19974, B2 => 
                           n25245, ZN => n13934);
   U553 : OAI22_X1 port map( A1 => n18345, A2 => n25211, B1 => n19973, B2 => 
                           n25245, ZN => n13935);
   U554 : OAI22_X1 port map( A1 => n18345, A2 => n25199, B1 => n19972, B2 => 
                           n25245, ZN => n13936);
   U555 : OAI22_X1 port map( A1 => n18345, A2 => n25196, B1 => n19971, B2 => 
                           n25245, ZN => n13937);
   U556 : OAI22_X1 port map( A1 => n18345, A2 => n25229, B1 => n19970, B2 => 
                           n25245, ZN => n13938);
   U557 : OAI22_X1 port map( A1 => n18345, A2 => n25195, B1 => n19969, B2 => 
                           n25245, ZN => n13939);
   U558 : OAI22_X1 port map( A1 => n18345, A2 => n25223, B1 => n19968, B2 => 
                           n25245, ZN => n13940);
   U559 : OAI22_X1 port map( A1 => n18345, A2 => n25202, B1 => n19967, B2 => 
                           n25245, ZN => n13941);
   U560 : OAI22_X1 port map( A1 => n18345, A2 => n25206, B1 => n19966, B2 => 
                           n25245, ZN => n13942);
   U561 : OAI22_X1 port map( A1 => n18345, A2 => n25198, B1 => n19965, B2 => 
                           n25245, ZN => n13943);
   U562 : OAI22_X1 port map( A1 => n18336, A2 => n25198, B1 => n19964, B2 => 
                           n25231, ZN => n13944);
   U563 : OAI22_X1 port map( A1 => n18335, A2 => n25222, B1 => n19963, B2 => 
                           n25239, ZN => n13945);
   U564 : OAI22_X1 port map( A1 => n18336, A2 => n25222, B1 => n19962, B2 => 
                           n25231, ZN => n13946);
   U565 : OAI22_X1 port map( A1 => n18337, A2 => n25198, B1 => n19961, B2 => 
                           n25235, ZN => n13947);
   U566 : OAI22_X1 port map( A1 => n18335, A2 => n25197, B1 => n19960, B2 => 
                           n25239, ZN => n13948);
   U567 : OAI22_X1 port map( A1 => n18336, A2 => n25197, B1 => n19959, B2 => 
                           n25231, ZN => n13949);
   U568 : OAI22_X1 port map( A1 => n18337, A2 => n25197, B1 => n19958, B2 => 
                           n25235, ZN => n13950);
   U569 : OAI22_X1 port map( A1 => n18337, A2 => n25222, B1 => n19957, B2 => 
                           n25235, ZN => n13951);
   U570 : OAI22_X1 port map( A1 => n18335, A2 => n25223, B1 => n19956, B2 => 
                           n25239, ZN => n13952);
   U571 : OAI22_X1 port map( A1 => n18336, A2 => n25223, B1 => n19955, B2 => 
                           n25231, ZN => n13953);
   U572 : OAI22_X1 port map( A1 => n18337, A2 => n25223, B1 => n19954, B2 => 
                           n25235, ZN => n13954);
   U573 : OAI22_X1 port map( A1 => n18336, A2 => n25224, B1 => n19953, B2 => 
                           n25231, ZN => n13955);
   U574 : OAI22_X1 port map( A1 => n18337, A2 => n25224, B1 => n19952, B2 => 
                           n25235, ZN => n13956);
   U575 : OAI22_X1 port map( A1 => n18335, A2 => n25224, B1 => n19951, B2 => 
                           n25239, ZN => n13957);
   U576 : OAI22_X1 port map( A1 => n18336, A2 => n25196, B1 => n19950, B2 => 
                           n25231, ZN => n13958);
   U577 : OAI22_X1 port map( A1 => n18337, A2 => n25196, B1 => n19949, B2 => 
                           n25235, ZN => n13959);
   U578 : OAI22_X1 port map( A1 => n18335, A2 => n25196, B1 => n19948, B2 => 
                           n25239, ZN => n13960);
   U579 : OAI22_X1 port map( A1 => n18331, A2 => n25198, B1 => n19947, B2 => 
                           n25242, ZN => n13961);
   U580 : OAI22_X1 port map( A1 => n18331, A2 => n25196, B1 => n19946, B2 => 
                           n25242, ZN => n13962);
   U581 : OAI22_X1 port map( A1 => n18331, A2 => n25197, B1 => n19945, B2 => 
                           n25242, ZN => n13963);
   U582 : OAI22_X1 port map( A1 => n18331, A2 => n25222, B1 => n19944, B2 => 
                           n25242, ZN => n13964);
   U583 : OAI22_X1 port map( A1 => n18331, A2 => n25224, B1 => n19943, B2 => 
                           n25242, ZN => n13965);
   U584 : OAI22_X1 port map( A1 => n18331, A2 => n25223, B1 => n19942, B2 => 
                           n25242, ZN => n13966);
   U585 : OAI22_X1 port map( A1 => n18336, A2 => n25210, B1 => n19941, B2 => 
                           n25231, ZN => n13967);
   U586 : OAI22_X1 port map( A1 => n18332, A2 => n25198, B1 => n19940, B2 => 
                           n25243, ZN => n13968);
   U587 : OAI22_X1 port map( A1 => n18332, A2 => n25196, B1 => n19939, B2 => 
                           n25243, ZN => n13969);
   U588 : OAI22_X1 port map( A1 => n18332, A2 => n25197, B1 => n19938, B2 => 
                           n25243, ZN => n13970);
   U589 : OAI22_X1 port map( A1 => n18332, A2 => n25222, B1 => n19937, B2 => 
                           n25243, ZN => n13971);
   U590 : OAI22_X1 port map( A1 => n18332, A2 => n25224, B1 => n19936, B2 => 
                           n25243, ZN => n13972);
   U591 : OAI22_X1 port map( A1 => n18332, A2 => n25223, B1 => n19935, B2 => 
                           n25243, ZN => n13973);
   U592 : OAI22_X1 port map( A1 => n18336, A2 => n25195, B1 => n19934, B2 => 
                           n25231, ZN => n13974);
   U593 : OAI22_X1 port map( A1 => n18337, A2 => n25195, B1 => n19933, B2 => 
                           n25235, ZN => n13975);
   U594 : OAI22_X1 port map( A1 => n18338, A2 => n25195, B1 => n19932, B2 => 
                           n25214, ZN => n13976);
   U595 : OAI22_X1 port map( A1 => n18333, A2 => n25198, B1 => n19931, B2 => 
                           n25213, ZN => n13977);
   U596 : OAI22_X1 port map( A1 => n18331, A2 => n25195, B1 => n19930, B2 => 
                           n25242, ZN => n13978);
   U597 : OAI22_X1 port map( A1 => n18332, A2 => n25195, B1 => n19929, B2 => 
                           n25243, ZN => n13979);
   U598 : OAI22_X1 port map( A1 => n18333, A2 => n25195, B1 => n19928, B2 => 
                           n25213, ZN => n13980);
   U599 : OAI22_X1 port map( A1 => n18333, A2 => n25196, B1 => n19927, B2 => 
                           n25213, ZN => n13981);
   U600 : OAI22_X1 port map( A1 => n18333, A2 => n25197, B1 => n19926, B2 => 
                           n25213, ZN => n13982);
   U601 : OAI22_X1 port map( A1 => n18333, A2 => n25222, B1 => n19925, B2 => 
                           n25213, ZN => n13983);
   U602 : OAI22_X1 port map( A1 => n18333, A2 => n25224, B1 => n19924, B2 => 
                           n25213, ZN => n13984);
   U603 : OAI22_X1 port map( A1 => n18333, A2 => n25223, B1 => n19923, B2 => 
                           n25213, ZN => n13985);
   U604 : OAI22_X1 port map( A1 => n18337, A2 => n25202, B1 => n19922, B2 => 
                           n25235, ZN => n13986);
   U605 : OAI22_X1 port map( A1 => n18338, A2 => n25202, B1 => n19921, B2 => 
                           n25214, ZN => n13987);
   U606 : OAI22_X1 port map( A1 => n18332, A2 => n25202, B1 => n19920, B2 => 
                           n25243, ZN => n13988);
   U607 : OAI22_X1 port map( A1 => n18333, A2 => n25202, B1 => n19919, B2 => 
                           n25213, ZN => n13989);
   U608 : OAI22_X1 port map( A1 => n18336, A2 => n25202, B1 => n19918, B2 => 
                           n25231, ZN => n13990);
   U609 : OAI22_X1 port map( A1 => n18338, A2 => n25216, B1 => n19917, B2 => 
                           n25214, ZN => n13991);
   U610 : OAI22_X1 port map( A1 => n18337, A2 => n25204, B1 => n19916, B2 => 
                           n25235, ZN => n13992);
   U611 : OAI22_X1 port map( A1 => n18336, A2 => n25204, B1 => n19915, B2 => 
                           n25231, ZN => n13993);
   U612 : OAI22_X1 port map( A1 => n18333, A2 => n25204, B1 => n19914, B2 => 
                           n25213, ZN => n13994);
   U613 : OAI22_X1 port map( A1 => n18332, A2 => n25204, B1 => n19913, B2 => 
                           n25243, ZN => n13995);
   U614 : OAI22_X1 port map( A1 => n18331, A2 => n25204, B1 => n19912, B2 => 
                           n25242, ZN => n13996);
   U615 : OAI22_X1 port map( A1 => n18335, A2 => n25204, B1 => n19911, B2 => 
                           n25239, ZN => n13997);
   U616 : OAI22_X1 port map( A1 => n18335, A2 => n25198, B1 => n19910, B2 => 
                           n25239, ZN => n13998);
   U617 : OAI22_X1 port map( A1 => n18335, A2 => n25202, B1 => n19909, B2 => 
                           n25239, ZN => n13999);
   U618 : OAI22_X1 port map( A1 => n18335, A2 => n25195, B1 => n19908, B2 => 
                           n25239, ZN => n14000);
   U619 : OAI22_X1 port map( A1 => n18337, A2 => n25199, B1 => n19907, B2 => 
                           n25235, ZN => n14001);
   U620 : OAI22_X1 port map( A1 => n18336, A2 => n25199, B1 => n19906, B2 => 
                           n25231, ZN => n14002);
   U621 : OAI22_X1 port map( A1 => n18335, A2 => n25199, B1 => n19905, B2 => 
                           n25239, ZN => n14003);
   U622 : OAI22_X1 port map( A1 => n18333, A2 => n25199, B1 => n19904, B2 => 
                           n25213, ZN => n14004);
   U623 : OAI22_X1 port map( A1 => n18332, A2 => n25199, B1 => n19903, B2 => 
                           n25243, ZN => n14005);
   U624 : OAI22_X1 port map( A1 => n18331, A2 => n25199, B1 => n19902, B2 => 
                           n25242, ZN => n14006);
   U625 : OAI22_X1 port map( A1 => n18334, A2 => n25223, B1 => n19901, B2 => 
                           n25244, ZN => n14007);
   U626 : OAI22_X1 port map( A1 => n18337, A2 => n25200, B1 => n19900, B2 => 
                           n25235, ZN => n14008);
   U627 : OAI22_X1 port map( A1 => n18336, A2 => n25200, B1 => n19899, B2 => 
                           n25231, ZN => n14009);
   U628 : OAI22_X1 port map( A1 => n18335, A2 => n25200, B1 => n19898, B2 => 
                           n25239, ZN => n14010);
   U629 : OAI22_X1 port map( A1 => n18333, A2 => n25200, B1 => n19897, B2 => 
                           n25213, ZN => n14011);
   U630 : OAI22_X1 port map( A1 => n18332, A2 => n25200, B1 => n19896, B2 => 
                           n25243, ZN => n14012);
   U631 : OAI22_X1 port map( A1 => n18331, A2 => n25200, B1 => n19895, B2 => 
                           n25242, ZN => n14013);
   U632 : OAI22_X1 port map( A1 => n18334, A2 => n25224, B1 => n19894, B2 => 
                           n25244, ZN => n14014);
   U633 : OAI22_X1 port map( A1 => n18334, A2 => n25222, B1 => n19893, B2 => 
                           n25244, ZN => n14015);
   U634 : OAI22_X1 port map( A1 => n18334, A2 => n25197, B1 => n19892, B2 => 
                           n25244, ZN => n14016);
   U635 : OAI22_X1 port map( A1 => n18334, A2 => n25196, B1 => n19891, B2 => 
                           n25244, ZN => n14017);
   U636 : OAI22_X1 port map( A1 => n18334, A2 => n25204, B1 => n19890, B2 => 
                           n25244, ZN => n14018);
   U637 : OAI22_X1 port map( A1 => n18334, A2 => n25198, B1 => n19889, B2 => 
                           n25244, ZN => n14019);
   U638 : OAI22_X1 port map( A1 => n18334, A2 => n25199, B1 => n19888, B2 => 
                           n25244, ZN => n14020);
   U639 : OAI22_X1 port map( A1 => n18334, A2 => n25200, B1 => n19887, B2 => 
                           n25244, ZN => n14021);
   U640 : OAI22_X1 port map( A1 => n18337, A2 => n25201, B1 => n19886, B2 => 
                           n25235, ZN => n14022);
   U641 : OAI22_X1 port map( A1 => n18336, A2 => n25201, B1 => n19885, B2 => 
                           n25231, ZN => n14023);
   U642 : OAI22_X1 port map( A1 => n18335, A2 => n25201, B1 => n19884, B2 => 
                           n25239, ZN => n14024);
   U643 : OAI22_X1 port map( A1 => n18334, A2 => n25201, B1 => n19883, B2 => 
                           n25244, ZN => n14025);
   U644 : OAI22_X1 port map( A1 => n18333, A2 => n25201, B1 => n19882, B2 => 
                           n25213, ZN => n14026);
   U645 : OAI22_X1 port map( A1 => n18332, A2 => n25201, B1 => n19881, B2 => 
                           n25243, ZN => n14027);
   U646 : CLKBUF_X1 port map( A => n25201, Z => n25208);
   U647 : OAI22_X1 port map( A1 => n18331, A2 => n25208, B1 => n19880, B2 => 
                           n25242, ZN => n14028);
   U648 : OAI22_X1 port map( A1 => n18334, A2 => n25202, B1 => n19879, B2 => 
                           n25244, ZN => n14029);
   U649 : OAI22_X1 port map( A1 => n18334, A2 => n25195, B1 => n19878, B2 => 
                           n25244, ZN => n14030);
   U650 : OAI22_X1 port map( A1 => n18337, A2 => n25216, B1 => n19877, B2 => 
                           n25235, ZN => n14031);
   U651 : OAI22_X1 port map( A1 => n18335, A2 => n25216, B1 => n19876, B2 => 
                           n25239, ZN => n14032);
   U652 : OAI22_X1 port map( A1 => n18334, A2 => n25216, B1 => n19875, B2 => 
                           n25244, ZN => n14033);
   U653 : OAI22_X1 port map( A1 => n18333, A2 => n25216, B1 => n19874, B2 => 
                           n25213, ZN => n14034);
   U654 : OAI22_X1 port map( A1 => n18332, A2 => n25216, B1 => n19873, B2 => 
                           n25243, ZN => n14035);
   U655 : OAI22_X1 port map( A1 => n18331, A2 => n25216, B1 => n19872, B2 => 
                           n25242, ZN => n14036);
   U656 : OAI22_X1 port map( A1 => n18331, A2 => n25202, B1 => n19871, B2 => 
                           n25242, ZN => n14037);
   U657 : OAI22_X1 port map( A1 => n18331, A2 => n25226, B1 => n19870, B2 => 
                           n25242, ZN => n14038);
   U658 : OAI22_X1 port map( A1 => n18333, A2 => n25226, B1 => n19869, B2 => 
                           n25213, ZN => n14039);
   U659 : OAI22_X1 port map( A1 => n18334, A2 => n25226, B1 => n19868, B2 => 
                           n25244, ZN => n14040);
   U660 : OAI22_X1 port map( A1 => n18335, A2 => n25226, B1 => n19867, B2 => 
                           n25239, ZN => n14041);
   U661 : OAI22_X1 port map( A1 => n18340, A2 => n25195, B1 => n19866, B2 => 
                           n25240, ZN => n14042);
   U662 : OAI22_X1 port map( A1 => n18340, A2 => n25202, B1 => n19865, B2 => 
                           n25240, ZN => n14043);
   U663 : OAI22_X1 port map( A1 => n18340, A2 => n25216, B1 => n19864, B2 => 
                           n25240, ZN => n14044);
   U664 : OAI22_X1 port map( A1 => n18340, A2 => n25208, B1 => n19863, B2 => 
                           n25240, ZN => n14045);
   U665 : OAI22_X1 port map( A1 => n18340, A2 => n25200, B1 => n19862, B2 => 
                           n25240, ZN => n14046);
   U666 : OAI22_X1 port map( A1 => n18340, A2 => n25199, B1 => n19861, B2 => 
                           n25240, ZN => n14047);
   U667 : OAI22_X1 port map( A1 => n18340, A2 => n25198, B1 => n19860, B2 => 
                           n25240, ZN => n14048);
   U668 : OAI22_X1 port map( A1 => n18344, A2 => n25203, B1 => n19859, B2 => 
                           n25238, ZN => n14049);
   U669 : OAI22_X1 port map( A1 => n18340, A2 => n25204, B1 => n19858, B2 => 
                           n25240, ZN => n14050);
   U670 : OAI22_X1 port map( A1 => n18340, A2 => n25196, B1 => n19857, B2 => 
                           n25240, ZN => n14051);
   U671 : OAI22_X1 port map( A1 => n18331, A2 => n25203, B1 => n19856, B2 => 
                           n25242, ZN => n14052);
   U672 : OAI22_X1 port map( A1 => n18332, A2 => n25203, B1 => n19855, B2 => 
                           n25243, ZN => n14053);
   U673 : OAI22_X1 port map( A1 => n18333, A2 => n25203, B1 => n19854, B2 => 
                           n25213, ZN => n14054);
   U674 : OAI22_X1 port map( A1 => n18334, A2 => n25203, B1 => n19853, B2 => 
                           n25244, ZN => n14055);
   U675 : OAI22_X1 port map( A1 => n18335, A2 => n25203, B1 => n19852, B2 => 
                           n25239, ZN => n14056);
   U676 : OAI22_X1 port map( A1 => n18336, A2 => n25203, B1 => n19851, B2 => 
                           n25231, ZN => n14057);
   U677 : OAI22_X1 port map( A1 => n18337, A2 => n25203, B1 => n19850, B2 => 
                           n25235, ZN => n14058);
   U678 : OAI22_X1 port map( A1 => n18344, A2 => n25223, B1 => n19849, B2 => 
                           n25238, ZN => n14059);
   U679 : OAI22_X1 port map( A1 => n18339, A2 => n25203, B1 => n19848, B2 => 
                           n25225, ZN => n14060);
   U680 : OAI22_X1 port map( A1 => n18340, A2 => n25197, B1 => n19847, B2 => 
                           n25240, ZN => n14061);
   U681 : OAI22_X1 port map( A1 => n18340, A2 => n25222, B1 => n19846, B2 => 
                           n25240, ZN => n14062);
   U682 : OAI22_X1 port map( A1 => n18340, A2 => n25224, B1 => n19845, B2 => 
                           n25240, ZN => n14063);
   U683 : OAI22_X1 port map( A1 => n18340, A2 => n25223, B1 => n19844, B2 => 
                           n25240, ZN => n14064);
   U684 : OAI22_X1 port map( A1 => n18344, A2 => n25224, B1 => n19843, B2 => 
                           n25238, ZN => n14065);
   U685 : OAI22_X1 port map( A1 => n18344, A2 => n25222, B1 => n19842, B2 => 
                           n25238, ZN => n14066);
   U686 : OAI22_X1 port map( A1 => n18344, A2 => n25197, B1 => n19841, B2 => 
                           n25238, ZN => n14067);
   U687 : OAI22_X1 port map( A1 => n18340, A2 => n25203, B1 => n19840, B2 => 
                           n25240, ZN => n14068);
   U688 : OAI22_X1 port map( A1 => n18344, A2 => n25196, B1 => n19839, B2 => 
                           n25238, ZN => n14069);
   U689 : OAI22_X1 port map( A1 => n18344, A2 => n25204, B1 => n19838, B2 => 
                           n25238, ZN => n14070);
   U690 : OAI22_X1 port map( A1 => n18334, A2 => n25229, B1 => n19837, B2 => 
                           n25244, ZN => n14071);
   U691 : OAI22_X1 port map( A1 => n18335, A2 => n25229, B1 => n19836, B2 => 
                           n25239, ZN => n14072);
   U692 : OAI22_X1 port map( A1 => n18344, A2 => n25198, B1 => n19835, B2 => 
                           n25238, ZN => n14073);
   U693 : OAI22_X1 port map( A1 => n18344, A2 => n25199, B1 => n19834, B2 => 
                           n25238, ZN => n14074);
   U694 : OAI22_X1 port map( A1 => n18344, A2 => n25200, B1 => n19833, B2 => 
                           n25238, ZN => n14075);
   U695 : OAI22_X1 port map( A1 => n18344, A2 => n25208, B1 => n19832, B2 => 
                           n25238, ZN => n14076);
   U696 : OAI22_X1 port map( A1 => n18337, A2 => n25229, B1 => n19831, B2 => 
                           n25235, ZN => n14077);
   U697 : OAI22_X1 port map( A1 => n18339, A2 => n25229, B1 => n19830, B2 => 
                           n25225, ZN => n14078);
   U698 : OAI22_X1 port map( A1 => n18344, A2 => n25216, B1 => n19829, B2 => 
                           n25238, ZN => n14079);
   U699 : OAI22_X1 port map( A1 => n18344, A2 => n25229, B1 => n19828, B2 => 
                           n25238, ZN => n14080);
   U700 : OAI22_X1 port map( A1 => n18344, A2 => n25202, B1 => n19827, B2 => 
                           n25238, ZN => n14081);
   U701 : OAI22_X1 port map( A1 => n18331, A2 => n25229, B1 => n19826, B2 => 
                           n25242, ZN => n14082);
   U702 : OAI22_X1 port map( A1 => n18344, A2 => n25195, B1 => n19825, B2 => 
                           n25238, ZN => n14083);
   U703 : OAI22_X1 port map( A1 => n18333, A2 => n25229, B1 => n19824, B2 => 
                           n25213, ZN => n14084);
   U704 : OAI22_X1 port map( A1 => n18335, A2 => n25230, B1 => n19823, B2 => 
                           n25239, ZN => n14085);
   U705 : OAI22_X1 port map( A1 => n18337, A2 => n25230, B1 => n19822, B2 => 
                           n25235, ZN => n14086);
   U706 : OAI22_X1 port map( A1 => n18339, A2 => n25230, B1 => n19821, B2 => 
                           n25225, ZN => n14087);
   U707 : OAI22_X1 port map( A1 => n18340, A2 => n25230, B1 => n19820, B2 => 
                           n25240, ZN => n14088);
   U708 : OAI22_X1 port map( A1 => n18344, A2 => n25230, B1 => n19819, B2 => 
                           n25238, ZN => n14089);
   U709 : OAI22_X1 port map( A1 => n18331, A2 => n25230, B1 => n19818, B2 => 
                           n25242, ZN => n14090);
   U710 : OAI22_X1 port map( A1 => n18333, A2 => n25230, B1 => n19817, B2 => 
                           n25213, ZN => n14091);
   U711 : OAI22_X1 port map( A1 => n18334, A2 => n25230, B1 => n19816, B2 => 
                           n25244, ZN => n14092);
   U712 : OAI22_X1 port map( A1 => n18343, A2 => n25203, B1 => n19815, B2 => 
                           n25236, ZN => n14094);
   U713 : OAI22_X1 port map( A1 => n18344, A2 => n25228, B1 => n19814, B2 => 
                           n25238, ZN => n14095);
   U714 : OAI22_X1 port map( A1 => n18333, A2 => n25228, B1 => n19813, B2 => 
                           n25213, ZN => n14096);
   U715 : OAI22_X1 port map( A1 => n18344, A2 => n25226, B1 => n19812, B2 => 
                           n25238, ZN => n14097);
   U716 : OAI22_X1 port map( A1 => n18334, A2 => n25228, B1 => n19811, B2 => 
                           n25244, ZN => n14098);
   U717 : OAI22_X1 port map( A1 => n18335, A2 => n25228, B1 => n19810, B2 => 
                           n25239, ZN => n14099);
   U718 : OAI22_X1 port map( A1 => n18337, A2 => n25228, B1 => n19809, B2 => 
                           n25235, ZN => n14100);
   U719 : OAI22_X1 port map( A1 => n18339, A2 => n25228, B1 => n19808, B2 => 
                           n25225, ZN => n14101);
   U720 : OAI22_X1 port map( A1 => n18340, A2 => n25229, B1 => n19807, B2 => 
                           n25240, ZN => n14102);
   U721 : OAI22_X1 port map( A1 => n18331, A2 => n25228, B1 => n19806, B2 => 
                           n25242, ZN => n14103);
   U722 : OAI22_X1 port map( A1 => n18340, A2 => n25228, B1 => n19805, B2 => 
                           n25240, ZN => n14104);
   U723 : OAI22_X1 port map( A1 => n18343, A2 => n25197, B1 => n19804, B2 => 
                           n25236, ZN => n14105);
   U724 : OAI22_X1 port map( A1 => n18343, A2 => n25196, B1 => n19803, B2 => 
                           n25236, ZN => n14106);
   U725 : OAI22_X1 port map( A1 => n18343, A2 => n25204, B1 => n19802, B2 => 
                           n25236, ZN => n14107);
   U726 : OAI22_X1 port map( A1 => n18333, A2 => n25205, B1 => n19801, B2 => 
                           n25213, ZN => n14108);
   U727 : OAI22_X1 port map( A1 => n18334, A2 => n25205, B1 => n19800, B2 => 
                           n25244, ZN => n14109);
   U728 : OAI22_X1 port map( A1 => n18335, A2 => n25205, B1 => n19799, B2 => 
                           n25239, ZN => n14110);
   U729 : OAI22_X1 port map( A1 => n18336, A2 => n25205, B1 => n19798, B2 => 
                           n25231, ZN => n14111);
   U730 : OAI22_X1 port map( A1 => n18337, A2 => n25205, B1 => n19797, B2 => 
                           n25235, ZN => n14112);
   U731 : OAI22_X1 port map( A1 => n18339, A2 => n25205, B1 => n19796, B2 => 
                           n25225, ZN => n14113);
   U732 : OAI22_X1 port map( A1 => n18343, A2 => n25198, B1 => n19795, B2 => 
                           n25236, ZN => n14114);
   U733 : OAI22_X1 port map( A1 => n18340, A2 => n25212, B1 => n19794, B2 => 
                           n25240, ZN => n14115);
   U734 : OAI22_X1 port map( A1 => n18343, A2 => n25212, B1 => n19793, B2 => 
                           n25236, ZN => n14116);
   U735 : OAI22_X1 port map( A1 => n18343, A2 => n25199, B1 => n19792, B2 => 
                           n25236, ZN => n14117);
   U736 : OAI22_X1 port map( A1 => n18343, A2 => n25200, B1 => n19791, B2 => 
                           n25236, ZN => n14118);
   U737 : OAI22_X1 port map( A1 => n18341, A2 => n25195, B1 => n19790, B2 => 
                           n25227, ZN => n14119);
   U738 : OAI22_X1 port map( A1 => n18341, A2 => n25202, B1 => n19789, B2 => 
                           n25227, ZN => n14120);
   U739 : OAI22_X1 port map( A1 => n18331, A2 => n25212, B1 => n19788, B2 => 
                           n25242, ZN => n14121);
   U740 : OAI22_X1 port map( A1 => n18332, A2 => n25212, B1 => n19787, B2 => 
                           n25243, ZN => n14123);
   U741 : OAI22_X1 port map( A1 => n18343, A2 => n25208, B1 => n19786, B2 => 
                           n25236, ZN => n14124);
   U742 : OAI22_X1 port map( A1 => n18343, A2 => n25202, B1 => n19785, B2 => 
                           n25236, ZN => n14126);
   U743 : OAI22_X1 port map( A1 => n18343, A2 => n25195, B1 => n19784, B2 => 
                           n25236, ZN => n14128);
   U744 : OAI22_X1 port map( A1 => n18341, A2 => n25208, B1 => n19783, B2 => 
                           n25227, ZN => n14130);
   U745 : OAI22_X1 port map( A1 => n18341, A2 => n25200, B1 => n19782, B2 => 
                           n25227, ZN => n14132);
   U746 : OAI22_X1 port map( A1 => n18341, A2 => n25199, B1 => n19781, B2 => 
                           n25227, ZN => n14133);
   U747 : OAI22_X1 port map( A1 => n18342, A2 => n25228, B1 => n19780, B2 => 
                           n25241, ZN => n14134);
   U748 : OAI22_X1 port map( A1 => n18342, A2 => n25212, B1 => n19779, B2 => 
                           n25241, ZN => n14135);
   U749 : OAI22_X1 port map( A1 => n18342, A2 => n25229, B1 => n19778, B2 => 
                           n25241, ZN => n14136);
   U750 : OAI22_X1 port map( A1 => n18342, A2 => n25230, B1 => n19777, B2 => 
                           n25241, ZN => n14137);
   U751 : OAI22_X1 port map( A1 => n18342, A2 => n25203, B1 => n19776, B2 => 
                           n25241, ZN => n14138);
   U752 : OAI22_X1 port map( A1 => n18341, A2 => n25198, B1 => n19775, B2 => 
                           n25227, ZN => n14139);
   U753 : OAI22_X1 port map( A1 => n18341, A2 => n25204, B1 => n19774, B2 => 
                           n25227, ZN => n14140);
   U754 : OAI22_X1 port map( A1 => n18341, A2 => n25196, B1 => n19773, B2 => 
                           n25227, ZN => n14141);
   U755 : OAI22_X1 port map( A1 => n18341, A2 => n25197, B1 => n19772, B2 => 
                           n25227, ZN => n14142);
   U756 : OAI22_X1 port map( A1 => n18341, A2 => n25222, B1 => n19771, B2 => 
                           n25227, ZN => n14143);
   U757 : OAI22_X1 port map( A1 => n18341, A2 => n25224, B1 => n19770, B2 => 
                           n25227, ZN => n14144);
   U758 : OAI22_X1 port map( A1 => n18342, A2 => n25206, B1 => n19769, B2 => 
                           n25241, ZN => n14145);
   U759 : OAI22_X1 port map( A1 => n18343, A2 => n25206, B1 => n19768, B2 => 
                           n25236, ZN => n14146);
   U760 : OAI22_X1 port map( A1 => n18344, A2 => n25206, B1 => n19767, B2 => 
                           n25238, ZN => n14147);
   U761 : OAI22_X1 port map( A1 => n18341, A2 => n25223, B1 => n19766, B2 => 
                           n25227, ZN => n14148);
   U762 : OAI22_X1 port map( A1 => n18341, A2 => n25203, B1 => n19765, B2 => 
                           n25227, ZN => n14149);
   U763 : OAI22_X1 port map( A1 => n18331, A2 => n25206, B1 => n19764, B2 => 
                           n25242, ZN => n14150);
   U764 : OAI22_X1 port map( A1 => n18332, A2 => n25206, B1 => n19763, B2 => 
                           n25243, ZN => n14151);
   U765 : OAI22_X1 port map( A1 => n18333, A2 => n25206, B1 => n19762, B2 => 
                           n25213, ZN => n14152);
   U766 : OAI22_X1 port map( A1 => n18334, A2 => n25206, B1 => n19761, B2 => 
                           n25244, ZN => n14153);
   U767 : OAI22_X1 port map( A1 => n18335, A2 => n25206, B1 => n19760, B2 => 
                           n25239, ZN => n14154);
   U768 : OAI22_X1 port map( A1 => n18336, A2 => n25206, B1 => n19759, B2 => 
                           n25231, ZN => n14155);
   U769 : OAI22_X1 port map( A1 => n18337, A2 => n25206, B1 => n19758, B2 => 
                           n25235, ZN => n14156);
   U770 : OAI22_X1 port map( A1 => n18339, A2 => n25206, B1 => n19757, B2 => 
                           n25225, ZN => n14157);
   U771 : OAI22_X1 port map( A1 => n18340, A2 => n25206, B1 => n19756, B2 => 
                           n25240, ZN => n14158);
   U772 : OAI22_X1 port map( A1 => n18341, A2 => n25230, B1 => n19755, B2 => 
                           n25227, ZN => n14159);
   U773 : OAI22_X1 port map( A1 => n18341, A2 => n25229, B1 => n19754, B2 => 
                           n25227, ZN => n14160);
   U774 : OAI22_X1 port map( A1 => n18341, A2 => n25212, B1 => n19753, B2 => 
                           n25227, ZN => n14161);
   U775 : OAI22_X1 port map( A1 => n18341, A2 => n25228, B1 => n19752, B2 => 
                           n25227, ZN => n14162);
   U776 : OAI22_X1 port map( A1 => n18341, A2 => n25206, B1 => n19751, B2 => 
                           n25227, ZN => n14164);
   U777 : OAI22_X1 port map( A1 => n18342, A2 => n25197, B1 => n19750, B2 => 
                           n25241, ZN => n14166);
   U778 : OAI22_X1 port map( A1 => n18342, A2 => n25196, B1 => n19749, B2 => 
                           n25241, ZN => n14168);
   U779 : OAI22_X1 port map( A1 => n18342, A2 => n25204, B1 => n19748, B2 => 
                           n25241, ZN => n14170);
   U780 : OAI22_X1 port map( A1 => n18342, A2 => n25198, B1 => n19747, B2 => 
                           n25241, ZN => n14172);
   U781 : OAI22_X1 port map( A1 => n18342, A2 => n25199, B1 => n19746, B2 => 
                           n25241, ZN => n14174);
   U782 : OAI22_X1 port map( A1 => n18342, A2 => n25200, B1 => n19745, B2 => 
                           n25241, ZN => n14175);
   U783 : OAI22_X1 port map( A1 => n18342, A2 => n25208, B1 => n19744, B2 => 
                           n25241, ZN => n14176);
   U784 : OAI22_X1 port map( A1 => n18342, A2 => n25195, B1 => n19743, B2 => 
                           n25241, ZN => n14177);
   U785 : OAI22_X1 port map( A1 => n18342, A2 => n25202, B1 => n19742, B2 => 
                           n25241, ZN => n14178);
   U786 : OAI22_X1 port map( A1 => n18342, A2 => n25216, B1 => n19741, B2 => 
                           n25241, ZN => n14179);
   U787 : OAI22_X1 port map( A1 => n18339, A2 => n25226, B1 => n19740, B2 => 
                           n25225, ZN => n14180);
   U788 : OAI22_X1 port map( A1 => n18340, A2 => n25226, B1 => n19739, B2 => 
                           n25240, ZN => n14181);
   U789 : OAI22_X1 port map( A1 => n18337, A2 => n25226, B1 => n19738, B2 => 
                           n25235, ZN => n14182);
   U790 : OAI22_X1 port map( A1 => n18336, A2 => n25207, B1 => n19737, B2 => 
                           n25231, ZN => n14183);
   U791 : OAI22_X1 port map( A1 => n18335, A2 => n25207, B1 => n19736, B2 => 
                           n25239, ZN => n14184);
   U792 : OAI22_X1 port map( A1 => n18334, A2 => n25207, B1 => n19735, B2 => 
                           n25244, ZN => n14185);
   U793 : OAI22_X1 port map( A1 => n18333, A2 => n25207, B1 => n19734, B2 => 
                           n25213, ZN => n14186);
   U794 : OAI22_X1 port map( A1 => n18332, A2 => n25207, B1 => n19733, B2 => 
                           n25243, ZN => n14187);
   U795 : OAI22_X1 port map( A1 => n18331, A2 => n25207, B1 => n19732, B2 => 
                           n25242, ZN => n14188);
   U796 : OAI22_X1 port map( A1 => n18339, A2 => n25223, B1 => n19731, B2 => 
                           n25225, ZN => n14189);
   U797 : OAI22_X1 port map( A1 => n18339, A2 => n25224, B1 => n19730, B2 => 
                           n25225, ZN => n14190);
   U798 : OAI22_X1 port map( A1 => n18339, A2 => n25222, B1 => n19729, B2 => 
                           n25225, ZN => n14191);
   U799 : OAI22_X1 port map( A1 => n18339, A2 => n25197, B1 => n19728, B2 => 
                           n25225, ZN => n14192);
   U800 : OAI22_X1 port map( A1 => n18344, A2 => n25207, B1 => n19727, B2 => 
                           n25238, ZN => n14193);
   U801 : OAI22_X1 port map( A1 => n18343, A2 => n25207, B1 => n19726, B2 => 
                           n25236, ZN => n14194);
   U802 : OAI22_X1 port map( A1 => n18342, A2 => n25207, B1 => n19725, B2 => 
                           n25241, ZN => n14196);
   U803 : OAI22_X1 port map( A1 => n18341, A2 => n25207, B1 => n19724, B2 => 
                           n25227, ZN => n14197);
   U804 : OAI22_X1 port map( A1 => n18340, A2 => n25207, B1 => n19723, B2 => 
                           n25240, ZN => n14198);
   U805 : OAI22_X1 port map( A1 => n18339, A2 => n25207, B1 => n19722, B2 => 
                           n25225, ZN => n14199);
   U806 : OAI22_X1 port map( A1 => n18337, A2 => n25207, B1 => n19721, B2 => 
                           n25235, ZN => n14200);
   U807 : OAI22_X1 port map( A1 => n18339, A2 => n25196, B1 => n19720, B2 => 
                           n25225, ZN => n14201);
   U808 : OAI22_X1 port map( A1 => n18339, A2 => n25204, B1 => n19719, B2 => 
                           n25225, ZN => n14202);
   U809 : OAI22_X1 port map( A1 => n18339, A2 => n25198, B1 => n19718, B2 => 
                           n25225, ZN => n14203);
   U810 : OAI22_X1 port map( A1 => n18341, A2 => n25226, B1 => n19717, B2 => 
                           n25227, ZN => n14204);
   U811 : OAI22_X1 port map( A1 => n18339, A2 => n25199, B1 => n19716, B2 => 
                           n25225, ZN => n14205);
   U812 : OAI22_X1 port map( A1 => n18339, A2 => n25200, B1 => n19715, B2 => 
                           n25225, ZN => n14206);
   U813 : OAI22_X1 port map( A1 => n18339, A2 => n25208, B1 => n19714, B2 => 
                           n25225, ZN => n14207);
   U814 : OAI22_X1 port map( A1 => n18339, A2 => n25216, B1 => n19713, B2 => 
                           n25225, ZN => n14208);
   U815 : OAI22_X1 port map( A1 => n18337, A2 => n25209, B1 => n19712, B2 => 
                           n25235, ZN => n14209);
   U816 : OAI22_X1 port map( A1 => n18338, A2 => n25208, B1 => n19711, B2 => 
                           n25214, ZN => n14211);
   U817 : OAI22_X1 port map( A1 => n18336, A2 => n25209, B1 => n19710, B2 => 
                           n25231, ZN => n14212);
   U818 : OAI22_X1 port map( A1 => n18335, A2 => n25209, B1 => n19709, B2 => 
                           n25239, ZN => n14213);
   U819 : OAI22_X1 port map( A1 => n18334, A2 => n25209, B1 => n19708, B2 => 
                           n25244, ZN => n14214);
   U820 : OAI22_X1 port map( A1 => n18333, A2 => n25209, B1 => n19707, B2 => 
                           n25213, ZN => n14215);
   U821 : OAI22_X1 port map( A1 => n18332, A2 => n25209, B1 => n19706, B2 => 
                           n25243, ZN => n14216);
   U822 : OAI22_X1 port map( A1 => n18331, A2 => n25209, B1 => n19705, B2 => 
                           n25242, ZN => n14217);
   U823 : OAI22_X1 port map( A1 => n18339, A2 => n25202, B1 => n19704, B2 => 
                           n25225, ZN => n14219);
   U824 : OAI22_X1 port map( A1 => n18339, A2 => n25195, B1 => n19703, B2 => 
                           n25225, ZN => n14221);
   U825 : OAI22_X1 port map( A1 => n18344, A2 => n25209, B1 => n19702, B2 => 
                           n25238, ZN => n14222);
   U826 : OAI22_X1 port map( A1 => n18343, A2 => n25209, B1 => n19701, B2 => 
                           n25236, ZN => n14223);
   U827 : OAI22_X1 port map( A1 => n18342, A2 => n25209, B1 => n19700, B2 => 
                           n25241, ZN => n14225);
   U828 : OAI22_X1 port map( A1 => n18341, A2 => n25209, B1 => n19699, B2 => 
                           n25227, ZN => n14226);
   U829 : OAI22_X1 port map( A1 => n18340, A2 => n25209, B1 => n19698, B2 => 
                           n25240, ZN => n14227);
   U830 : OAI22_X1 port map( A1 => n18339, A2 => n25209, B1 => n19697, B2 => 
                           n25225, ZN => n14228);
   U831 : OAI22_X1 port map( A1 => n18338, A2 => n25206, B1 => n19696, B2 => 
                           n25214, ZN => n14230);
   U832 : OAI22_X1 port map( A1 => n18338, A2 => n25228, B1 => n19695, B2 => 
                           n25214, ZN => n14231);
   U833 : OAI22_X1 port map( A1 => n18338, A2 => n25212, B1 => n19694, B2 => 
                           n25214, ZN => n14232);
   U834 : OAI22_X1 port map( A1 => n18337, A2 => n25210, B1 => n19693, B2 => 
                           n25235, ZN => n14233);
   U835 : OAI22_X1 port map( A1 => n18335, A2 => n25210, B1 => n19692, B2 => 
                           n25239, ZN => n14234);
   U836 : OAI22_X1 port map( A1 => n18334, A2 => n25210, B1 => n19691, B2 => 
                           n25244, ZN => n14235);
   U837 : OAI22_X1 port map( A1 => n18333, A2 => n25210, B1 => n19690, B2 => 
                           n25213, ZN => n14236);
   U838 : OAI22_X1 port map( A1 => n18332, A2 => n25210, B1 => n19689, B2 => 
                           n25243, ZN => n14237);
   U839 : OAI22_X1 port map( A1 => n18331, A2 => n25210, B1 => n19688, B2 => 
                           n25242, ZN => n14238);
   U840 : OAI22_X1 port map( A1 => n18338, A2 => n25229, B1 => n19687, B2 => 
                           n25214, ZN => n14239);
   U841 : OAI22_X1 port map( A1 => n18338, A2 => n25230, B1 => n19686, B2 => 
                           n25214, ZN => n14240);
   U842 : OAI22_X1 port map( A1 => n18338, A2 => n25203, B1 => n19685, B2 => 
                           n25214, ZN => n14242);
   U843 : OAI22_X1 port map( A1 => n18338, A2 => n25226, B1 => n19684, B2 => 
                           n25214, ZN => n14243);
   U844 : OAI22_X1 port map( A1 => n18344, A2 => n25210, B1 => n19683, B2 => 
                           n25238, ZN => n14244);
   U845 : OAI22_X1 port map( A1 => n18344, A2 => n25211, B1 => n19682, B2 => 
                           n25238, ZN => n14245);
   U846 : OAI22_X1 port map( A1 => n18343, A2 => n25211, B1 => n19681, B2 => 
                           n25236, ZN => n14246);
   U847 : OAI22_X1 port map( A1 => n18342, A2 => n25211, B1 => n19680, B2 => 
                           n25241, ZN => n14248);
   U848 : OAI22_X1 port map( A1 => n18341, A2 => n25211, B1 => n19679, B2 => 
                           n25227, ZN => n14249);
   U849 : OAI22_X1 port map( A1 => n18334, A2 => n25211, B1 => n19678, B2 => 
                           n25244, ZN => n14250);
   U850 : OAI22_X1 port map( A1 => n18340, A2 => n25211, B1 => n19677, B2 => 
                           n25240, ZN => n14251);
   U851 : OAI22_X1 port map( A1 => n18339, A2 => n25211, B1 => n19676, B2 => 
                           n25225, ZN => n14252);
   U852 : OAI22_X1 port map( A1 => n18343, A2 => n25210, B1 => n19675, B2 => 
                           n25236, ZN => n14254);
   U853 : OAI22_X1 port map( A1 => n18342, A2 => n25210, B1 => n19674, B2 => 
                           n25241, ZN => n14255);
   U854 : OAI22_X1 port map( A1 => n18341, A2 => n25210, B1 => n19673, B2 => 
                           n25227, ZN => n14256);
   U855 : OAI22_X1 port map( A1 => n18335, A2 => n25211, B1 => n19672, B2 => 
                           n25239, ZN => n14257);
   U856 : OAI22_X1 port map( A1 => n18340, A2 => n25210, B1 => n19671, B2 => 
                           n25240, ZN => n14258);
   U857 : OAI22_X1 port map( A1 => n18339, A2 => n25210, B1 => n19670, B2 => 
                           n25225, ZN => n14259);
   U858 : OAI22_X1 port map( A1 => n18338, A2 => n25209, B1 => n19669, B2 => 
                           n25214, ZN => n14260);
   U859 : OAI22_X1 port map( A1 => n18344, A2 => n25212, B1 => n19668, B2 => 
                           n25238, ZN => n14262);
   U860 : OAI22_X1 port map( A1 => n18333, A2 => n25211, B1 => n19667, B2 => 
                           n25213, ZN => n14263);
   U861 : OAI22_X1 port map( A1 => n18332, A2 => n25211, B1 => n19666, B2 => 
                           n25243, ZN => n14264);
   U862 : OAI22_X1 port map( A1 => n18342, A2 => n25226, B1 => n19665, B2 => 
                           n25241, ZN => n14265);
   U863 : OAI22_X1 port map( A1 => n18331, A2 => n25211, B1 => n19664, B2 => 
                           n25242, ZN => n14266);
   U864 : OAI22_X1 port map( A1 => n18338, A2 => n25210, B1 => n19663, B2 => 
                           n25214, ZN => n14268);
   U865 : OAI22_X1 port map( A1 => n18338, A2 => n25223, B1 => n19662, B2 => 
                           n25214, ZN => n14269);
   U866 : OAI22_X1 port map( A1 => n18338, A2 => n25224, B1 => n19661, B2 => 
                           n25214, ZN => n14270);
   U867 : OAI22_X1 port map( A1 => n18338, A2 => n25207, B1 => n19660, B2 => 
                           n25214, ZN => n14272);
   U868 : OAI22_X1 port map( A1 => n18338, A2 => n25222, B1 => n19659, B2 => 
                           n25214, ZN => n14273);
   U869 : OAI22_X1 port map( A1 => n18338, A2 => n25197, B1 => n19658, B2 => 
                           n25214, ZN => n14275);
   U870 : OAI22_X1 port map( A1 => n18338, A2 => n25196, B1 => n19657, B2 => 
                           n25214, ZN => n14277);
   U871 : OAI22_X1 port map( A1 => n18338, A2 => n25204, B1 => n19656, B2 => 
                           n25214, ZN => n14278);
   U872 : OAI22_X1 port map( A1 => n18338, A2 => n25211, B1 => n19655, B2 => 
                           n25214, ZN => n14279);
   U873 : OAI22_X1 port map( A1 => n18338, A2 => n25199, B1 => n19654, B2 => 
                           n25214, ZN => n14281);
   U874 : OAI22_X1 port map( A1 => n18338, A2 => n25198, B1 => n19653, B2 => 
                           n25214, ZN => n14283);
   U875 : OAI22_X1 port map( A1 => n18336, A2 => n25211, B1 => n19652, B2 => 
                           n25231, ZN => n14284);
   U876 : OAI22_X1 port map( A1 => n18337, A2 => n25211, B1 => n19651, B2 => 
                           n25235, ZN => n14286);
   U877 : OAI22_X1 port map( A1 => n18338, A2 => n25200, B1 => n19650, B2 => 
                           n25214, ZN => n14288);
   U878 : OAI22_X1 port map( A1 => n18347, A2 => n25237, B1 => n19649, B2 => 
                           n25232, ZN => n14290);
   U879 : OAI22_X1 port map( A1 => n18346, A2 => n25237, B1 => n19648, B2 => 
                           n25233, ZN => n14292);
   U880 : OAI22_X1 port map( A1 => n18348, A2 => n25237, B1 => n19647, B2 => 
                           n25234, ZN => n14294);
   U881 : OAI22_X1 port map( A1 => n18353, A2 => n25216, B1 => n19646, B2 => 
                           n25215, ZN => n14296);
   U882 : OAI22_X1 port map( A1 => n18343, A2 => n25216, B1 => n19645, B2 => 
                           n25236, ZN => n14297);
   U883 : OAI22_X1 port map( A1 => n18349, A2 => n25216, B1 => n19644, B2 => 
                           n25219, ZN => n14298);
   U884 : OAI22_X1 port map( A1 => n18355, A2 => n25216, B1 => n19643, B2 => 
                           n25221, ZN => n14299);
   U885 : OAI22_X1 port map( A1 => n18341, A2 => n25216, B1 => n19642, B2 => 
                           n25227, ZN => n14300);
   U886 : OAI22_X1 port map( A1 => n18351, A2 => n25216, B1 => n19641, B2 => 
                           n25218, ZN => n14301);
   U887 : OAI22_X1 port map( A1 => n18354, A2 => n25216, B1 => n19640, B2 => 
                           n25217, ZN => n14302);
   U888 : OAI22_X1 port map( A1 => n18357, A2 => n25216, B1 => n19639, B2 => 
                           n25220, ZN => n14303);
   U889 : OAI22_X1 port map( A1 => n18336, A2 => n25216, B1 => n19638, B2 => 
                           n25231, ZN => n14304);
   U890 : OAI22_X1 port map( A1 => n18360, A2 => n25216, B1 => n19637, B2 => 
                           n25193, ZN => n14305);
   U891 : OAI22_X1 port map( A1 => n18359, A2 => n25216, B1 => n19636, B2 => 
                           n25194, ZN => n14307);
   U892 : OAI22_X1 port map( A1 => n18345, A2 => n25237, B1 => n19635, B2 => 
                           n25245, ZN => n14309);
   U893 : OAI22_X1 port map( A1 => n18354, A2 => n25253, B1 => n19634, B2 => 
                           n25217, ZN => n14310);
   U894 : OAI22_X1 port map( A1 => n18351, A2 => n25253, B1 => n19633, B2 => 
                           n25218, ZN => n14311);
   U895 : OAI22_X1 port map( A1 => n18349, A2 => n25253, B1 => n19632, B2 => 
                           n25219, ZN => n14312);
   U896 : OAI22_X1 port map( A1 => n18359, A2 => n25253, B1 => n19631, B2 => 
                           n25194, ZN => n14313);
   U897 : OAI22_X1 port map( A1 => n18354, A2 => n25222, B1 => n19630, B2 => 
                           n25217, ZN => n14315);
   U898 : OAI22_X1 port map( A1 => n18351, A2 => n25222, B1 => n19629, B2 => 
                           n25218, ZN => n14317);
   U899 : OAI22_X1 port map( A1 => n18349, A2 => n25222, B1 => n19628, B2 => 
                           n25219, ZN => n14319);
   U900 : OAI22_X1 port map( A1 => n18359, A2 => n25222, B1 => n19627, B2 => 
                           n25194, ZN => n14321);
   U901 : OAI22_X1 port map( A1 => n18353, A2 => n25253, B1 => n19626, B2 => 
                           n25215, ZN => n14322);
   U902 : OAI22_X1 port map( A1 => n18353, A2 => n25222, B1 => n19625, B2 => 
                           n25215, ZN => n14324);
   U903 : OAI22_X1 port map( A1 => n18357, A2 => n25253, B1 => n19624, B2 => 
                           n25220, ZN => n14325);
   U904 : OAI22_X1 port map( A1 => n18355, A2 => n25253, B1 => n19623, B2 => 
                           n25221, ZN => n14326);
   U905 : OAI22_X1 port map( A1 => n18355, A2 => n25222, B1 => n19622, B2 => 
                           n25221, ZN => n14328);
   U906 : OAI22_X1 port map( A1 => n18360, A2 => n25222, B1 => n19621, B2 => 
                           n25193, ZN => n14329);
   U907 : OAI22_X1 port map( A1 => n18360, A2 => n25253, B1 => n19620, B2 => 
                           n25193, ZN => n14331);
   U908 : OAI22_X1 port map( A1 => n18357, A2 => n25222, B1 => n19619, B2 => 
                           n25220, ZN => n14333);
   U909 : OAI22_X1 port map( A1 => n18349, A2 => n25223, B1 => n19618, B2 => 
                           n25219, ZN => n14335);
   U910 : OAI22_X1 port map( A1 => n18343, A2 => n25223, B1 => n19617, B2 => 
                           n25236, ZN => n14336);
   U911 : OAI22_X1 port map( A1 => n18349, A2 => n25224, B1 => n19616, B2 => 
                           n25219, ZN => n14338);
   U912 : OAI22_X1 port map( A1 => n18351, A2 => n25223, B1 => n19615, B2 => 
                           n25218, ZN => n14339);
   U913 : OAI22_X1 port map( A1 => n18351, A2 => n25224, B1 => n19614, B2 => 
                           n25218, ZN => n14340);
   U914 : OAI22_X1 port map( A1 => n18353, A2 => n25223, B1 => n19613, B2 => 
                           n25215, ZN => n14341);
   U915 : OAI22_X1 port map( A1 => n18354, A2 => n25223, B1 => n19612, B2 => 
                           n25217, ZN => n14342);
   U916 : OAI22_X1 port map( A1 => n18353, A2 => n25224, B1 => n19611, B2 => 
                           n25215, ZN => n14343);
   U917 : OAI22_X1 port map( A1 => n18357, A2 => n25226, B1 => n19610, B2 => 
                           n25220, ZN => n14345);
   U918 : OAI22_X1 port map( A1 => n18354, A2 => n25224, B1 => n19609, B2 => 
                           n25217, ZN => n14346);
   U919 : OAI22_X1 port map( A1 => n18342, A2 => n25223, B1 => n19608, B2 => 
                           n25241, ZN => n14347);
   U920 : OAI22_X1 port map( A1 => n18355, A2 => n25224, B1 => n19607, B2 => 
                           n25221, ZN => n14348);
   U921 : OAI22_X1 port map( A1 => n18357, A2 => n25224, B1 => n19606, B2 => 
                           n25220, ZN => n14349);
   U922 : OAI22_X1 port map( A1 => n18359, A2 => n25224, B1 => n19605, B2 => 
                           n25194, ZN => n14350);
   U923 : OAI22_X1 port map( A1 => n18360, A2 => n25224, B1 => n19604, B2 => 
                           n25193, ZN => n14351);
   U924 : OAI22_X1 port map( A1 => n18342, A2 => n25224, B1 => n19603, B2 => 
                           n25241, ZN => n14352);
   U925 : OAI22_X1 port map( A1 => n18339, A2 => n25237, B1 => n19602, B2 => 
                           n25225, ZN => n14354);
   U926 : OAI22_X1 port map( A1 => n18343, A2 => n25224, B1 => n19601, B2 => 
                           n25236, ZN => n14356);
   U927 : OAI22_X1 port map( A1 => n18355, A2 => n25226, B1 => n19600, B2 => 
                           n25221, ZN => n14357);
   U928 : OAI22_X1 port map( A1 => n18360, A2 => n25223, B1 => n19599, B2 => 
                           n25193, ZN => n14359);
   U929 : OAI22_X1 port map( A1 => n18343, A2 => n25222, B1 => n19598, B2 => 
                           n25236, ZN => n14360);
   U930 : CLKBUF_X1 port map( A => n25227, Z => n25252);
   U931 : OAI22_X1 port map( A1 => n18341, A2 => n25237, B1 => n19597, B2 => 
                           n25252, ZN => n14362);
   U932 : OAI22_X1 port map( A1 => n18330, A2 => n25228, B1 => n19596, B2 => 
                           n25188, ZN => n14364);
   U933 : OAI22_X1 port map( A1 => n18359, A2 => n25223, B1 => n19595, B2 => 
                           n25194, ZN => n14366);
   U934 : OAI22_X1 port map( A1 => n18357, A2 => n25223, B1 => n19594, B2 => 
                           n25220, ZN => n14367);
   U935 : OAI22_X1 port map( A1 => n18332, A2 => n25228, B1 => n19593, B2 => 
                           n25243, ZN => n14368);
   U936 : OAI22_X1 port map( A1 => n18355, A2 => n25228, B1 => n19592, B2 => 
                           n25221, ZN => n14369);
   U937 : OAI22_X1 port map( A1 => n18354, A2 => n25228, B1 => n19591, B2 => 
                           n25217, ZN => n14370);
   U938 : OAI22_X1 port map( A1 => n18353, A2 => n25228, B1 => n19590, B2 => 
                           n25215, ZN => n14371);
   U939 : OAI22_X1 port map( A1 => n18351, A2 => n25228, B1 => n19589, B2 => 
                           n25218, ZN => n14372);
   U940 : OAI22_X1 port map( A1 => n18336, A2 => n25237, B1 => n19588, B2 => 
                           n25231, ZN => n14374);
   U941 : OAI22_X1 port map( A1 => n18349, A2 => n25229, B1 => n19587, B2 => 
                           n25219, ZN => n14376);
   U942 : OAI22_X1 port map( A1 => n18349, A2 => n25228, B1 => n19586, B2 => 
                           n25219, ZN => n14377);
   U943 : OAI22_X1 port map( A1 => n18351, A2 => n25229, B1 => n19585, B2 => 
                           n25218, ZN => n14378);
   U944 : OAI22_X1 port map( A1 => n18353, A2 => n25229, B1 => n19584, B2 => 
                           n25215, ZN => n14379);
   U945 : OAI22_X1 port map( A1 => n18354, A2 => n25229, B1 => n19583, B2 => 
                           n25217, ZN => n14380);
   U946 : OAI22_X1 port map( A1 => n18355, A2 => n25223, B1 => n19582, B2 => 
                           n25221, ZN => n14382);
   U947 : OAI22_X1 port map( A1 => n18336, A2 => n25228, B1 => n19581, B2 => 
                           n25231, ZN => n14383);
   U948 : OAI22_X1 port map( A1 => n18336, A2 => n25230, B1 => n19580, B2 => 
                           n25231, ZN => n14385);
   U949 : OAI22_X1 port map( A1 => n18343, A2 => n25226, B1 => n19579, B2 => 
                           n25236, ZN => n14386);
   U950 : OAI22_X1 port map( A1 => n18355, A2 => n25229, B1 => n19578, B2 => 
                           n25221, ZN => n14387);
   U951 : OAI22_X1 port map( A1 => n18357, A2 => n25229, B1 => n19577, B2 => 
                           n25220, ZN => n14388);
   U952 : OAI22_X1 port map( A1 => n18343, A2 => n25228, B1 => n19576, B2 => 
                           n25236, ZN => n14389);
   U953 : OAI22_X1 port map( A1 => n18332, A2 => n25230, B1 => n19575, B2 => 
                           n25243, ZN => n14390);
   U954 : OAI22_X1 port map( A1 => n18330, A2 => n25230, B1 => n19574, B2 => 
                           n25188, ZN => n14391);
   U955 : OAI22_X1 port map( A1 => n18336, A2 => n25229, B1 => n19573, B2 => 
                           n25231, ZN => n14392);
   U956 : OAI22_X1 port map( A1 => n18343, A2 => n25229, B1 => n19572, B2 => 
                           n25236, ZN => n14393);
   U957 : OAI22_X1 port map( A1 => n18330, A2 => n25229, B1 => n19571, B2 => 
                           n25188, ZN => n14394);
   U958 : OAI22_X1 port map( A1 => n18332, A2 => n25229, B1 => n19570, B2 => 
                           n25243, ZN => n14396);
   U959 : OAI22_X1 port map( A1 => n18349, A2 => n25230, B1 => n19569, B2 => 
                           n25219, ZN => n14397);
   U960 : OAI22_X1 port map( A1 => n18343, A2 => n25230, B1 => n19568, B2 => 
                           n25236, ZN => n14398);
   U961 : OAI22_X1 port map( A1 => n18351, A2 => n25230, B1 => n19567, B2 => 
                           n25218, ZN => n14399);
   U962 : OAI22_X1 port map( A1 => n18357, A2 => n25228, B1 => n19566, B2 => 
                           n25220, ZN => n14401);
   U963 : OAI22_X1 port map( A1 => n18353, A2 => n25230, B1 => n19565, B2 => 
                           n25215, ZN => n14402);
   U964 : OAI22_X1 port map( A1 => n18354, A2 => n25230, B1 => n19564, B2 => 
                           n25217, ZN => n14403);
   U965 : OAI22_X1 port map( A1 => n18354, A2 => n25226, B1 => n19563, B2 => 
                           n25217, ZN => n14405);
   U966 : OAI22_X1 port map( A1 => n18357, A2 => n25230, B1 => n19562, B2 => 
                           n25220, ZN => n14407);
   U967 : OAI22_X1 port map( A1 => n18353, A2 => n25226, B1 => n19561, B2 => 
                           n25215, ZN => n14409);
   U968 : OAI22_X1 port map( A1 => n18349, A2 => n25226, B1 => n19560, B2 => 
                           n25219, ZN => n14411);
   U969 : OAI22_X1 port map( A1 => n18342, A2 => n25222, B1 => n19559, B2 => 
                           n25241, ZN => n14413);
   U970 : OAI22_X1 port map( A1 => n18330, A2 => n25226, B1 => n19558, B2 => 
                           n25188, ZN => n14415);
   U971 : OAI22_X1 port map( A1 => n18332, A2 => n25226, B1 => n19557, B2 => 
                           n25243, ZN => n14416);
   U972 : OAI22_X1 port map( A1 => n18336, A2 => n25226, B1 => n19556, B2 => 
                           n25231, ZN => n14418);
   U973 : OAI22_X1 port map( A1 => n18351, A2 => n25226, B1 => n19555, B2 => 
                           n25218, ZN => n14421);
   U974 : OAI22_X1 port map( A1 => n18355, A2 => n25230, B1 => n19554, B2 => 
                           n25221, ZN => n14424);
   U975 : OAI22_X1 port map( A1 => n18346, A2 => n25249, B1 => n19553, B2 => 
                           n25233, ZN => n14425);
   U976 : OAI22_X1 port map( A1 => n18347, A2 => n25249, B1 => n19552, B2 => 
                           n25232, ZN => n14426);
   U977 : OAI22_X1 port map( A1 => n18347, A2 => n25222, B1 => n19551, B2 => 
                           n25232, ZN => n14427);
   U978 : OAI22_X1 port map( A1 => n18347, A2 => n25209, B1 => n19550, B2 => 
                           n25232, ZN => n14428);
   U979 : OAI22_X1 port map( A1 => n18347, A2 => n25204, B1 => n19549, B2 => 
                           n25232, ZN => n14429);
   U980 : OAI22_X1 port map( A1 => n18346, A2 => n25222, B1 => n19548, B2 => 
                           n25233, ZN => n14430);
   U981 : OAI22_X1 port map( A1 => n18346, A2 => n25209, B1 => n19547, B2 => 
                           n25233, ZN => n14431);
   U982 : OAI22_X1 port map( A1 => n18348, A2 => n25249, B1 => n19546, B2 => 
                           n25234, ZN => n14432);
   U983 : OAI22_X1 port map( A1 => n18347, A2 => n25247, B1 => n19545, B2 => 
                           n25232, ZN => n14433);
   U984 : OAI22_X1 port map( A1 => n18348, A2 => n25222, B1 => n19544, B2 => 
                           n25234, ZN => n14434);
   U985 : OAI22_X1 port map( A1 => n18348, A2 => n25251, B1 => n19543, B2 => 
                           n25234, ZN => n14435);
   U986 : OAI22_X1 port map( A1 => n18348, A2 => n25253, B1 => n19542, B2 => 
                           n25234, ZN => n14436);
   U987 : OAI22_X1 port map( A1 => n18348, A2 => n25247, B1 => n19541, B2 => 
                           n25234, ZN => n14437);
   U988 : OAI22_X1 port map( A1 => n18347, A2 => n25248, B1 => n19540, B2 => 
                           n25232, ZN => n14438);
   U989 : OAI22_X1 port map( A1 => n18347, A2 => n25253, B1 => n19539, B2 => 
                           n25232, ZN => n14439);
   U990 : OAI22_X1 port map( A1 => n18347, A2 => n25250, B1 => n19538, B2 => 
                           n25232, ZN => n14440);
   U991 : OAI22_X1 port map( A1 => n18346, A2 => n25253, B1 => n19537, B2 => 
                           n25233, ZN => n14441);
   U992 : OAI22_X1 port map( A1 => n18348, A2 => n25246, B1 => n19536, B2 => 
                           n25234, ZN => n14442);
   U993 : OAI22_X1 port map( A1 => n18348, A2 => n25204, B1 => n19535, B2 => 
                           n25234, ZN => n14443);
   U994 : OAI22_X1 port map( A1 => n18346, A2 => n25247, B1 => n19534, B2 => 
                           n25233, ZN => n14444);
   U995 : OAI22_X1 port map( A1 => n18346, A2 => n25204, B1 => n19533, B2 => 
                           n25233, ZN => n14445);
   U996 : OAI22_X1 port map( A1 => n18348, A2 => n25209, B1 => n19532, B2 => 
                           n25234, ZN => n14446);
   U997 : OAI22_X1 port map( A1 => n18346, A2 => n25248, B1 => n19531, B2 => 
                           n25233, ZN => n14447);
   U998 : OAI22_X1 port map( A1 => n18347, A2 => n25246, B1 => n19530, B2 => 
                           n25232, ZN => n14448);
   U999 : OAI22_X1 port map( A1 => n18348, A2 => n25248, B1 => n19529, B2 => 
                           n25234, ZN => n14449);
   U1000 : OAI22_X1 port map( A1 => n18347, A2 => n25251, B1 => n19528, B2 => 
                           n25232, ZN => n14451);
   U1001 : OAI22_X1 port map( A1 => n18346, A2 => n25251, B1 => n19527, B2 => 
                           n25233, ZN => n14452);
   U1002 : OAI22_X1 port map( A1 => n18346, A2 => n25246, B1 => n19526, B2 => 
                           n25233, ZN => n14453);
   U1003 : OAI22_X1 port map( A1 => n18348, A2 => n25250, B1 => n19525, B2 => 
                           n25234, ZN => n14455);
   U1004 : OAI22_X1 port map( A1 => n18346, A2 => n25250, B1 => n19524, B2 => 
                           n25233, ZN => n14457);
   U1005 : CLKBUF_X1 port map( A => n25235, Z => n25254);
   U1006 : OAI22_X1 port map( A1 => n18337, A2 => n25237, B1 => n19523, B2 => 
                           n25254, ZN => n14459);
   U1007 : OAI22_X1 port map( A1 => n18333, A2 => n25237, B1 => n19522, B2 => 
                           n25213, ZN => n14461);
   U1008 : OAI22_X1 port map( A1 => n18343, A2 => n25237, B1 => n19521, B2 => 
                           n25236, ZN => n14463);
   U1009 : OAI22_X1 port map( A1 => n18344, A2 => n25237, B1 => n19520, B2 => 
                           n25238, ZN => n14465);
   U1010 : OAI22_X1 port map( A1 => n18335, A2 => n25237, B1 => n19519, B2 => 
                           n25239, ZN => n14467);
   U1011 : OAI22_X1 port map( A1 => n18340, A2 => n25237, B1 => n19518, B2 => 
                           n25240, ZN => n14469);
   U1012 : OAI22_X1 port map( A1 => n18338, A2 => n25237, B1 => n19517, B2 => 
                           n25214, ZN => n14471);
   U1013 : OAI22_X1 port map( A1 => n18342, A2 => n25237, B1 => n19516, B2 => 
                           n25241, ZN => n14473);
   U1014 : OAI22_X1 port map( A1 => n18331, A2 => n25237, B1 => n19515, B2 => 
                           n25242, ZN => n14475);
   U1015 : OAI22_X1 port map( A1 => n18332, A2 => n25237, B1 => n19514, B2 => 
                           n25243, ZN => n14477);
   U1016 : OAI22_X1 port map( A1 => n18334, A2 => n25237, B1 => n19513, B2 => 
                           n25244, ZN => n14480);
   U1017 : OAI22_X1 port map( A1 => n18345, A2 => n25247, B1 => n19512, B2 => 
                           n25245, ZN => n14481);
   U1018 : OAI22_X1 port map( A1 => n18345, A2 => n25253, B1 => n19511, B2 => 
                           n25245, ZN => n14482);
   U1019 : OAI22_X1 port map( A1 => n18345, A2 => n25249, B1 => n19510, B2 => 
                           n25245, ZN => n14483);
   U1020 : OAI22_X1 port map( A1 => n18345, A2 => n25204, B1 => n19509, B2 => 
                           n25245, ZN => n14485);
   U1021 : OAI22_X1 port map( A1 => n18345, A2 => n25250, B1 => n19508, B2 => 
                           n25245, ZN => n14486);
   U1022 : OAI22_X1 port map( A1 => n18345, A2 => n25251, B1 => n19507, B2 => 
                           n25245, ZN => n14487);
   U1023 : OAI22_X1 port map( A1 => n18345, A2 => n25222, B1 => n19506, B2 => 
                           n25245, ZN => n14489);
   U1024 : OAI22_X1 port map( A1 => n18345, A2 => n25209, B1 => n19505, B2 => 
                           n25245, ZN => n14491);
   U1025 : OAI22_X1 port map( A1 => n18345, A2 => n25248, B1 => n19504, B2 => 
                           n25245, ZN => n14492);
   U1026 : OAI22_X1 port map( A1 => n18345, A2 => n25246, B1 => n19503, B2 => 
                           n25245, ZN => n14494);
   U1027 : OAI22_X1 port map( A1 => n18342, A2 => n25251, B1 => n19502, B2 => 
                           n25241, ZN => n14495);
   U1028 : OAI22_X1 port map( A1 => n18342, A2 => n25253, B1 => n19501, B2 => 
                           n25241, ZN => n14496);
   U1029 : OAI22_X1 port map( A1 => n18343, A2 => n25249, B1 => n19500, B2 => 
                           n25236, ZN => n14497);
   U1030 : OAI22_X1 port map( A1 => n18342, A2 => n25248, B1 => n19499, B2 => 
                           n25241, ZN => n14498);
   U1031 : OAI22_X1 port map( A1 => n18343, A2 => n25253, B1 => n19498, B2 => 
                           n25236, ZN => n14500);
   U1032 : OAI22_X1 port map( A1 => n18342, A2 => n25250, B1 => n19497, B2 => 
                           n25241, ZN => n14501);
   U1033 : OAI22_X1 port map( A1 => n18343, A2 => n25250, B1 => n19496, B2 => 
                           n25236, ZN => n14503);
   U1034 : OAI22_X1 port map( A1 => n18342, A2 => n25246, B1 => n19495, B2 => 
                           n25241, ZN => n14504);
   U1035 : OAI22_X1 port map( A1 => n18342, A2 => n25249, B1 => n19494, B2 => 
                           n25241, ZN => n14506);
   U1036 : OAI22_X1 port map( A1 => n18343, A2 => n25247, B1 => n19493, B2 => 
                           n25236, ZN => n14507);
   U1037 : OAI22_X1 port map( A1 => n18343, A2 => n25251, B1 => n19492, B2 => 
                           n25236, ZN => n14509);
   U1038 : OAI22_X1 port map( A1 => n18342, A2 => n25247, B1 => n19491, B2 => 
                           n25241, ZN => n14512);
   U1039 : OAI22_X1 port map( A1 => n18343, A2 => n25246, B1 => n19490, B2 => 
                           n25236, ZN => n14514);
   U1040 : OAI22_X1 port map( A1 => n18343, A2 => n25248, B1 => n19489, B2 => 
                           n25236, ZN => n14517);
   U1041 : OAI22_X1 port map( A1 => n18339, A2 => n25248, B1 => n19488, B2 => 
                           n25225, ZN => n14518);
   U1042 : OAI22_X1 port map( A1 => n18337, A2 => n25248, B1 => n19487, B2 => 
                           n25254, ZN => n14519);
   U1043 : OAI22_X1 port map( A1 => n18340, A2 => n25246, B1 => n19486, B2 => 
                           n25240, ZN => n14520);
   U1044 : OAI22_X1 port map( A1 => n18339, A2 => n25246, B1 => n19485, B2 => 
                           n25225, ZN => n14521);
   U1045 : OAI22_X1 port map( A1 => n18337, A2 => n25246, B1 => n19484, B2 => 
                           n25254, ZN => n14522);
   U1046 : OAI22_X1 port map( A1 => n18336, A2 => n25248, B1 => n19483, B2 => 
                           n25231, ZN => n14523);
   U1047 : OAI22_X1 port map( A1 => n18336, A2 => n25246, B1 => n19482, B2 => 
                           n25231, ZN => n14524);
   U1048 : OAI22_X1 port map( A1 => n18339, A2 => n25247, B1 => n19481, B2 => 
                           n25225, ZN => n14525);
   U1049 : OAI22_X1 port map( A1 => n18340, A2 => n25249, B1 => n19480, B2 => 
                           n25240, ZN => n14526);
   U1050 : OAI22_X1 port map( A1 => n18337, A2 => n25247, B1 => n19479, B2 => 
                           n25254, ZN => n14527);
   U1051 : OAI22_X1 port map( A1 => n18336, A2 => n25247, B1 => n19478, B2 => 
                           n25231, ZN => n14528);
   U1052 : OAI22_X1 port map( A1 => n18339, A2 => n25249, B1 => n19477, B2 => 
                           n25225, ZN => n14529);
   U1053 : OAI22_X1 port map( A1 => n18338, A2 => n25247, B1 => n19476, B2 => 
                           n25214, ZN => n14530);
   U1054 : OAI22_X1 port map( A1 => n18331, A2 => n25247, B1 => n19475, B2 => 
                           n25242, ZN => n14531);
   U1055 : OAI22_X1 port map( A1 => n18331, A2 => n25246, B1 => n19474, B2 => 
                           n25242, ZN => n14532);
   U1056 : OAI22_X1 port map( A1 => n18341, A2 => n25253, B1 => n19473, B2 => 
                           n25252, ZN => n14533);
   U1057 : OAI22_X1 port map( A1 => n18341, A2 => n25248, B1 => n19472, B2 => 
                           n25252, ZN => n14534);
   U1058 : OAI22_X1 port map( A1 => n18332, A2 => n25246, B1 => n19471, B2 => 
                           n25243, ZN => n14535);
   U1059 : OAI22_X1 port map( A1 => n18334, A2 => n25246, B1 => n19470, B2 => 
                           n25244, ZN => n14536);
   U1060 : OAI22_X1 port map( A1 => n18332, A2 => n25247, B1 => n19469, B2 => 
                           n25243, ZN => n14537);
   U1061 : OAI22_X1 port map( A1 => n18334, A2 => n25247, B1 => n19468, B2 => 
                           n25244, ZN => n14538);
   U1062 : OAI22_X1 port map( A1 => n18332, A2 => n25248, B1 => n19467, B2 => 
                           n25243, ZN => n14539);
   U1063 : OAI22_X1 port map( A1 => n18334, A2 => n25248, B1 => n19466, B2 => 
                           n25244, ZN => n14540);
   U1064 : OAI22_X1 port map( A1 => n18338, A2 => n25248, B1 => n19465, B2 => 
                           n25214, ZN => n14541);
   U1065 : OAI22_X1 port map( A1 => n18331, A2 => n25248, B1 => n19464, B2 => 
                           n25242, ZN => n14542);
   U1066 : OAI22_X1 port map( A1 => n18341, A2 => n25247, B1 => n19463, B2 => 
                           n25252, ZN => n14543);
   U1067 : OAI22_X1 port map( A1 => n18341, A2 => n25249, B1 => n19462, B2 => 
                           n25252, ZN => n14544);
   U1068 : OAI22_X1 port map( A1 => n18341, A2 => n25246, B1 => n19461, B2 => 
                           n25252, ZN => n14545);
   U1069 : OAI22_X1 port map( A1 => n18334, A2 => n25250, B1 => n19460, B2 => 
                           n25244, ZN => n14546);
   U1070 : OAI22_X1 port map( A1 => n18344, A2 => n25246, B1 => n19459, B2 => 
                           n25238, ZN => n14547);
   U1071 : OAI22_X1 port map( A1 => n18336, A2 => n25250, B1 => n19458, B2 => 
                           n25231, ZN => n14548);
   U1072 : OAI22_X1 port map( A1 => n18344, A2 => n25249, B1 => n19457, B2 => 
                           n25238, ZN => n14549);
   U1073 : OAI22_X1 port map( A1 => n18337, A2 => n25250, B1 => n19456, B2 => 
                           n25254, ZN => n14550);
   U1074 : OAI22_X1 port map( A1 => n18339, A2 => n25250, B1 => n19455, B2 => 
                           n25225, ZN => n14551);
   U1075 : OAI22_X1 port map( A1 => n18344, A2 => n25247, B1 => n19454, B2 => 
                           n25238, ZN => n14552);
   U1076 : OAI22_X1 port map( A1 => n18344, A2 => n25248, B1 => n19453, B2 => 
                           n25238, ZN => n14553);
   U1077 : OAI22_X1 port map( A1 => n18344, A2 => n25250, B1 => n19452, B2 => 
                           n25238, ZN => n14554);
   U1078 : OAI22_X1 port map( A1 => n18335, A2 => n25246, B1 => n19451, B2 => 
                           n25239, ZN => n14555);
   U1079 : OAI22_X1 port map( A1 => n18341, A2 => n25250, B1 => n19450, B2 => 
                           n25252, ZN => n14556);
   U1080 : OAI22_X1 port map( A1 => n18338, A2 => n25246, B1 => n19449, B2 => 
                           n25214, ZN => n14557);
   U1081 : OAI22_X1 port map( A1 => n18338, A2 => n25250, B1 => n19448, B2 => 
                           n25214, ZN => n14558);
   U1082 : OAI22_X1 port map( A1 => n18331, A2 => n25250, B1 => n19447, B2 => 
                           n25242, ZN => n14559);
   U1083 : OAI22_X1 port map( A1 => n18335, A2 => n25247, B1 => n19446, B2 => 
                           n25239, ZN => n14560);
   U1084 : OAI22_X1 port map( A1 => n18332, A2 => n25250, B1 => n19445, B2 => 
                           n25243, ZN => n14561);
   U1085 : OAI22_X1 port map( A1 => n18333, A2 => n25250, B1 => n19444, B2 => 
                           n25213, ZN => n14562);
   U1086 : OAI22_X1 port map( A1 => n18333, A2 => n25248, B1 => n19443, B2 => 
                           n25213, ZN => n14563);
   U1087 : OAI22_X1 port map( A1 => n18333, A2 => n25247, B1 => n19442, B2 => 
                           n25213, ZN => n14564);
   U1088 : OAI22_X1 port map( A1 => n18334, A2 => n25251, B1 => n19441, B2 => 
                           n25244, ZN => n14565);
   U1089 : OAI22_X1 port map( A1 => n18335, A2 => n25248, B1 => n19440, B2 => 
                           n25239, ZN => n14566);
   U1090 : OAI22_X1 port map( A1 => n18335, A2 => n25250, B1 => n19439, B2 => 
                           n25239, ZN => n14567);
   U1091 : OAI22_X1 port map( A1 => n18335, A2 => n25251, B1 => n19438, B2 => 
                           n25239, ZN => n14568);
   U1092 : OAI22_X1 port map( A1 => n18332, A2 => n25251, B1 => n19437, B2 => 
                           n25243, ZN => n14569);
   U1093 : OAI22_X1 port map( A1 => n18336, A2 => n25251, B1 => n19436, B2 => 
                           n25231, ZN => n14570);
   U1094 : OAI22_X1 port map( A1 => n18337, A2 => n25251, B1 => n19435, B2 => 
                           n25254, ZN => n14571);
   U1095 : OAI22_X1 port map( A1 => n18340, A2 => n25253, B1 => n19434, B2 => 
                           n25240, ZN => n14572);
   U1096 : OAI22_X1 port map( A1 => n18340, A2 => n25250, B1 => n19433, B2 => 
                           n25240, ZN => n14574);
   U1097 : OAI22_X1 port map( A1 => n18338, A2 => n25249, B1 => n19432, B2 => 
                           n25214, ZN => n14575);
   U1098 : OAI22_X1 port map( A1 => n18339, A2 => n25251, B1 => n19431, B2 => 
                           n25225, ZN => n14576);
   U1099 : OAI22_X1 port map( A1 => n18337, A2 => n25249, B1 => n19430, B2 => 
                           n25254, ZN => n14577);
   U1100 : OAI22_X1 port map( A1 => n18336, A2 => n25249, B1 => n19429, B2 => 
                           n25231, ZN => n14578);
   U1101 : OAI22_X1 port map( A1 => n18340, A2 => n25251, B1 => n19428, B2 => 
                           n25240, ZN => n14579);
   U1102 : OAI22_X1 port map( A1 => n18341, A2 => n25251, B1 => n19427, B2 => 
                           n25252, ZN => n14581);
   U1103 : OAI22_X1 port map( A1 => n18344, A2 => n25251, B1 => n19426, B2 => 
                           n25238, ZN => n14582);
   U1104 : OAI22_X1 port map( A1 => n18339, A2 => n25253, B1 => n19425, B2 => 
                           n25225, ZN => n14584);
   U1105 : OAI22_X1 port map( A1 => n18331, A2 => n25249, B1 => n19424, B2 => 
                           n25242, ZN => n14585);
   U1106 : OAI22_X1 port map( A1 => n18335, A2 => n25249, B1 => n19423, B2 => 
                           n25239, ZN => n14586);
   U1107 : OAI22_X1 port map( A1 => n18334, A2 => n25253, B1 => n19422, B2 => 
                           n25244, ZN => n14587);
   U1108 : OAI22_X1 port map( A1 => n18334, A2 => n25249, B1 => n19421, B2 => 
                           n25244, ZN => n14589);
   U1109 : OAI22_X1 port map( A1 => n18333, A2 => n25253, B1 => n19420, B2 => 
                           n25213, ZN => n14590);
   U1110 : OAI22_X1 port map( A1 => n18333, A2 => n25246, B1 => n19419, B2 => 
                           n25213, ZN => n14592);
   U1111 : OAI22_X1 port map( A1 => n18333, A2 => n25249, B1 => n19418, B2 => 
                           n25213, ZN => n14593);
   U1112 : OAI22_X1 port map( A1 => n18332, A2 => n25249, B1 => n19417, B2 => 
                           n25243, ZN => n14595);
   U1113 : OAI22_X1 port map( A1 => n18331, A2 => n25251, B1 => n19416, B2 => 
                           n25242, ZN => n14596);
   U1114 : OAI22_X1 port map( A1 => n18337, A2 => n25253, B1 => n19415, B2 => 
                           n25254, ZN => n14598);
   U1115 : OAI22_X1 port map( A1 => n18340, A2 => n25247, B1 => n19414, B2 => 
                           n25240, ZN => n14600);
   U1116 : OAI22_X1 port map( A1 => n18333, A2 => n25251, B1 => n19413, B2 => 
                           n25213, ZN => n14602);
   U1117 : OAI22_X1 port map( A1 => n18340, A2 => n25248, B1 => n19412, B2 => 
                           n25240, ZN => n14605);
   U1118 : OAI22_X1 port map( A1 => n18332, A2 => n25253, B1 => n19411, B2 => 
                           n25243, ZN => n14607);
   U1119 : OAI22_X1 port map( A1 => n18331, A2 => n25253, B1 => n19410, B2 => 
                           n25242, ZN => n14609);
   U1120 : OAI22_X1 port map( A1 => n18338, A2 => n25251, B1 => n19409, B2 => 
                           n25214, ZN => n14611);
   U1121 : OAI22_X1 port map( A1 => n18344, A2 => n25253, B1 => n19408, B2 => 
                           n25238, ZN => n14613);
   U1122 : OAI22_X1 port map( A1 => n18338, A2 => n25253, B1 => n19407, B2 => 
                           n25214, ZN => n14615);
   U1123 : OAI22_X1 port map( A1 => n18335, A2 => n25253, B1 => n19406, B2 => 
                           n25239, ZN => n14617);
   U1124 : OAI22_X1 port map( A1 => n18336, A2 => n25253, B1 => n19405, B2 => 
                           n25231, ZN => n14620);
   U1125 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1),
                           ZN => n14632);
   U1126 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n19404, ZN => 
                           n25261);
   U1127 : NOR2_X1 port map( A1 => n20466, A2 => n25261, ZN => n25259);
   U1128 : NAND2_X1 port map( A1 => n18284, A2 => n25259, ZN => n10102);
   U1129 : INV_X1 port map( A => ADD_WR(0), ZN => n25255);
   U1130 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n25255, ZN
                           => n14633);
   U1131 : NAND2_X1 port map( A1 => n25259, A2 => n18283, ZN => n10101);
   U1132 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n25255, ZN => n25256);
   U1133 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n25256, ZN => n14634);
   U1134 : NAND2_X1 port map( A1 => n25259, A2 => n18358, ZN => n10100);
   U1135 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n25257);
   U1136 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n25257, ZN => n14635);
   U1137 : NAND2_X1 port map( A1 => n25259, A2 => n18356, ZN => n10099);
   U1138 : INV_X1 port map( A => ADD_WR(2), ZN => n25258);
   U1139 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n25258, ZN
                           => n14636);
   U1140 : NAND2_X1 port map( A1 => n25259, A2 => n18282, ZN => n10098);
   U1141 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n25255, A3 => n25258, ZN =>
                           n14637);
   U1142 : NAND2_X1 port map( A1 => n25259, A2 => n18281, ZN => n10097);
   U1143 : NOR2_X1 port map( A1 => n25258, A2 => n25256, ZN => n14638);
   U1144 : NAND2_X1 port map( A1 => n25259, A2 => n18352, ZN => n10096);
   U1145 : NOR2_X1 port map( A1 => n25258, A2 => n25257, ZN => n14640);
   U1146 : NAND2_X1 port map( A1 => n25259, A2 => n18350, ZN => n10095);
   U1147 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n20465, ZN => 
                           n25263);
   U1148 : NOR2_X1 port map( A1 => n20466, A2 => n25263, ZN => n25260);
   U1149 : NAND2_X1 port map( A1 => n18284, A2 => n25260, ZN => n10094);
   U1150 : NAND2_X1 port map( A1 => n18283, A2 => n25260, ZN => n10093);
   U1151 : NAND2_X1 port map( A1 => n18358, A2 => n25260, ZN => n10092);
   U1152 : NAND2_X1 port map( A1 => n18356, A2 => n25260, ZN => n10091);
   U1153 : NAND2_X1 port map( A1 => n18282, A2 => n25260, ZN => n10090);
   U1154 : NAND2_X1 port map( A1 => n18281, A2 => n25260, ZN => n10089);
   U1155 : NAND2_X1 port map( A1 => n18352, A2 => n25260, ZN => n10088);
   U1156 : NAND2_X1 port map( A1 => n18350, A2 => n25260, ZN => n10087);
   U1157 : NOR2_X1 port map( A1 => n19403, A2 => n25261, ZN => n25262);
   U1158 : NAND2_X1 port map( A1 => n18284, A2 => n25262, ZN => n10086);
   U1159 : NAND2_X1 port map( A1 => n18283, A2 => n25262, ZN => n10085);
   U1160 : NAND2_X1 port map( A1 => n18358, A2 => n25262, ZN => n10084);
   U1161 : NAND2_X1 port map( A1 => n18356, A2 => n25262, ZN => n10083);
   U1162 : NAND2_X1 port map( A1 => n18282, A2 => n25262, ZN => n10082);
   U1163 : NAND2_X1 port map( A1 => n18281, A2 => n25262, ZN => n10081);
   U1164 : NAND2_X1 port map( A1 => n18352, A2 => n25262, ZN => n10080);
   U1165 : NAND2_X1 port map( A1 => n18350, A2 => n25262, ZN => n10079);
   U1166 : NOR2_X1 port map( A1 => n19403, A2 => n25263, ZN => n25264);
   U1167 : NAND2_X1 port map( A1 => n18284, A2 => n25264, ZN => n10078);
   U1168 : NAND2_X1 port map( A1 => n18283, A2 => n25264, ZN => n10077);
   U1169 : NAND2_X1 port map( A1 => n18358, A2 => n25264, ZN => n10076);
   U1170 : NAND2_X1 port map( A1 => n18356, A2 => n25264, ZN => n10075);
   U1171 : NAND2_X1 port map( A1 => n18282, A2 => n25264, ZN => n10074);
   U1172 : NAND2_X1 port map( A1 => n18281, A2 => n25264, ZN => n10073);
   U1173 : NAND2_X1 port map( A1 => n18352, A2 => n25264, ZN => n10072);
   U1174 : NAND2_X1 port map( A1 => n18350, A2 => n25264, ZN => n10071);
   U1175 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => n25266, A3 => n25269, ZN 
                           => n25144);
   U1176 : INV_X1 port map( A => ADD_RD2(3), ZN => n25265);
   U1177 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n25265, ZN => n25271);
   U1178 : NOR2_X1 port map( A1 => n25271, A2 => n25144, ZN => n11175);
   U1179 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n25266,
                           ZN => n25145);
   U1180 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n25270)
                           ;
   U1181 : NOR2_X1 port map( A1 => n25145, A2 => n25270, ZN => n11174);
   U1182 : NOR2_X1 port map( A1 => n25270, A2 => n1521, ZN => n11173);
   U1183 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => 
                           ADD_RD2(2), ZN => n25147);
   U1184 : NOR2_X1 port map( A1 => n25270, A2 => n25147, ZN => n11191);
   U1185 : NOR2_X1 port map( A1 => n25271, A2 => n1521, ZN => n11168);
   U1186 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => n25269, ZN => n25267);
   U1187 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n25267, ZN => n25146);
   U1188 : NOR2_X1 port map( A1 => n25270, A2 => n25146, ZN => n11172);
   U1189 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n25268, ZN => n25143);
   U1190 : NOR2_X1 port map( A1 => n25270, A2 => n25143, ZN => n11166);
   U1191 : NOR2_X1 port map( A1 => n25271, A2 => n25147, ZN => n11165);
   U1192 : NOR2_X1 port map( A1 => n25271, A2 => n1520, ZN => n11167);
   U1193 : NOR2_X1 port map( A1 => n25144, A2 => n25270, ZN => n11190);
   U1194 : NOR2_X1 port map( A1 => n25270, A2 => n1520, ZN => n11157);
   U1195 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n25269,
                           ZN => n25148);
   U1196 : NOR2_X1 port map( A1 => n25270, A2 => n25148, ZN => n11189);
   U1197 : NOR2_X1 port map( A1 => n25271, A2 => n25148, ZN => n11188);
   U1198 : NOR2_X1 port map( A1 => n25271, A2 => n25146, ZN => n11187);
   U1199 : NOR2_X1 port map( A1 => n25271, A2 => n25145, ZN => n11186);
   U1200 : NOR2_X1 port map( A1 => n25271, A2 => n25143, ZN => n11162);
   U1201 : AOI22_X1 port map( A1 => n18977, A2 => n18311, B1 => n19201, B2 => 
                           n18322, ZN => n25275);
   U1202 : CLKBUF_X1 port map( A => n18314, Z => n25982);
   U1203 : CLKBUF_X1 port map( A => n18317, Z => n25950);
   U1204 : AOI22_X1 port map( A1 => n19137, A2 => n25982, B1 => n19105, B2 => 
                           n25950, ZN => n25274);
   U1205 : AOI22_X1 port map( A1 => n19233, A2 => n18319, B1 => n19329, B2 => 
                           n18323, ZN => n25273);
   U1206 : CLKBUF_X1 port map( A => n18320, Z => n25902);
   U1207 : AOI22_X1 port map( A1 => n19297, A2 => n18313, B1 => n18945, B2 => 
                           n25902, ZN => n25272);
   U1208 : NAND4_X1 port map( A1 => n25275, A2 => n25274, A3 => n25273, A4 => 
                           n25272, ZN => n25281);
   U1209 : AOI22_X1 port map( A1 => n18913, A2 => n18309, B1 => n19169, B2 => 
                           n18318, ZN => n25279);
   U1210 : CLKBUF_X1 port map( A => n18316, Z => n25922);
   U1211 : AOI22_X1 port map( A1 => n19041, A2 => n18312, B1 => n18881, B2 => 
                           n25922, ZN => n25278);
   U1212 : CLKBUF_X1 port map( A => n18321, Z => n25974);
   U1213 : CLKBUF_X1 port map( A => n18310, Z => n25829);
   U1214 : AOI22_X1 port map( A1 => n19361, A2 => n25974, B1 => n19073, B2 => 
                           n25829, ZN => n25277);
   U1215 : CLKBUF_X1 port map( A => n18315, Z => n25949);
   U1216 : AOI22_X1 port map( A1 => n19009, A2 => n18324, B1 => n19265, B2 => 
                           n25949, ZN => n25276);
   U1217 : NAND4_X1 port map( A1 => n25279, A2 => n25278, A3 => n25277, A4 => 
                           n25276, ZN => n25280);
   U1218 : NOR2_X1 port map( A1 => n25281, A2 => n25280, ZN => n25293);
   U1219 : NOR3_X1 port map( A1 => n18370, A2 => n20463, A3 => n25828, ZN => 
                           n25734);
   U1220 : CLKBUF_X1 port map( A => n25734, Z => n25780);
   U1221 : INV_X1 port map( A => n25151, ZN => n25797);
   U1222 : CLKBUF_X1 port map( A => n26754, Z => n25994);
   U1223 : AOI22_X1 port map( A1 => n18498, A2 => n25797, B1 => n18562, B2 => 
                           n25994, ZN => n25285);
   U1224 : AOI22_X1 port map( A1 => n18530, A2 => n26757, B1 => n18434, B2 => 
                           n18288, ZN => n25284);
   U1225 : CLKBUF_X1 port map( A => n18291, Z => n25961);
   U1226 : AOI22_X1 port map( A1 => n18594, A2 => n26755, B1 => n18371, B2 => 
                           n25961, ZN => n25283);
   U1227 : INV_X1 port map( A => n25150, ZN => n25992);
   U1228 : AOI22_X1 port map( A1 => n18402, A2 => n25992, B1 => n18466, B2 => 
                           n26756, ZN => n25282);
   U1229 : NAND4_X1 port map( A1 => n25285, A2 => n25284, A3 => n25283, A4 => 
                           n25282, ZN => n25291);
   U1230 : NOR3_X1 port map( A1 => n20463, A2 => n20429, A3 => n25828, ZN => 
                           n25533);
   U1231 : CLKBUF_X1 port map( A => n25533, Z => n26007);
   U1232 : INV_X1 port map( A => n25155, ZN => n25993);
   U1233 : CLKBUF_X1 port map( A => n25993, Z => n25866);
   U1234 : AOI22_X1 port map( A1 => n18721, A2 => n25866, B1 => n18753, B2 => 
                           n26759, ZN => n25289);
   U1235 : AOI22_X1 port map( A1 => n19402, A2 => n18689, B1 => n18785, B2 => 
                           n26757, ZN => n25288);
   U1236 : CLKBUF_X1 port map( A => n26755, Z => n25995);
   U1237 : AOI22_X1 port map( A1 => n19401, A2 => n18625, B1 => n18849, B2 => 
                           n25995, ZN => n25287);
   U1238 : CLKBUF_X1 port map( A => n26754, Z => n25705);
   U1239 : AOI22_X1 port map( A1 => n18657, A2 => n26758, B1 => n18817, B2 => 
                           n25705, ZN => n25286);
   U1240 : NAND4_X1 port map( A1 => n25289, A2 => n25288, A3 => n25287, A4 => 
                           n25286, ZN => n25290);
   U1241 : AOI22_X1 port map( A1 => n25780, A2 => n25291, B1 => n26007, B2 => 
                           n25290, ZN => n25292);
   U1242 : OAI21_X1 port map( B1 => n25828, B2 => n25293, A => n25292, ZN => 
                           OUT2(31));
   U1243 : AOI22_X1 port map( A1 => n18318, A2 => n19170, B1 => n18311, B2 => 
                           n18978, ZN => n25297);
   U1244 : AOI22_X1 port map( A1 => n18309, A2 => n18914, B1 => n18319, B2 => 
                           n19234, ZN => n25296);
   U1245 : AOI22_X1 port map( A1 => n18316, A2 => n18882, B1 => n25950, B2 => 
                           n19106, ZN => n25295);
   U1246 : CLKBUF_X1 port map( A => n18313, Z => n25985);
   U1247 : AOI22_X1 port map( A1 => n25985, A2 => n19298, B1 => n25902, B2 => 
                           n18946, ZN => n25294);
   U1248 : NAND4_X1 port map( A1 => n25297, A2 => n25296, A3 => n25295, A4 => 
                           n25294, ZN => n25303);
   U1249 : CLKBUF_X1 port map( A => n18312, Z => n25928);
   U1250 : AOI22_X1 port map( A1 => n25928, A2 => n19042, B1 => n25974, B2 => 
                           n19362, ZN => n25301);
   U1251 : CLKBUF_X1 port map( A => n18324, Z => n25984);
   U1252 : AOI22_X1 port map( A1 => n25984, A2 => n19010, B1 => n18310, B2 => 
                           n19074, ZN => n25300);
   U1253 : AOI22_X1 port map( A1 => n18314, A2 => n19138, B1 => n18322, B2 => 
                           n19202, ZN => n25299);
   U1254 : AOI22_X1 port map( A1 => n18315, A2 => n19266, B1 => n18323, B2 => 
                           n19330, ZN => n25298);
   U1255 : NAND4_X1 port map( A1 => n25301, A2 => n25300, A3 => n25299, A4 => 
                           n25298, ZN => n25302);
   U1256 : NOR2_X1 port map( A1 => n25303, A2 => n25302, ZN => n25315);
   U1257 : AOI22_X1 port map( A1 => n18595, A2 => n26755, B1 => n18531, B2 => 
                           n26757, ZN => n25307);
   U1258 : AOI22_X1 port map( A1 => n25961, A2 => n18372, B1 => n19402, B2 => 
                           n18435, ZN => n25306);
   U1259 : CLKBUF_X1 port map( A => n25992, Z => n25769);
   U1260 : AOI22_X1 port map( A1 => n18403, A2 => n25769, B1 => n18499, B2 => 
                           n26759, ZN => n25305);
   U1261 : AOI22_X1 port map( A1 => n18467, A2 => n25866, B1 => n18563, B2 => 
                           n26754, ZN => n25304);
   U1262 : NAND4_X1 port map( A1 => n25307, A2 => n25306, A3 => n25305, A4 => 
                           n25304, ZN => n25313);
   U1263 : AOI22_X1 port map( A1 => n18658, A2 => n25769, B1 => n18818, B2 => 
                           n26754, ZN => n25311);
   U1264 : AOI22_X1 port map( A1 => n18722, A2 => n25866, B1 => n18754, B2 => 
                           n26759, ZN => n25310);
   U1265 : CLKBUF_X1 port map( A => n18288, Z => n26001);
   U1266 : AOI22_X1 port map( A1 => n26001, A2 => n18690, B1 => n19401, B2 => 
                           n18626, ZN => n25309);
   U1267 : INV_X1 port map( A => n25154, ZN => n25940);
   U1268 : AOI22_X1 port map( A1 => n18850, A2 => n26755, B1 => n18786, B2 => 
                           n25940, ZN => n25308);
   U1269 : NAND4_X1 port map( A1 => n25311, A2 => n25310, A3 => n25309, A4 => 
                           n25308, ZN => n25312);
   U1270 : AOI22_X1 port map( A1 => n25780, A2 => n25313, B1 => n26007, B2 => 
                           n25312, ZN => n25314);
   U1271 : OAI21_X1 port map( B1 => n25828, B2 => n25315, A => n25314, ZN => 
                           OUT2(30));
   U1272 : CLKBUF_X1 port map( A => n18322, Z => n25976);
   U1273 : AOI22_X1 port map( A1 => n25976, A2 => n19203, B1 => n18320, B2 => 
                           n18947, ZN => n25319);
   U1274 : AOI22_X1 port map( A1 => n18324, A2 => n19011, B1 => n25829, B2 => 
                           n19075, ZN => n25318);
   U1275 : AOI22_X1 port map( A1 => n18316, A2 => n18883, B1 => n25982, B2 => 
                           n19139, ZN => n25317);
   U1276 : AOI22_X1 port map( A1 => n18313, A2 => n19299, B1 => n18319, B2 => 
                           n19235, ZN => n25316);
   U1277 : NAND4_X1 port map( A1 => n25319, A2 => n25318, A3 => n25317, A4 => 
                           n25316, ZN => n25325);
   U1278 : AOI22_X1 port map( A1 => n18317, A2 => n19107, B1 => n18311, B2 => 
                           n18979, ZN => n25323);
   U1279 : AOI22_X1 port map( A1 => n18318, A2 => n19171, B1 => n25974, B2 => 
                           n19363, ZN => n25322);
   U1280 : CLKBUF_X1 port map( A => n18309, Z => n25975);
   U1281 : CLKBUF_X1 port map( A => n18323, Z => n25923);
   U1282 : AOI22_X1 port map( A1 => n25975, A2 => n18915, B1 => n25923, B2 => 
                           n19331, ZN => n25321);
   U1283 : AOI22_X1 port map( A1 => n18312, A2 => n19043, B1 => n25949, B2 => 
                           n19267, ZN => n25320);
   U1284 : NAND4_X1 port map( A1 => n25323, A2 => n25322, A3 => n25321, A4 => 
                           n25320, ZN => n25324);
   U1285 : NOR2_X1 port map( A1 => n25325, A2 => n25324, ZN => n25337);
   U1286 : AOI22_X1 port map( A1 => n18468, A2 => n25866, B1 => n18564, B2 => 
                           n25994, ZN => n25329);
   U1287 : CLKBUF_X1 port map( A => n25797, Z => n25939);
   U1288 : AOI22_X1 port map( A1 => n18596, A2 => n26755, B1 => n18500, B2 => 
                           n25939, ZN => n25328);
   U1289 : AOI22_X1 port map( A1 => n18436, A2 => n19402, B1 => n18532, B2 => 
                           n25940, ZN => n25327);
   U1290 : AOI22_X1 port map( A1 => n18291, A2 => n18373, B1 => n18404, B2 => 
                           n25992, ZN => n25326);
   U1291 : NAND4_X1 port map( A1 => n25329, A2 => n25328, A3 => n25327, A4 => 
                           n25326, ZN => n25335);
   U1292 : AOI22_X1 port map( A1 => n18851, A2 => n26755, B1 => n18787, B2 => 
                           n25940, ZN => n25333);
   U1293 : AOI22_X1 port map( A1 => n18819, A2 => n25994, B1 => n18755, B2 => 
                           n26759, ZN => n25332);
   U1294 : AOI22_X1 port map( A1 => n18288, A2 => n18691, B1 => n19401, B2 => 
                           n18627, ZN => n25331);
   U1295 : AOI22_X1 port map( A1 => n18723, A2 => n26756, B1 => n18659, B2 => 
                           n25992, ZN => n25330);
   U1296 : NAND4_X1 port map( A1 => n25333, A2 => n25332, A3 => n25331, A4 => 
                           n25330, ZN => n25334);
   U1297 : AOI22_X1 port map( A1 => n25780, A2 => n25335, B1 => n26007, B2 => 
                           n25334, ZN => n25336);
   U1298 : OAI21_X1 port map( B1 => n25828, B2 => n25337, A => n25336, ZN => 
                           OUT2(29));
   U1299 : AOI22_X1 port map( A1 => n25949, A2 => n19268, B1 => n18311, B2 => 
                           n18980, ZN => n25341);
   U1300 : AOI22_X1 port map( A1 => n25829, A2 => n19076, B1 => n18323, B2 => 
                           n19332, ZN => n25340);
   U1301 : AOI22_X1 port map( A1 => n18318, A2 => n19172, B1 => n18321, B2 => 
                           n19364, ZN => n25339);
   U1302 : AOI22_X1 port map( A1 => n18316, A2 => n18884, B1 => n18322, B2 => 
                           n19204, ZN => n25338);
   U1303 : NAND4_X1 port map( A1 => n25341, A2 => n25340, A3 => n25339, A4 => 
                           n25338, ZN => n25347);
   U1304 : AOI22_X1 port map( A1 => n18309, A2 => n18916, B1 => n18320, B2 => 
                           n18948, ZN => n25345);
   U1305 : AOI22_X1 port map( A1 => n25984, A2 => n19012, B1 => n25985, B2 => 
                           n19300, ZN => n25344);
   U1306 : CLKBUF_X1 port map( A => n18319, Z => n25981);
   U1307 : AOI22_X1 port map( A1 => n18317, A2 => n19108, B1 => n25981, B2 => 
                           n19236, ZN => n25343);
   U1308 : AOI22_X1 port map( A1 => n18312, A2 => n19044, B1 => n25982, B2 => 
                           n19140, ZN => n25342);
   U1309 : NAND4_X1 port map( A1 => n25345, A2 => n25344, A3 => n25343, A4 => 
                           n25342, ZN => n25346);
   U1310 : NOR2_X1 port map( A1 => n25347, A2 => n25346, ZN => n25359);
   U1311 : AOI22_X1 port map( A1 => n18405, A2 => n26758, B1 => n18501, B2 => 
                           n25797, ZN => n25351);
   U1312 : AOI22_X1 port map( A1 => n18437, A2 => n18288, B1 => n18565, B2 => 
                           n25705, ZN => n25350);
   U1313 : AOI22_X1 port map( A1 => n18597, A2 => n26755, B1 => n18533, B2 => 
                           n26757, ZN => n25349);
   U1314 : AOI22_X1 port map( A1 => n18291, A2 => n18374, B1 => n18469, B2 => 
                           n25993, ZN => n25348);
   U1315 : NAND4_X1 port map( A1 => n25351, A2 => n25350, A3 => n25349, A4 => 
                           n25348, ZN => n25357);
   U1316 : CLKBUF_X1 port map( A => n26755, Z => n26000);
   U1317 : AOI22_X1 port map( A1 => n18724, A2 => n26756, B1 => n18852, B2 => 
                           n26000, ZN => n25355);
   U1318 : AOI22_X1 port map( A1 => n19402, A2 => n18692, B1 => n19401, B2 => 
                           n18628, ZN => n25354);
   U1319 : AOI22_X1 port map( A1 => n18660, A2 => n26758, B1 => n18756, B2 => 
                           n26759, ZN => n25353);
   U1320 : CLKBUF_X1 port map( A => n25940, Z => n25889);
   U1321 : AOI22_X1 port map( A1 => n18788, A2 => n25889, B1 => n18820, B2 => 
                           n25705, ZN => n25352);
   U1322 : NAND4_X1 port map( A1 => n25355, A2 => n25354, A3 => n25353, A4 => 
                           n25352, ZN => n25356);
   U1323 : AOI22_X1 port map( A1 => n25780, A2 => n25357, B1 => n26007, B2 => 
                           n25356, ZN => n25358);
   U1324 : OAI21_X1 port map( B1 => n25828, B2 => n25359, A => n25358, ZN => 
                           OUT2(28));
   U1325 : AOI22_X1 port map( A1 => n25982, A2 => n19141, B1 => n18323, B2 => 
                           n19333, ZN => n25363);
   U1326 : AOI22_X1 port map( A1 => n18312, A2 => n19045, B1 => n25981, B2 => 
                           n19237, ZN => n25362);
   U1327 : AOI22_X1 port map( A1 => n18313, A2 => n19301, B1 => n18320, B2 => 
                           n18949, ZN => n25361);
   U1328 : AOI22_X1 port map( A1 => n18315, A2 => n19269, B1 => n18317, B2 => 
                           n19109, ZN => n25360);
   U1329 : NAND4_X1 port map( A1 => n25363, A2 => n25362, A3 => n25361, A4 => 
                           n25360, ZN => n25369);
   U1330 : AOI22_X1 port map( A1 => n18318, A2 => n19173, B1 => n18321, B2 => 
                           n19365, ZN => n25367);
   U1331 : AOI22_X1 port map( A1 => n18316, A2 => n18885, B1 => n18324, B2 => 
                           n19013, ZN => n25366);
   U1332 : CLKBUF_X1 port map( A => n18311, Z => n25903);
   U1333 : AOI22_X1 port map( A1 => n18309, A2 => n18917, B1 => n25903, B2 => 
                           n18981, ZN => n25365);
   U1334 : AOI22_X1 port map( A1 => n18310, A2 => n19077, B1 => n18322, B2 => 
                           n19205, ZN => n25364);
   U1335 : NAND4_X1 port map( A1 => n25367, A2 => n25366, A3 => n25365, A4 => 
                           n25364, ZN => n25368);
   U1336 : NOR2_X1 port map( A1 => n25369, A2 => n25368, ZN => n25381);
   U1337 : AOI22_X1 port map( A1 => n18470, A2 => n25866, B1 => n18406, B2 => 
                           n25769, ZN => n25373);
   U1338 : AOI22_X1 port map( A1 => n18438, A2 => n19402, B1 => n18566, B2 => 
                           n26754, ZN => n25372);
   U1339 : AOI22_X1 port map( A1 => n18534, A2 => n25889, B1 => n18502, B2 => 
                           n26759, ZN => n25371);
   U1340 : AOI22_X1 port map( A1 => n18375, A2 => n25961, B1 => n18598, B2 => 
                           n26000, ZN => n25370);
   U1341 : NAND4_X1 port map( A1 => n25373, A2 => n25372, A3 => n25371, A4 => 
                           n25370, ZN => n25379);
   U1342 : AOI22_X1 port map( A1 => n18629, A2 => n19401, B1 => n18821, B2 => 
                           n25705, ZN => n25377);
   U1343 : AOI22_X1 port map( A1 => n18789, A2 => n25889, B1 => n18757, B2 => 
                           n26759, ZN => n25376);
   U1344 : AOI22_X1 port map( A1 => n26001, A2 => n18693, B1 => n18725, B2 => 
                           n25993, ZN => n25375);
   U1345 : AOI22_X1 port map( A1 => n18661, A2 => n26758, B1 => n18853, B2 => 
                           n25995, ZN => n25374);
   U1346 : NAND4_X1 port map( A1 => n25377, A2 => n25376, A3 => n25375, A4 => 
                           n25374, ZN => n25378);
   U1347 : AOI22_X1 port map( A1 => n25780, A2 => n25379, B1 => n26007, B2 => 
                           n25378, ZN => n25380);
   U1348 : OAI21_X1 port map( B1 => n25828, B2 => n25381, A => n25380, ZN => 
                           OUT2(27));
   U1349 : AOI22_X1 port map( A1 => n18314, A2 => n19142, B1 => n18323, B2 => 
                           n19334, ZN => n25385);
   U1350 : AOI22_X1 port map( A1 => n18318, A2 => n19174, B1 => n18324, B2 => 
                           n19014, ZN => n25384);
   U1351 : AOI22_X1 port map( A1 => n18309, A2 => n18918, B1 => n18319, B2 => 
                           n19238, ZN => n25383);
   U1352 : AOI22_X1 port map( A1 => n18321, A2 => n19366, B1 => n25902, B2 => 
                           n18950, ZN => n25382);
   U1353 : NAND4_X1 port map( A1 => n25385, A2 => n25384, A3 => n25383, A4 => 
                           n25382, ZN => n25391);
   U1354 : AOI22_X1 port map( A1 => n18310, A2 => n19078, B1 => n25903, B2 => 
                           n18982, ZN => n25389);
   U1355 : AOI22_X1 port map( A1 => n25928, A2 => n19046, B1 => n25950, B2 => 
                           n19110, ZN => n25388);
   U1356 : AOI22_X1 port map( A1 => n18315, A2 => n19270, B1 => n25976, B2 => 
                           n19206, ZN => n25387);
   U1357 : AOI22_X1 port map( A1 => n18316, A2 => n18886, B1 => n18313, B2 => 
                           n19302, ZN => n25386);
   U1358 : NAND4_X1 port map( A1 => n25389, A2 => n25388, A3 => n25387, A4 => 
                           n25386, ZN => n25390);
   U1359 : NOR2_X1 port map( A1 => n25391, A2 => n25390, ZN => n25403);
   U1360 : AOI22_X1 port map( A1 => n18407, A2 => n26758, B1 => n18599, B2 => 
                           n25995, ZN => n25395);
   U1361 : AOI22_X1 port map( A1 => n18376, A2 => n25961, B1 => n18567, B2 => 
                           n26754, ZN => n25394);
   U1362 : AOI22_X1 port map( A1 => n18439, A2 => n18288, B1 => n18503, B2 => 
                           n26759, ZN => n25393);
   U1363 : AOI22_X1 port map( A1 => n18471, A2 => n26756, B1 => n18535, B2 => 
                           n25940, ZN => n25392);
   U1364 : NAND4_X1 port map( A1 => n25395, A2 => n25394, A3 => n25393, A4 => 
                           n25392, ZN => n25401);
   U1365 : AOI22_X1 port map( A1 => n18694, A2 => n19402, B1 => n18662, B2 => 
                           n25992, ZN => n25399);
   U1366 : AOI22_X1 port map( A1 => n18630, A2 => n25961, B1 => n18758, B2 => 
                           n26759, ZN => n25398);
   U1367 : AOI22_X1 port map( A1 => n18726, A2 => n26756, B1 => n18822, B2 => 
                           n26754, ZN => n25397);
   U1368 : AOI22_X1 port map( A1 => n18854, A2 => n25995, B1 => n18790, B2 => 
                           n26757, ZN => n25396);
   U1369 : NAND4_X1 port map( A1 => n25399, A2 => n25398, A3 => n25397, A4 => 
                           n25396, ZN => n25400);
   U1370 : AOI22_X1 port map( A1 => n25780, A2 => n25401, B1 => n25533, B2 => 
                           n25400, ZN => n25402);
   U1371 : OAI21_X1 port map( B1 => n25828, B2 => n25403, A => n25402, ZN => 
                           OUT2(26));
   U1372 : AOI22_X1 port map( A1 => n18324, A2 => n19015, B1 => n25974, B2 => 
                           n19367, ZN => n25407);
   U1373 : AOI22_X1 port map( A1 => n18318, A2 => n19175, B1 => n25985, B2 => 
                           n19303, ZN => n25406);
   U1374 : AOI22_X1 port map( A1 => n18312, A2 => n19047, B1 => n18317, B2 => 
                           n19111, ZN => n25405);
   U1375 : AOI22_X1 port map( A1 => n18310, A2 => n19079, B1 => n18319, B2 => 
                           n19239, ZN => n25404);
   U1376 : NAND4_X1 port map( A1 => n25407, A2 => n25406, A3 => n25405, A4 => 
                           n25404, ZN => n25413);
   U1377 : AOI22_X1 port map( A1 => n18314, A2 => n19143, B1 => n18320, B2 => 
                           n18951, ZN => n25411);
   U1378 : AOI22_X1 port map( A1 => n25903, A2 => n18983, B1 => n25976, B2 => 
                           n19207, ZN => n25410);
   U1379 : AOI22_X1 port map( A1 => n25922, A2 => n18887, B1 => n25923, B2 => 
                           n19335, ZN => n25409);
   U1380 : AOI22_X1 port map( A1 => n25975, A2 => n18919, B1 => n18315, B2 => 
                           n19271, ZN => n25408);
   U1381 : NAND4_X1 port map( A1 => n25411, A2 => n25410, A3 => n25409, A4 => 
                           n25408, ZN => n25412);
   U1382 : NOR2_X1 port map( A1 => n25413, A2 => n25412, ZN => n25425);
   U1383 : AOI22_X1 port map( A1 => n18440, A2 => n19402, B1 => n18504, B2 => 
                           n25939, ZN => n25417);
   U1384 : AOI22_X1 port map( A1 => n18472, A2 => n25866, B1 => n18408, B2 => 
                           n25769, ZN => n25416);
   U1385 : AOI22_X1 port map( A1 => n18536, A2 => n25889, B1 => n18568, B2 => 
                           n26754, ZN => n25415);
   U1386 : AOI22_X1 port map( A1 => n18377, A2 => n19401, B1 => n18600, B2 => 
                           n25995, ZN => n25414);
   U1387 : NAND4_X1 port map( A1 => n25417, A2 => n25416, A3 => n25415, A4 => 
                           n25414, ZN => n25423);
   U1388 : AOI22_X1 port map( A1 => n26001, A2 => n18695, B1 => n18855, B2 => 
                           n26000, ZN => n25421);
   U1389 : AOI22_X1 port map( A1 => n18791, A2 => n25889, B1 => n18823, B2 => 
                           n26754, ZN => n25420);
   U1390 : AOI22_X1 port map( A1 => n18727, A2 => n26756, B1 => n18759, B2 => 
                           n25797, ZN => n25419);
   U1391 : AOI22_X1 port map( A1 => n18631, A2 => n19401, B1 => n18663, B2 => 
                           n25992, ZN => n25418);
   U1392 : NAND4_X1 port map( A1 => n25421, A2 => n25420, A3 => n25419, A4 => 
                           n25418, ZN => n25422);
   U1393 : AOI22_X1 port map( A1 => n25780, A2 => n25423, B1 => n25533, B2 => 
                           n25422, ZN => n25424);
   U1394 : OAI21_X1 port map( B1 => n25828, B2 => n25425, A => n25424, ZN => 
                           OUT2(25));
   U1395 : AOI22_X1 port map( A1 => n25975, A2 => n18920, B1 => n25984, B2 => 
                           n19016, ZN => n25429);
   U1396 : AOI22_X1 port map( A1 => n25922, A2 => n18888, B1 => n18321, B2 => 
                           n19368, ZN => n25428);
   U1397 : AOI22_X1 port map( A1 => n18312, A2 => n19048, B1 => n25923, B2 => 
                           n19336, ZN => n25427);
   U1398 : AOI22_X1 port map( A1 => n18315, A2 => n19272, B1 => n18320, B2 => 
                           n18952, ZN => n25426);
   U1399 : NAND4_X1 port map( A1 => n25429, A2 => n25428, A3 => n25427, A4 => 
                           n25426, ZN => n25435);
   U1400 : AOI22_X1 port map( A1 => n25950, A2 => n19112, B1 => n25976, B2 => 
                           n19208, ZN => n25433);
   U1401 : AOI22_X1 port map( A1 => n18314, A2 => n19144, B1 => n18313, B2 => 
                           n19304, ZN => n25432);
   U1402 : CLKBUF_X1 port map( A => n18318, Z => n25983);
   U1403 : AOI22_X1 port map( A1 => n25983, A2 => n19176, B1 => n25829, B2 => 
                           n19080, ZN => n25431);
   U1404 : AOI22_X1 port map( A1 => n18311, A2 => n18984, B1 => n25981, B2 => 
                           n19240, ZN => n25430);
   U1405 : NAND4_X1 port map( A1 => n25433, A2 => n25432, A3 => n25431, A4 => 
                           n25430, ZN => n25434);
   U1406 : NOR2_X1 port map( A1 => n25435, A2 => n25434, ZN => n25447);
   U1407 : AOI22_X1 port map( A1 => n18288, A2 => n18441, B1 => n18473, B2 => 
                           n25866, ZN => n25439);
   U1408 : AOI22_X1 port map( A1 => n18601, A2 => n26755, B1 => n18505, B2 => 
                           n25797, ZN => n25438);
   U1409 : AOI22_X1 port map( A1 => n19394, A2 => n18291, B1 => n18569, B2 => 
                           n25705, ZN => n25437);
   U1410 : AOI22_X1 port map( A1 => n18409, A2 => n26758, B1 => n18537, B2 => 
                           n25940, ZN => n25436);
   U1411 : NAND4_X1 port map( A1 => n25439, A2 => n25438, A3 => n25437, A4 => 
                           n25436, ZN => n25445);
   U1412 : AOI22_X1 port map( A1 => n18696, A2 => n18288, B1 => n18792, B2 => 
                           n25940, ZN => n25443);
   U1413 : AOI22_X1 port map( A1 => n18632, A2 => n19401, B1 => n18728, B2 => 
                           n25993, ZN => n25442);
   U1414 : AOI22_X1 port map( A1 => n18856, A2 => n25995, B1 => n18760, B2 => 
                           n25797, ZN => n25441);
   U1415 : AOI22_X1 port map( A1 => n18664, A2 => n26758, B1 => n18824, B2 => 
                           n25705, ZN => n25440);
   U1416 : NAND4_X1 port map( A1 => n25443, A2 => n25442, A3 => n25441, A4 => 
                           n25440, ZN => n25444);
   U1417 : AOI22_X1 port map( A1 => n25780, A2 => n25445, B1 => n25533, B2 => 
                           n25444, ZN => n25446);
   U1418 : OAI21_X1 port map( B1 => n25828, B2 => n25447, A => n25446, ZN => 
                           OUT2(24));
   U1419 : AOI22_X1 port map( A1 => n18312, A2 => n19049, B1 => n18309, B2 => 
                           n18921, ZN => n25451);
   U1420 : AOI22_X1 port map( A1 => n18315, A2 => n19273, B1 => n18323, B2 => 
                           n19337, ZN => n25450);
   U1421 : AOI22_X1 port map( A1 => n18317, A2 => n19113, B1 => n25985, B2 => 
                           n19305, ZN => n25449);
   U1422 : AOI22_X1 port map( A1 => n18322, A2 => n19209, B1 => n18320, B2 => 
                           n18953, ZN => n25448);
   U1423 : NAND4_X1 port map( A1 => n25451, A2 => n25450, A3 => n25449, A4 => 
                           n25448, ZN => n25457);
   U1424 : AOI22_X1 port map( A1 => n18321, A2 => n19369, B1 => n25981, B2 => 
                           n19241, ZN => n25455);
   U1425 : AOI22_X1 port map( A1 => n25983, A2 => n19177, B1 => n18314, B2 => 
                           n19145, ZN => n25454);
   U1426 : AOI22_X1 port map( A1 => n25829, A2 => n19081, B1 => n25903, B2 => 
                           n18985, ZN => n25453);
   U1427 : AOI22_X1 port map( A1 => n25922, A2 => n18889, B1 => n25984, B2 => 
                           n19017, ZN => n25452);
   U1428 : NAND4_X1 port map( A1 => n25455, A2 => n25454, A3 => n25453, A4 => 
                           n25452, ZN => n25456);
   U1429 : NOR2_X1 port map( A1 => n25457, A2 => n25456, ZN => n25469);
   U1430 : AOI22_X1 port map( A1 => n18378, A2 => n18291, B1 => n18570, B2 => 
                           n25705, ZN => n25461);
   U1431 : AOI22_X1 port map( A1 => n18442, A2 => n19402, B1 => n18410, B2 => 
                           n25769, ZN => n25460);
   U1432 : AOI22_X1 port map( A1 => n18474, A2 => n25866, B1 => n18538, B2 => 
                           n25889, ZN => n25459);
   U1433 : AOI22_X1 port map( A1 => n18602, A2 => n26755, B1 => n18506, B2 => 
                           n25797, ZN => n25458);
   U1434 : NAND4_X1 port map( A1 => n25461, A2 => n25460, A3 => n25459, A4 => 
                           n25458, ZN => n25467);
   U1435 : AOI22_X1 port map( A1 => n18633, A2 => n25961, B1 => n18857, B2 => 
                           n25995, ZN => n25465);
   U1436 : AOI22_X1 port map( A1 => n18729, A2 => n26756, B1 => n18825, B2 => 
                           n26754, ZN => n25464);
   U1437 : AOI22_X1 port map( A1 => n18665, A2 => n26758, B1 => n18793, B2 => 
                           n25889, ZN => n25463);
   U1438 : AOI22_X1 port map( A1 => n18697, A2 => n19402, B1 => n18761, B2 => 
                           n25797, ZN => n25462);
   U1439 : NAND4_X1 port map( A1 => n25465, A2 => n25464, A3 => n25463, A4 => 
                           n25462, ZN => n25466);
   U1440 : AOI22_X1 port map( A1 => n25780, A2 => n25467, B1 => n25533, B2 => 
                           n25466, ZN => n25468);
   U1441 : OAI21_X1 port map( B1 => n26012, B2 => n25469, A => n25468, ZN => 
                           OUT2(23));
   U1442 : AOI22_X1 port map( A1 => n25983, A2 => n19178, B1 => n25902, B2 => 
                           n18954, ZN => n25473);
   U1443 : AOI22_X1 port map( A1 => n25949, A2 => n19274, B1 => n18317, B2 => 
                           n19114, ZN => n25472);
   U1444 : AOI22_X1 port map( A1 => n18309, A2 => n18922, B1 => n25829, B2 => 
                           n19082, ZN => n25471);
   U1445 : AOI22_X1 port map( A1 => n25928, A2 => n19050, B1 => n18311, B2 => 
                           n18986, ZN => n25470);
   U1446 : NAND4_X1 port map( A1 => n25473, A2 => n25472, A3 => n25471, A4 => 
                           n25470, ZN => n25479);
   U1447 : AOI22_X1 port map( A1 => n18314, A2 => n19146, B1 => n25923, B2 => 
                           n19338, ZN => n25477);
   U1448 : AOI22_X1 port map( A1 => n18321, A2 => n19370, B1 => n18319, B2 => 
                           n19242, ZN => n25476);
   U1449 : AOI22_X1 port map( A1 => n18316, A2 => n18890, B1 => n18313, B2 => 
                           n19306, ZN => n25475);
   U1450 : AOI22_X1 port map( A1 => n25984, A2 => n19018, B1 => n25976, B2 => 
                           n19210, ZN => n25474);
   U1451 : NAND4_X1 port map( A1 => n25477, A2 => n25476, A3 => n25475, A4 => 
                           n25474, ZN => n25478);
   U1452 : NOR2_X1 port map( A1 => n25479, A2 => n25478, ZN => n25491);
   U1453 : AOI22_X1 port map( A1 => n18603, A2 => n26755, B1 => n18507, B2 => 
                           n25797, ZN => n25483);
   U1454 : AOI22_X1 port map( A1 => n18443, A2 => n19402, B1 => n18475, B2 => 
                           n25993, ZN => n25482);
   U1455 : AOI22_X1 port map( A1 => n18379, A2 => n19401, B1 => n18539, B2 => 
                           n25889, ZN => n25481);
   U1456 : AOI22_X1 port map( A1 => n18411, A2 => n26758, B1 => n18571, B2 => 
                           n25705, ZN => n25480);
   U1457 : NAND4_X1 port map( A1 => n25483, A2 => n25482, A3 => n25481, A4 => 
                           n25480, ZN => n25489);
   U1458 : AOI22_X1 port map( A1 => n18826, A2 => n25705, B1 => n18762, B2 => 
                           n25797, ZN => n25487);
   U1459 : AOI22_X1 port map( A1 => n26001, A2 => n18698, B1 => n18730, B2 => 
                           n25993, ZN => n25486);
   U1460 : AOI22_X1 port map( A1 => n18634, A2 => n19401, B1 => n18794, B2 => 
                           n25940, ZN => n25485);
   U1461 : AOI22_X1 port map( A1 => n18666, A2 => n26758, B1 => n18858, B2 => 
                           n26755, ZN => n25484);
   U1462 : NAND4_X1 port map( A1 => n25487, A2 => n25486, A3 => n25485, A4 => 
                           n25484, ZN => n25488);
   U1463 : AOI22_X1 port map( A1 => n25780, A2 => n25489, B1 => n25533, B2 => 
                           n25488, ZN => n25490);
   U1464 : OAI21_X1 port map( B1 => n26012, B2 => n25491, A => n25490, ZN => 
                           OUT2(22));
   U1465 : AOI22_X1 port map( A1 => n25975, A2 => n18923, B1 => n18324, B2 => 
                           n19019, ZN => n25495);
   U1466 : AOI22_X1 port map( A1 => n18321, A2 => n19371, B1 => n18310, B2 => 
                           n19083, ZN => n25494);
   U1467 : AOI22_X1 port map( A1 => n18315, A2 => n19275, B1 => n18317, B2 => 
                           n19115, ZN => n25493);
   U1468 : AOI22_X1 port map( A1 => n18316, A2 => n18891, B1 => n18319, B2 => 
                           n19243, ZN => n25492);
   U1469 : NAND4_X1 port map( A1 => n25495, A2 => n25494, A3 => n25493, A4 => 
                           n25492, ZN => n25501);
   U1470 : AOI22_X1 port map( A1 => n18311, A2 => n18987, B1 => n18313, B2 => 
                           n19307, ZN => n25499);
   U1471 : AOI22_X1 port map( A1 => n25976, A2 => n19211, B1 => n18323, B2 => 
                           n19339, ZN => n25498);
   U1472 : AOI22_X1 port map( A1 => n18318, A2 => n19179, B1 => n18314, B2 => 
                           n19147, ZN => n25497);
   U1473 : AOI22_X1 port map( A1 => n25928, A2 => n19051, B1 => n25902, B2 => 
                           n18955, ZN => n25496);
   U1474 : NAND4_X1 port map( A1 => n25499, A2 => n25498, A3 => n25497, A4 => 
                           n25496, ZN => n25500);
   U1475 : NOR2_X1 port map( A1 => n25501, A2 => n25500, ZN => n25513);
   U1476 : AOI22_X1 port map( A1 => n18476, A2 => n26756, B1 => n18540, B2 => 
                           n25889, ZN => n25505);
   U1477 : AOI22_X1 port map( A1 => n18604, A2 => n26000, B1 => n18572, B2 => 
                           n25705, ZN => n25504);
   U1478 : AOI22_X1 port map( A1 => n18380, A2 => n18291, B1 => n18508, B2 => 
                           n25797, ZN => n25503);
   U1479 : AOI22_X1 port map( A1 => n18288, A2 => n18444, B1 => n18412, B2 => 
                           n25769, ZN => n25502);
   U1480 : NAND4_X1 port map( A1 => n25505, A2 => n25504, A3 => n25503, A4 => 
                           n25502, ZN => n25511);
   U1481 : AOI22_X1 port map( A1 => n18635, A2 => n19401, B1 => n18795, B2 => 
                           n26757, ZN => n25509);
   U1482 : AOI22_X1 port map( A1 => n18827, A2 => n25994, B1 => n18763, B2 => 
                           n25797, ZN => n25508);
   U1483 : AOI22_X1 port map( A1 => n18699, A2 => n19402, B1 => n18731, B2 => 
                           n25993, ZN => n25507);
   U1484 : AOI22_X1 port map( A1 => n18667, A2 => n26758, B1 => n18859, B2 => 
                           n26755, ZN => n25506);
   U1485 : NAND4_X1 port map( A1 => n25509, A2 => n25508, A3 => n25507, A4 => 
                           n25506, ZN => n25510);
   U1486 : AOI22_X1 port map( A1 => n25780, A2 => n25511, B1 => n25533, B2 => 
                           n25510, ZN => n25512);
   U1487 : OAI21_X1 port map( B1 => n26012, B2 => n25513, A => n25512, ZN => 
                           OUT2(21));
   U1488 : AOI22_X1 port map( A1 => n18310, A2 => n19084, B1 => n18320, B2 => 
                           n18956, ZN => n25517);
   U1489 : AOI22_X1 port map( A1 => n18312, A2 => n19052, B1 => n18315, B2 => 
                           n19276, ZN => n25516);
   U1490 : AOI22_X1 port map( A1 => n25982, A2 => n19148, B1 => n18317, B2 => 
                           n19116, ZN => n25515);
   U1491 : AOI22_X1 port map( A1 => n18324, A2 => n19020, B1 => n18311, B2 => 
                           n18988, ZN => n25514);
   U1492 : NAND4_X1 port map( A1 => n25517, A2 => n25516, A3 => n25515, A4 => 
                           n25514, ZN => n25523);
   U1493 : AOI22_X1 port map( A1 => n18309, A2 => n18924, B1 => n18319, B2 => 
                           n19244, ZN => n25521);
   U1494 : AOI22_X1 port map( A1 => n25974, A2 => n19372, B1 => n25923, B2 => 
                           n19340, ZN => n25520);
   U1495 : AOI22_X1 port map( A1 => n18318, A2 => n19180, B1 => n18322, B2 => 
                           n19212, ZN => n25519);
   U1496 : AOI22_X1 port map( A1 => n18316, A2 => n18892, B1 => n18313, B2 => 
                           n19308, ZN => n25518);
   U1497 : NAND4_X1 port map( A1 => n25521, A2 => n25520, A3 => n25519, A4 => 
                           n25518, ZN => n25522);
   U1498 : NOR2_X1 port map( A1 => n25523, A2 => n25522, ZN => n25536);
   U1499 : AOI22_X1 port map( A1 => n25961, A2 => n18381, B1 => n19402, B2 => 
                           n18445, ZN => n25527);
   U1500 : AOI22_X1 port map( A1 => n18477, A2 => n26756, B1 => n18413, B2 => 
                           n25769, ZN => n25526);
   U1501 : AOI22_X1 port map( A1 => n18605, A2 => n26755, B1 => n18541, B2 => 
                           n25940, ZN => n25525);
   U1502 : AOI22_X1 port map( A1 => n18573, A2 => n26754, B1 => n18509, B2 => 
                           n25797, ZN => n25524);
   U1503 : NAND4_X1 port map( A1 => n25527, A2 => n25526, A3 => n25525, A4 => 
                           n25524, ZN => n25534);
   U1504 : AOI22_X1 port map( A1 => n18668, A2 => n26758, B1 => n18828, B2 => 
                           n25705, ZN => n25531);
   U1505 : AOI22_X1 port map( A1 => n26001, A2 => n18700, B1 => n18732, B2 => 
                           n25993, ZN => n25530);
   U1506 : AOI22_X1 port map( A1 => n18796, A2 => n25889, B1 => n18764, B2 => 
                           n25797, ZN => n25529);
   U1507 : AOI22_X1 port map( A1 => n18636, A2 => n19401, B1 => n18860, B2 => 
                           n26755, ZN => n25528);
   U1508 : NAND4_X1 port map( A1 => n25531, A2 => n25530, A3 => n25529, A4 => 
                           n25528, ZN => n25532);
   U1509 : AOI22_X1 port map( A1 => n25780, A2 => n25534, B1 => n25533, B2 => 
                           n25532, ZN => n25535);
   U1510 : OAI21_X1 port map( B1 => n26012, B2 => n25536, A => n25535, ZN => 
                           OUT2(20));
   U1511 : AOI22_X1 port map( A1 => n18312, A2 => n19053, B1 => n18321, B2 => 
                           n19373, ZN => n25540);
   U1512 : AOI22_X1 port map( A1 => n18314, A2 => n19149, B1 => n18323, B2 => 
                           n19341, ZN => n25539);
   U1513 : AOI22_X1 port map( A1 => n25949, A2 => n19277, B1 => n18320, B2 => 
                           n18957, ZN => n25538);
   U1514 : AOI22_X1 port map( A1 => n25975, A2 => n18925, B1 => n25981, B2 => 
                           n19245, ZN => n25537);
   U1515 : NAND4_X1 port map( A1 => n25540, A2 => n25539, A3 => n25538, A4 => 
                           n25537, ZN => n25546);
   U1516 : AOI22_X1 port map( A1 => n18324, A2 => n19021, B1 => n18322, B2 => 
                           n19213, ZN => n25544);
   U1517 : AOI22_X1 port map( A1 => n25950, A2 => n19117, B1 => n25903, B2 => 
                           n18989, ZN => n25543);
   U1518 : AOI22_X1 port map( A1 => n18318, A2 => n19181, B1 => n18310, B2 => 
                           n19085, ZN => n25542);
   U1519 : AOI22_X1 port map( A1 => n25922, A2 => n18893, B1 => n25985, B2 => 
                           n19309, ZN => n25541);
   U1520 : NAND4_X1 port map( A1 => n25544, A2 => n25543, A3 => n25542, A4 => 
                           n25541, ZN => n25545);
   U1521 : NOR2_X1 port map( A1 => n25546, A2 => n25545, ZN => n25558);
   U1522 : AOI22_X1 port map( A1 => n18382, A2 => n25961, B1 => n18574, B2 => 
                           n25705, ZN => n25550);
   U1523 : AOI22_X1 port map( A1 => n18414, A2 => n26758, B1 => n18606, B2 => 
                           n25995, ZN => n25549);
   U1524 : AOI22_X1 port map( A1 => n18542, A2 => n25889, B1 => n18510, B2 => 
                           n26759, ZN => n25548);
   U1525 : AOI22_X1 port map( A1 => n18288, A2 => n18446, B1 => n18478, B2 => 
                           n25866, ZN => n25547);
   U1526 : NAND4_X1 port map( A1 => n25550, A2 => n25549, A3 => n25548, A4 => 
                           n25547, ZN => n25556);
   U1527 : AOI22_X1 port map( A1 => n18669, A2 => n26758, B1 => n18765, B2 => 
                           n26759, ZN => n25554);
   U1528 : AOI22_X1 port map( A1 => n18797, A2 => n25889, B1 => n18829, B2 => 
                           n25705, ZN => n25553);
   U1529 : AOI22_X1 port map( A1 => n18637, A2 => n18291, B1 => n18861, B2 => 
                           n26755, ZN => n25552);
   U1530 : AOI22_X1 port map( A1 => n26001, A2 => n18701, B1 => n18733, B2 => 
                           n25866, ZN => n25551);
   U1531 : NAND4_X1 port map( A1 => n25554, A2 => n25553, A3 => n25552, A4 => 
                           n25551, ZN => n25555);
   U1532 : AOI22_X1 port map( A1 => n25780, A2 => n25556, B1 => n26007, B2 => 
                           n25555, ZN => n25557);
   U1533 : OAI21_X1 port map( B1 => n26012, B2 => n25558, A => n25557, ZN => 
                           OUT2(19));
   U1534 : AOI22_X1 port map( A1 => n18317, A2 => n19118, B1 => n18311, B2 => 
                           n18990, ZN => n25562);
   U1535 : AOI22_X1 port map( A1 => n18309, A2 => n18926, B1 => n18322, B2 => 
                           n19214, ZN => n25561);
   U1536 : AOI22_X1 port map( A1 => n18315, A2 => n19278, B1 => n25985, B2 => 
                           n19310, ZN => n25560);
   U1537 : AOI22_X1 port map( A1 => n18312, A2 => n19054, B1 => n18316, B2 => 
                           n18894, ZN => n25559);
   U1538 : NAND4_X1 port map( A1 => n25562, A2 => n25561, A3 => n25560, A4 => 
                           n25559, ZN => n25568);
   U1539 : AOI22_X1 port map( A1 => n25982, A2 => n19150, B1 => n25902, B2 => 
                           n18958, ZN => n25566);
   U1540 : AOI22_X1 port map( A1 => n18321, A2 => n19374, B1 => n25981, B2 => 
                           n19246, ZN => n25565);
   U1541 : AOI22_X1 port map( A1 => n18324, A2 => n19022, B1 => n25829, B2 => 
                           n19086, ZN => n25564);
   U1542 : AOI22_X1 port map( A1 => n18318, A2 => n19182, B1 => n25923, B2 => 
                           n19342, ZN => n25563);
   U1543 : NAND4_X1 port map( A1 => n25566, A2 => n25565, A3 => n25564, A4 => 
                           n25563, ZN => n25567);
   U1544 : NOR2_X1 port map( A1 => n25568, A2 => n25567, ZN => n25580);
   U1545 : CLKBUF_X1 port map( A => n25734, Z => n26009);
   U1546 : AOI22_X1 port map( A1 => n18479, A2 => n26756, B1 => n18607, B2 => 
                           n26000, ZN => n25572);
   U1547 : AOI22_X1 port map( A1 => n18415, A2 => n26758, B1 => n18511, B2 => 
                           n26759, ZN => n25571);
   U1548 : AOI22_X1 port map( A1 => n18447, A2 => n26001, B1 => n18543, B2 => 
                           n25940, ZN => n25570);
   U1549 : AOI22_X1 port map( A1 => n18383, A2 => n25961, B1 => n18575, B2 => 
                           n25705, ZN => n25569);
   U1550 : NAND4_X1 port map( A1 => n25572, A2 => n25571, A3 => n25570, A4 => 
                           n25569, ZN => n25578);
   U1551 : AOI22_X1 port map( A1 => n18638, A2 => n19401, B1 => n18670, B2 => 
                           n25992, ZN => n25576);
   U1552 : AOI22_X1 port map( A1 => n18830, A2 => n25994, B1 => n18766, B2 => 
                           n26759, ZN => n25575);
   U1553 : AOI22_X1 port map( A1 => n18288, A2 => n18702, B1 => n18862, B2 => 
                           n26755, ZN => n25574);
   U1554 : AOI22_X1 port map( A1 => n18734, A2 => n26756, B1 => n18798, B2 => 
                           n25940, ZN => n25573);
   U1555 : NAND4_X1 port map( A1 => n25576, A2 => n25575, A3 => n25574, A4 => 
                           n25573, ZN => n25577);
   U1556 : AOI22_X1 port map( A1 => n26009, A2 => n25578, B1 => n26007, B2 => 
                           n25577, ZN => n25579);
   U1557 : OAI21_X1 port map( B1 => n26012, B2 => n25580, A => n25579, ZN => 
                           OUT2(18));
   U1558 : AOI22_X1 port map( A1 => n25949, A2 => n19279, B1 => n18323, B2 => 
                           n19343, ZN => n25584);
   U1559 : AOI22_X1 port map( A1 => n25928, A2 => n19055, B1 => n25983, B2 => 
                           n19183, ZN => n25583);
   U1560 : AOI22_X1 port map( A1 => n18324, A2 => n19023, B1 => n18310, B2 => 
                           n19087, ZN => n25582);
   U1561 : AOI22_X1 port map( A1 => n18309, A2 => n18927, B1 => n18321, B2 => 
                           n19375, ZN => n25581);
   U1562 : NAND4_X1 port map( A1 => n25584, A2 => n25583, A3 => n25582, A4 => 
                           n25581, ZN => n25590);
   U1563 : AOI22_X1 port map( A1 => n18311, A2 => n18991, B1 => n18322, B2 => 
                           n19215, ZN => n25588);
   U1564 : AOI22_X1 port map( A1 => n18314, A2 => n19151, B1 => n18319, B2 => 
                           n19247, ZN => n25587);
   U1565 : AOI22_X1 port map( A1 => n18316, A2 => n18895, B1 => n25902, B2 => 
                           n18959, ZN => n25586);
   U1566 : AOI22_X1 port map( A1 => n25950, A2 => n19119, B1 => n18313, B2 => 
                           n19311, ZN => n25585);
   U1567 : NAND4_X1 port map( A1 => n25588, A2 => n25587, A3 => n25586, A4 => 
                           n25585, ZN => n25589);
   U1568 : NOR2_X1 port map( A1 => n25590, A2 => n25589, ZN => n25602);
   U1569 : AOI22_X1 port map( A1 => n19393, A2 => n25995, B1 => n18544, B2 => 
                           n25940, ZN => n25594);
   U1570 : AOI22_X1 port map( A1 => n25961, A2 => n18384, B1 => n18416, B2 => 
                           n25769, ZN => n25593);
   U1571 : AOI22_X1 port map( A1 => n18576, A2 => n25994, B1 => n18512, B2 => 
                           n26759, ZN => n25592);
   U1572 : AOI22_X1 port map( A1 => n18288, A2 => n18448, B1 => n18480, B2 => 
                           n25866, ZN => n25591);
   U1573 : NAND4_X1 port map( A1 => n25594, A2 => n25593, A3 => n25592, A4 => 
                           n25591, ZN => n25600);
   U1574 : AOI22_X1 port map( A1 => n18735, A2 => n26756, B1 => n18767, B2 => 
                           n26759, ZN => n25598);
   U1575 : AOI22_X1 port map( A1 => n18671, A2 => n26758, B1 => n18831, B2 => 
                           n25705, ZN => n25597);
   U1576 : AOI22_X1 port map( A1 => n26001, A2 => n18703, B1 => n18863, B2 => 
                           n26755, ZN => n25596);
   U1577 : AOI22_X1 port map( A1 => n18639, A2 => n25961, B1 => n18799, B2 => 
                           n25940, ZN => n25595);
   U1578 : NAND4_X1 port map( A1 => n25598, A2 => n25597, A3 => n25596, A4 => 
                           n25595, ZN => n25599);
   U1579 : AOI22_X1 port map( A1 => n26009, A2 => n25600, B1 => n26007, B2 => 
                           n25599, ZN => n25601);
   U1580 : OAI21_X1 port map( B1 => n26012, B2 => n25602, A => n25601, ZN => 
                           OUT2(17));
   U1581 : AOI22_X1 port map( A1 => n18318, A2 => n19184, B1 => n25950, B2 => 
                           n19120, ZN => n25606);
   U1582 : AOI22_X1 port map( A1 => n25982, A2 => n19152, B1 => n18322, B2 => 
                           n19216, ZN => n25605);
   U1583 : AOI22_X1 port map( A1 => n18309, A2 => n18928, B1 => n25829, B2 => 
                           n19088, ZN => n25604);
   U1584 : AOI22_X1 port map( A1 => n18312, A2 => n19056, B1 => n18324, B2 => 
                           n19024, ZN => n25603);
   U1585 : NAND4_X1 port map( A1 => n25606, A2 => n25605, A3 => n25604, A4 => 
                           n25603, ZN => n25612);
   U1586 : AOI22_X1 port map( A1 => n18320, A2 => n18960, B1 => n18319, B2 => 
                           n19248, ZN => n25610);
   U1587 : AOI22_X1 port map( A1 => n18316, A2 => n18896, B1 => n18323, B2 => 
                           n19344, ZN => n25609);
   U1588 : AOI22_X1 port map( A1 => n18315, A2 => n19280, B1 => n18311, B2 => 
                           n18992, ZN => n25608);
   U1589 : AOI22_X1 port map( A1 => n25974, A2 => n19376, B1 => n25985, B2 => 
                           n19312, ZN => n25607);
   U1590 : NAND4_X1 port map( A1 => n25610, A2 => n25609, A3 => n25608, A4 => 
                           n25607, ZN => n25611);
   U1591 : NOR2_X1 port map( A1 => n25612, A2 => n25611, ZN => n25624);
   U1592 : AOI22_X1 port map( A1 => n18449, A2 => n19402, B1 => n18577, B2 => 
                           n25705, ZN => n25616);
   U1593 : AOI22_X1 port map( A1 => n18608, A2 => n26755, B1 => n18513, B2 => 
                           n26759, ZN => n25615);
   U1594 : AOI22_X1 port map( A1 => n18481, A2 => n26756, B1 => n18545, B2 => 
                           n25940, ZN => n25614);
   U1595 : AOI22_X1 port map( A1 => n18291, A2 => n18385, B1 => n18417, B2 => 
                           n25992, ZN => n25613);
   U1596 : NAND4_X1 port map( A1 => n25616, A2 => n25615, A3 => n25614, A4 => 
                           n25613, ZN => n25622);
   U1597 : AOI22_X1 port map( A1 => n18640, A2 => n19401, B1 => n18864, B2 => 
                           n26755, ZN => n25620);
   U1598 : AOI22_X1 port map( A1 => n18800, A2 => n26757, B1 => n18768, B2 => 
                           n26759, ZN => n25619);
   U1599 : AOI22_X1 port map( A1 => n18736, A2 => n26756, B1 => n18832, B2 => 
                           n25705, ZN => n25618);
   U1600 : AOI22_X1 port map( A1 => n18288, A2 => n18704, B1 => n18672, B2 => 
                           n25992, ZN => n25617);
   U1601 : NAND4_X1 port map( A1 => n25620, A2 => n25619, A3 => n25618, A4 => 
                           n25617, ZN => n25621);
   U1602 : AOI22_X1 port map( A1 => n25780, A2 => n25622, B1 => n26007, B2 => 
                           n25621, ZN => n25623);
   U1603 : OAI21_X1 port map( B1 => n26012, B2 => n25624, A => n25623, ZN => 
                           OUT2(16));
   U1604 : AOI22_X1 port map( A1 => n25922, A2 => n18897, B1 => n18309, B2 => 
                           n18929, ZN => n25628);
   U1605 : AOI22_X1 port map( A1 => n18310, A2 => n19089, B1 => n18313, B2 => 
                           n19313, ZN => n25627);
   U1606 : AOI22_X1 port map( A1 => n18314, A2 => n19153, B1 => n18320, B2 => 
                           n18961, ZN => n25626);
   U1607 : AOI22_X1 port map( A1 => n18315, A2 => n19281, B1 => n25923, B2 => 
                           n19345, ZN => n25625);
   U1608 : NAND4_X1 port map( A1 => n25628, A2 => n25627, A3 => n25626, A4 => 
                           n25625, ZN => n25634);
   U1609 : AOI22_X1 port map( A1 => n18312, A2 => n19057, B1 => n18324, B2 => 
                           n19025, ZN => n25632);
   U1610 : AOI22_X1 port map( A1 => n18321, A2 => n19377, B1 => n25981, B2 => 
                           n19249, ZN => n25631);
   U1611 : AOI22_X1 port map( A1 => n18318, A2 => n19185, B1 => n25950, B2 => 
                           n19121, ZN => n25630);
   U1612 : AOI22_X1 port map( A1 => n18311, A2 => n18993, B1 => n25976, B2 => 
                           n19217, ZN => n25629);
   U1613 : NAND4_X1 port map( A1 => n25632, A2 => n25631, A3 => n25630, A4 => 
                           n25629, ZN => n25633);
   U1614 : NOR2_X1 port map( A1 => n25634, A2 => n25633, ZN => n25646);
   U1615 : AOI22_X1 port map( A1 => n18450, A2 => n26001, B1 => n18514, B2 => 
                           n26759, ZN => n25638);
   U1616 : AOI22_X1 port map( A1 => n18482, A2 => n25993, B1 => n18418, B2 => 
                           n25769, ZN => n25637);
   U1617 : AOI22_X1 port map( A1 => n18609, A2 => n26755, B1 => n18546, B2 => 
                           n25940, ZN => n25636);
   U1618 : AOI22_X1 port map( A1 => n18386, A2 => n18291, B1 => n18578, B2 => 
                           n25705, ZN => n25635);
   U1619 : NAND4_X1 port map( A1 => n25638, A2 => n25637, A3 => n25636, A4 => 
                           n25635, ZN => n25644);
   U1620 : AOI22_X1 port map( A1 => n18737, A2 => n26756, B1 => n18833, B2 => 
                           n25705, ZN => n25642);
   U1621 : AOI22_X1 port map( A1 => n18673, A2 => n26758, B1 => n18769, B2 => 
                           n26759, ZN => n25641);
   U1622 : AOI22_X1 port map( A1 => n26001, A2 => n18705, B1 => n18865, B2 => 
                           n26000, ZN => n25640);
   U1623 : AOI22_X1 port map( A1 => n18641, A2 => n18291, B1 => n18801, B2 => 
                           n25940, ZN => n25639);
   U1624 : NAND4_X1 port map( A1 => n25642, A2 => n25641, A3 => n25640, A4 => 
                           n25639, ZN => n25643);
   U1625 : AOI22_X1 port map( A1 => n25780, A2 => n25644, B1 => n26007, B2 => 
                           n25643, ZN => n25645);
   U1626 : OAI21_X1 port map( B1 => n26012, B2 => n25646, A => n25645, ZN => 
                           OUT2(15));
   U1627 : AOI22_X1 port map( A1 => n25922, A2 => n18898, B1 => n18311, B2 => 
                           n18994, ZN => n25650);
   U1628 : AOI22_X1 port map( A1 => n18309, A2 => n18930, B1 => n25950, B2 => 
                           n19122, ZN => n25649);
   U1629 : AOI22_X1 port map( A1 => n18312, A2 => n19058, B1 => n25949, B2 => 
                           n19282, ZN => n25648);
   U1630 : AOI22_X1 port map( A1 => n25983, A2 => n19186, B1 => n25974, B2 => 
                           n19378, ZN => n25647);
   U1631 : NAND4_X1 port map( A1 => n25650, A2 => n25649, A3 => n25648, A4 => 
                           n25647, ZN => n25656);
   U1632 : AOI22_X1 port map( A1 => n18322, A2 => n19218, B1 => n18323, B2 => 
                           n19346, ZN => n25654);
   U1633 : AOI22_X1 port map( A1 => n18313, A2 => n19314, B1 => n18320, B2 => 
                           n18962, ZN => n25653);
   U1634 : AOI22_X1 port map( A1 => n25984, A2 => n19026, B1 => n25982, B2 => 
                           n19154, ZN => n25652);
   U1635 : AOI22_X1 port map( A1 => n18310, A2 => n19090, B1 => n25981, B2 => 
                           n19250, ZN => n25651);
   U1636 : NAND4_X1 port map( A1 => n25654, A2 => n25653, A3 => n25652, A4 => 
                           n25651, ZN => n25655);
   U1637 : NOR2_X1 port map( A1 => n25656, A2 => n25655, ZN => n25668);
   U1638 : AOI22_X1 port map( A1 => n18579, A2 => n26754, B1 => n18515, B2 => 
                           n26759, ZN => n25660);
   U1639 : AOI22_X1 port map( A1 => n18451, A2 => n26001, B1 => n18547, B2 => 
                           n25889, ZN => n25659);
   U1640 : AOI22_X1 port map( A1 => n18483, A2 => n26756, B1 => n18610, B2 => 
                           n26000, ZN => n25658);
   U1641 : AOI22_X1 port map( A1 => n18291, A2 => n18387, B1 => n18419, B2 => 
                           n25769, ZN => n25657);
   U1642 : NAND4_X1 port map( A1 => n25660, A2 => n25659, A3 => n25658, A4 => 
                           n25657, ZN => n25666);
   U1643 : AOI22_X1 port map( A1 => n18674, A2 => n26758, B1 => n18834, B2 => 
                           n25705, ZN => n25664);
   U1644 : AOI22_X1 port map( A1 => n18706, A2 => n18288, B1 => n18770, B2 => 
                           n26759, ZN => n25663);
   U1645 : AOI22_X1 port map( A1 => n18738, A2 => n26756, B1 => n18866, B2 => 
                           n26000, ZN => n25662);
   U1646 : AOI22_X1 port map( A1 => n18642, A2 => n19401, B1 => n18802, B2 => 
                           n26757, ZN => n25661);
   U1647 : NAND4_X1 port map( A1 => n25664, A2 => n25663, A3 => n25662, A4 => 
                           n25661, ZN => n25665);
   U1648 : AOI22_X1 port map( A1 => n25780, A2 => n25666, B1 => n26007, B2 => 
                           n25665, ZN => n25667);
   U1649 : OAI21_X1 port map( B1 => n26012, B2 => n25668, A => n25667, ZN => 
                           OUT2(14));
   U1650 : AOI22_X1 port map( A1 => n25922, A2 => n18899, B1 => n18310, B2 => 
                           n19091, ZN => n25672);
   U1651 : AOI22_X1 port map( A1 => n18317, A2 => n19123, B1 => n25903, B2 => 
                           n18995, ZN => n25671);
   U1652 : AOI22_X1 port map( A1 => n18324, A2 => n19027, B1 => n18319, B2 => 
                           n19251, ZN => n25670);
   U1653 : AOI22_X1 port map( A1 => n18314, A2 => n19155, B1 => n25976, B2 => 
                           n19219, ZN => n25669);
   U1654 : NAND4_X1 port map( A1 => n25672, A2 => n25671, A3 => n25670, A4 => 
                           n25669, ZN => n25678);
   U1655 : AOI22_X1 port map( A1 => n25975, A2 => n18931, B1 => n25985, B2 => 
                           n19315, ZN => n25676);
   U1656 : AOI22_X1 port map( A1 => n25928, A2 => n19059, B1 => n25949, B2 => 
                           n19283, ZN => n25675);
   U1657 : AOI22_X1 port map( A1 => n25983, A2 => n19187, B1 => n25974, B2 => 
                           n19379, ZN => n25674);
   U1658 : AOI22_X1 port map( A1 => n25902, A2 => n18963, B1 => n25923, B2 => 
                           n19347, ZN => n25673);
   U1659 : NAND4_X1 port map( A1 => n25676, A2 => n25675, A3 => n25674, A4 => 
                           n25673, ZN => n25677);
   U1660 : NOR2_X1 port map( A1 => n25678, A2 => n25677, ZN => n25690);
   U1661 : AOI22_X1 port map( A1 => n18288, A2 => n18452, B1 => n18291, B2 => 
                           n18388, ZN => n25682);
   U1662 : AOI22_X1 port map( A1 => n18548, A2 => n26757, B1 => n18580, B2 => 
                           n26754, ZN => n25681);
   U1663 : AOI22_X1 port map( A1 => n18420, A2 => n26758, B1 => n18516, B2 => 
                           n25797, ZN => n25680);
   U1664 : AOI22_X1 port map( A1 => n18484, A2 => n25993, B1 => n18611, B2 => 
                           n26000, ZN => n25679);
   U1665 : NAND4_X1 port map( A1 => n25682, A2 => n25681, A3 => n25680, A4 => 
                           n25679, ZN => n25688);
   U1666 : AOI22_X1 port map( A1 => n18803, A2 => n26757, B1 => n18771, B2 => 
                           n25797, ZN => n25686);
   U1667 : AOI22_X1 port map( A1 => n18643, A2 => n18291, B1 => n18835, B2 => 
                           n25705, ZN => n25685);
   U1668 : AOI22_X1 port map( A1 => n26001, A2 => n18707, B1 => n18739, B2 => 
                           n25866, ZN => n25684);
   U1669 : AOI22_X1 port map( A1 => n18675, A2 => n26758, B1 => n18867, B2 => 
                           n26000, ZN => n25683);
   U1670 : NAND4_X1 port map( A1 => n25686, A2 => n25685, A3 => n25684, A4 => 
                           n25683, ZN => n25687);
   U1671 : AOI22_X1 port map( A1 => n25780, A2 => n25688, B1 => n26007, B2 => 
                           n25687, ZN => n25689);
   U1672 : OAI21_X1 port map( B1 => n26012, B2 => n25690, A => n25689, ZN => 
                           OUT2(13));
   U1673 : AOI22_X1 port map( A1 => n18315, A2 => n19284, B1 => n18317, B2 => 
                           n19124, ZN => n25694);
   U1674 : AOI22_X1 port map( A1 => n18309, A2 => n18932, B1 => n18323, B2 => 
                           n19348, ZN => n25693);
   U1675 : AOI22_X1 port map( A1 => n25928, A2 => n19060, B1 => n18316, B2 => 
                           n18900, ZN => n25692);
   U1676 : AOI22_X1 port map( A1 => n25829, A2 => n19092, B1 => n18314, B2 => 
                           n19156, ZN => n25691);
   U1677 : NAND4_X1 port map( A1 => n25694, A2 => n25693, A3 => n25692, A4 => 
                           n25691, ZN => n25700);
   U1678 : AOI22_X1 port map( A1 => n25983, A2 => n19188, B1 => n25984, B2 => 
                           n19028, ZN => n25698);
   U1679 : AOI22_X1 port map( A1 => n18322, A2 => n19220, B1 => n18313, B2 => 
                           n19316, ZN => n25697);
   U1680 : AOI22_X1 port map( A1 => n25974, A2 => n19380, B1 => n25903, B2 => 
                           n18996, ZN => n25696);
   U1681 : AOI22_X1 port map( A1 => n18320, A2 => n18964, B1 => n18319, B2 => 
                           n19252, ZN => n25695);
   U1682 : NAND4_X1 port map( A1 => n25698, A2 => n25697, A3 => n25696, A4 => 
                           n25695, ZN => n25699);
   U1683 : NOR2_X1 port map( A1 => n25700, A2 => n25699, ZN => n25713);
   U1684 : AOI22_X1 port map( A1 => n18389, A2 => n25961, B1 => n18581, B2 => 
                           n26754, ZN => n25704);
   U1685 : AOI22_X1 port map( A1 => n18549, A2 => n26757, B1 => n18517, B2 => 
                           n25797, ZN => n25703);
   U1686 : AOI22_X1 port map( A1 => n18485, A2 => n26756, B1 => n18421, B2 => 
                           n25769, ZN => n25702);
   U1687 : AOI22_X1 port map( A1 => n18288, A2 => n18453, B1 => n18612, B2 => 
                           n26000, ZN => n25701);
   U1688 : NAND4_X1 port map( A1 => n25704, A2 => n25703, A3 => n25702, A4 => 
                           n25701, ZN => n25711);
   U1689 : AOI22_X1 port map( A1 => n18291, A2 => n18644, B1 => n18740, B2 => 
                           n25993, ZN => n25709);
   U1690 : AOI22_X1 port map( A1 => n18708, A2 => n18288, B1 => n18772, B2 => 
                           n25797, ZN => n25708);
   U1691 : AOI22_X1 port map( A1 => n18868, A2 => n25995, B1 => n18836, B2 => 
                           n25705, ZN => n25707);
   U1692 : AOI22_X1 port map( A1 => n18676, A2 => n26758, B1 => n18804, B2 => 
                           n26757, ZN => n25706);
   U1693 : NAND4_X1 port map( A1 => n25709, A2 => n25708, A3 => n25707, A4 => 
                           n25706, ZN => n25710);
   U1694 : AOI22_X1 port map( A1 => n25780, A2 => n25711, B1 => n26007, B2 => 
                           n25710, ZN => n25712);
   U1695 : OAI21_X1 port map( B1 => n26012, B2 => n25713, A => n25712, ZN => 
                           OUT2(12));
   U1696 : AOI22_X1 port map( A1 => n25829, A2 => n19093, B1 => n18314, B2 => 
                           n19157, ZN => n25717);
   U1697 : AOI22_X1 port map( A1 => n25975, A2 => n18933, B1 => n25984, B2 => 
                           n19029, ZN => n25716);
   U1698 : AOI22_X1 port map( A1 => n18320, A2 => n18965, B1 => n25923, B2 => 
                           n19349, ZN => n25715);
   U1699 : AOI22_X1 port map( A1 => n18311, A2 => n18997, B1 => n18319, B2 => 
                           n19253, ZN => n25714);
   U1700 : NAND4_X1 port map( A1 => n25717, A2 => n25716, A3 => n25715, A4 => 
                           n25714, ZN => n25723);
   U1701 : AOI22_X1 port map( A1 => n18315, A2 => n19285, B1 => n25976, B2 => 
                           n19221, ZN => n25721);
   U1702 : AOI22_X1 port map( A1 => n18312, A2 => n19061, B1 => n18317, B2 => 
                           n19125, ZN => n25720);
   U1703 : AOI22_X1 port map( A1 => n18316, A2 => n18901, B1 => n18321, B2 => 
                           n19381, ZN => n25719);
   U1704 : AOI22_X1 port map( A1 => n18318, A2 => n19189, B1 => n18313, B2 => 
                           n19317, ZN => n25718);
   U1705 : NAND4_X1 port map( A1 => n25721, A2 => n25720, A3 => n25719, A4 => 
                           n25718, ZN => n25722);
   U1706 : NOR2_X1 port map( A1 => n25723, A2 => n25722, ZN => n25736);
   U1707 : AOI22_X1 port map( A1 => n18613, A2 => n26755, B1 => n18518, B2 => 
                           n25797, ZN => n25727);
   U1708 : AOI22_X1 port map( A1 => n18390, A2 => n19401, B1 => n18582, B2 => 
                           n26754, ZN => n25726);
   U1709 : AOI22_X1 port map( A1 => n18288, A2 => n18454, B1 => n18486, B2 => 
                           n25866, ZN => n25725);
   U1710 : AOI22_X1 port map( A1 => n18422, A2 => n26758, B1 => n18550, B2 => 
                           n26757, ZN => n25724);
   U1711 : NAND4_X1 port map( A1 => n25727, A2 => n25726, A3 => n25725, A4 => 
                           n25724, ZN => n25733);
   U1712 : AOI22_X1 port map( A1 => n18741, A2 => n26756, B1 => n18773, B2 => 
                           n25797, ZN => n25731);
   U1713 : AOI22_X1 port map( A1 => n18869, A2 => n25995, B1 => n18837, B2 => 
                           n26754, ZN => n25730);
   U1714 : AOI22_X1 port map( A1 => n25961, A2 => n18645, B1 => n18677, B2 => 
                           n25769, ZN => n25729);
   U1715 : AOI22_X1 port map( A1 => n18709, A2 => n18288, B1 => n18805, B2 => 
                           n26757, ZN => n25728);
   U1716 : NAND4_X1 port map( A1 => n25731, A2 => n25730, A3 => n25729, A4 => 
                           n25728, ZN => n25732);
   U1717 : AOI22_X1 port map( A1 => n25734, A2 => n25733, B1 => n26007, B2 => 
                           n25732, ZN => n25735);
   U1718 : OAI21_X1 port map( B1 => n25828, B2 => n25736, A => n25735, ZN => 
                           OUT2(11));
   U1719 : AOI22_X1 port map( A1 => n18318, A2 => n19190, B1 => n18313, B2 => 
                           n19318, ZN => n25740);
   U1720 : AOI22_X1 port map( A1 => n25949, A2 => n19286, B1 => n25903, B2 => 
                           n18998, ZN => n25739);
   U1721 : AOI22_X1 port map( A1 => n18319, A2 => n19254, B1 => n18323, B2 => 
                           n19350, ZN => n25738);
   U1722 : AOI22_X1 port map( A1 => n18317, A2 => n19126, B1 => n18320, B2 => 
                           n18966, ZN => n25737);
   U1723 : NAND4_X1 port map( A1 => n25740, A2 => n25739, A3 => n25738, A4 => 
                           n25737, ZN => n25746);
   U1724 : AOI22_X1 port map( A1 => n18310, A2 => n19094, B1 => n25976, B2 => 
                           n19222, ZN => n25744);
   U1725 : AOI22_X1 port map( A1 => n18309, A2 => n18934, B1 => n18324, B2 => 
                           n19030, ZN => n25743);
   U1726 : AOI22_X1 port map( A1 => n18316, A2 => n18902, B1 => n25974, B2 => 
                           n19382, ZN => n25742);
   U1727 : AOI22_X1 port map( A1 => n25928, A2 => n19062, B1 => n18314, B2 => 
                           n19158, ZN => n25741);
   U1728 : NAND4_X1 port map( A1 => n25744, A2 => n25743, A3 => n25742, A4 => 
                           n25741, ZN => n25745);
   U1729 : NOR2_X1 port map( A1 => n25746, A2 => n25745, ZN => n25758);
   U1730 : AOI22_X1 port map( A1 => n26001, A2 => n18455, B1 => n18487, B2 => 
                           n25866, ZN => n25750);
   U1731 : AOI22_X1 port map( A1 => n18551, A2 => n26757, B1 => n18519, B2 => 
                           n25797, ZN => n25749);
   U1732 : AOI22_X1 port map( A1 => n18391, A2 => n19401, B1 => n18583, B2 => 
                           n26754, ZN => n25748);
   U1733 : AOI22_X1 port map( A1 => n18423, A2 => n26758, B1 => n18614, B2 => 
                           n26000, ZN => n25747);
   U1734 : NAND4_X1 port map( A1 => n25750, A2 => n25749, A3 => n25748, A4 => 
                           n25747, ZN => n25756);
   U1735 : AOI22_X1 port map( A1 => n18710, A2 => n26001, B1 => n18838, B2 => 
                           n26754, ZN => n25754);
   U1736 : AOI22_X1 port map( A1 => n18678, A2 => n25769, B1 => n18806, B2 => 
                           n26757, ZN => n25753);
   U1737 : AOI22_X1 port map( A1 => n18742, A2 => n26756, B1 => n18774, B2 => 
                           n25797, ZN => n25752);
   U1738 : AOI22_X1 port map( A1 => n18646, A2 => n25961, B1 => n18870, B2 => 
                           n26000, ZN => n25751);
   U1739 : NAND4_X1 port map( A1 => n25754, A2 => n25753, A3 => n25752, A4 => 
                           n25751, ZN => n25755);
   U1740 : AOI22_X1 port map( A1 => n25780, A2 => n25756, B1 => n26007, B2 => 
                           n25755, ZN => n25757);
   U1741 : OAI21_X1 port map( B1 => n25828, B2 => n25758, A => n25757, ZN => 
                           OUT2(10));
   U1742 : AOI22_X1 port map( A1 => n18315, A2 => n19287, B1 => n18321, B2 => 
                           n19383, ZN => n25762);
   U1743 : AOI22_X1 port map( A1 => n25975, A2 => n18935, B1 => n18313, B2 => 
                           n19319, ZN => n25761);
   U1744 : AOI22_X1 port map( A1 => n25984, A2 => n19031, B1 => n25950, B2 => 
                           n19127, ZN => n25760);
   U1745 : AOI22_X1 port map( A1 => n18322, A2 => n19223, B1 => n25902, B2 => 
                           n18967, ZN => n25759);
   U1746 : NAND4_X1 port map( A1 => n25762, A2 => n25761, A3 => n25760, A4 => 
                           n25759, ZN => n25768);
   U1747 : AOI22_X1 port map( A1 => n18312, A2 => n19063, B1 => n25922, B2 => 
                           n18903, ZN => n25766);
   U1748 : AOI22_X1 port map( A1 => n18310, A2 => n19095, B1 => n18323, B2 => 
                           n19351, ZN => n25765);
   U1749 : AOI22_X1 port map( A1 => n18318, A2 => n19191, B1 => n25981, B2 => 
                           n19255, ZN => n25764);
   U1750 : AOI22_X1 port map( A1 => n18314, A2 => n19159, B1 => n18311, B2 => 
                           n18999, ZN => n25763);
   U1751 : NAND4_X1 port map( A1 => n25766, A2 => n25765, A3 => n25764, A4 => 
                           n25763, ZN => n25767);
   U1752 : NOR2_X1 port map( A1 => n25768, A2 => n25767, ZN => n25782);
   U1753 : AOI22_X1 port map( A1 => n18615, A2 => n25995, B1 => n18520, B2 => 
                           n25797, ZN => n25773);
   U1754 : AOI22_X1 port map( A1 => n18488, A2 => n25993, B1 => n18424, B2 => 
                           n25769, ZN => n25772);
   U1755 : AOI22_X1 port map( A1 => n18288, A2 => n18456, B1 => n19401, B2 => 
                           n18392, ZN => n25771);
   U1756 : AOI22_X1 port map( A1 => n18552, A2 => n26757, B1 => n18584, B2 => 
                           n26754, ZN => n25770);
   U1757 : NAND4_X1 port map( A1 => n25773, A2 => n25772, A3 => n25771, A4 => 
                           n25770, ZN => n25779);
   U1758 : AOI22_X1 port map( A1 => n18743, A2 => n26756, B1 => n18871, B2 => 
                           n26000, ZN => n25777);
   U1759 : AOI22_X1 port map( A1 => n26001, A2 => n18711, B1 => n18679, B2 => 
                           n25992, ZN => n25776);
   U1760 : AOI22_X1 port map( A1 => n18807, A2 => n26757, B1 => n18775, B2 => 
                           n25797, ZN => n25775);
   U1761 : AOI22_X1 port map( A1 => n18647, A2 => n18291, B1 => n18839, B2 => 
                           n25994, ZN => n25774);
   U1762 : NAND4_X1 port map( A1 => n25777, A2 => n25776, A3 => n25775, A4 => 
                           n25774, ZN => n25778);
   U1763 : AOI22_X1 port map( A1 => n25780, A2 => n25779, B1 => n26007, B2 => 
                           n25778, ZN => n25781);
   U1764 : OAI21_X1 port map( B1 => n25828, B2 => n25782, A => n25781, ZN => 
                           OUT2(9));
   U1765 : AOI22_X1 port map( A1 => n18314, A2 => n19160, B1 => n18322, B2 => 
                           n19224, ZN => n25786);
   U1766 : AOI22_X1 port map( A1 => n18310, A2 => n19096, B1 => n18317, B2 => 
                           n19128, ZN => n25785);
   U1767 : AOI22_X1 port map( A1 => n18316, A2 => n18904, B1 => n18315, B2 => 
                           n19288, ZN => n25784);
   U1768 : AOI22_X1 port map( A1 => n18309, A2 => n18936, B1 => n25985, B2 => 
                           n19320, ZN => n25783);
   U1769 : NAND4_X1 port map( A1 => n25786, A2 => n25785, A3 => n25784, A4 => 
                           n25783, ZN => n25792);
   U1770 : AOI22_X1 port map( A1 => n18318, A2 => n19192, B1 => n18323, B2 => 
                           n19352, ZN => n25790);
   U1771 : AOI22_X1 port map( A1 => n25928, A2 => n19064, B1 => n18324, B2 => 
                           n19032, ZN => n25789);
   U1772 : AOI22_X1 port map( A1 => n18311, A2 => n19000, B1 => n25981, B2 => 
                           n19256, ZN => n25788);
   U1773 : AOI22_X1 port map( A1 => n18321, A2 => n19384, B1 => n25902, B2 => 
                           n18968, ZN => n25787);
   U1774 : NAND4_X1 port map( A1 => n25790, A2 => n25789, A3 => n25788, A4 => 
                           n25787, ZN => n25791);
   U1775 : NOR2_X1 port map( A1 => n25792, A2 => n25791, ZN => n25805);
   U1776 : AOI22_X1 port map( A1 => n18425, A2 => n25992, B1 => n18616, B2 => 
                           n26000, ZN => n25796);
   U1777 : AOI22_X1 port map( A1 => n18457, A2 => n18288, B1 => n18553, B2 => 
                           n25940, ZN => n25795);
   U1778 : AOI22_X1 port map( A1 => n18393, A2 => n18291, B1 => n18521, B2 => 
                           n25797, ZN => n25794);
   U1779 : AOI22_X1 port map( A1 => n18489, A2 => n25993, B1 => n18585, B2 => 
                           n25994, ZN => n25793);
   U1780 : NAND4_X1 port map( A1 => n25796, A2 => n25795, A3 => n25794, A4 => 
                           n25793, ZN => n25803);
   U1781 : AOI22_X1 port map( A1 => n18680, A2 => n25992, B1 => n18840, B2 => 
                           n25994, ZN => n25801);
   U1782 : AOI22_X1 port map( A1 => n18744, A2 => n25993, B1 => n18808, B2 => 
                           n26757, ZN => n25800);
   U1783 : AOI22_X1 port map( A1 => n18712, A2 => n19402, B1 => n18776, B2 => 
                           n25797, ZN => n25799);
   U1784 : AOI22_X1 port map( A1 => n18648, A2 => n19401, B1 => n18872, B2 => 
                           n25995, ZN => n25798);
   U1785 : NAND4_X1 port map( A1 => n25801, A2 => n25800, A3 => n25799, A4 => 
                           n25798, ZN => n25802);
   U1786 : AOI22_X1 port map( A1 => n26009, A2 => n25803, B1 => n26007, B2 => 
                           n25802, ZN => n25804);
   U1787 : OAI21_X1 port map( B1 => n25828, B2 => n25805, A => n25804, ZN => 
                           OUT2(8));
   U1788 : AOI22_X1 port map( A1 => n25982, A2 => n19161, B1 => n18323, B2 => 
                           n19353, ZN => n25809);
   U1789 : AOI22_X1 port map( A1 => n18324, A2 => n19033, B1 => n18313, B2 => 
                           n19321, ZN => n25808);
   U1790 : AOI22_X1 port map( A1 => n25903, A2 => n19001, B1 => n18322, B2 => 
                           n19225, ZN => n25807);
   U1791 : AOI22_X1 port map( A1 => n18316, A2 => n18905, B1 => n18317, B2 => 
                           n19129, ZN => n25806);
   U1792 : NAND4_X1 port map( A1 => n25809, A2 => n25808, A3 => n25807, A4 => 
                           n25806, ZN => n25815);
   U1793 : AOI22_X1 port map( A1 => n25949, A2 => n19289, B1 => n25974, B2 => 
                           n19385, ZN => n25813);
   U1794 : AOI22_X1 port map( A1 => n18312, A2 => n19065, B1 => n25983, B2 => 
                           n19193, ZN => n25812);
   U1795 : AOI22_X1 port map( A1 => n18320, A2 => n18969, B1 => n18319, B2 => 
                           n19257, ZN => n25811);
   U1796 : AOI22_X1 port map( A1 => n18309, A2 => n18937, B1 => n25829, B2 => 
                           n19097, ZN => n25810);
   U1797 : NAND4_X1 port map( A1 => n25813, A2 => n25812, A3 => n25811, A4 => 
                           n25810, ZN => n25814);
   U1798 : NOR2_X1 port map( A1 => n25815, A2 => n25814, ZN => n25827);
   U1799 : AOI22_X1 port map( A1 => n25961, A2 => n18394, B1 => n18426, B2 => 
                           n25992, ZN => n25819);
   U1800 : AOI22_X1 port map( A1 => n18458, A2 => n19402, B1 => n18554, B2 => 
                           n25940, ZN => n25818);
   U1801 : AOI22_X1 port map( A1 => n18586, A2 => n26754, B1 => n18522, B2 => 
                           n25939, ZN => n25817);
   U1802 : AOI22_X1 port map( A1 => n18490, A2 => n25993, B1 => n18617, B2 => 
                           n25995, ZN => n25816);
   U1803 : NAND4_X1 port map( A1 => n25819, A2 => n25818, A3 => n25817, A4 => 
                           n25816, ZN => n25825);
   U1804 : AOI22_X1 port map( A1 => n18291, A2 => n18649, B1 => n18681, B2 => 
                           n25992, ZN => n25823);
   U1805 : AOI22_X1 port map( A1 => n18745, A2 => n25993, B1 => n18841, B2 => 
                           n25994, ZN => n25822);
   U1806 : AOI22_X1 port map( A1 => n18873, A2 => n26755, B1 => n18809, B2 => 
                           n25940, ZN => n25821);
   U1807 : AOI22_X1 port map( A1 => n18713, A2 => n18288, B1 => n18777, B2 => 
                           n25939, ZN => n25820);
   U1808 : NAND4_X1 port map( A1 => n25823, A2 => n25822, A3 => n25821, A4 => 
                           n25820, ZN => n25824);
   U1809 : AOI22_X1 port map( A1 => n26009, A2 => n25825, B1 => n26007, B2 => 
                           n25824, ZN => n25826);
   U1810 : OAI21_X1 port map( B1 => n25828, B2 => n25827, A => n25826, ZN => 
                           OUT2(7));
   U1811 : AOI22_X1 port map( A1 => n18321, A2 => n19386, B1 => n18320, B2 => 
                           n18970, ZN => n25833);
   U1812 : AOI22_X1 port map( A1 => n18317, A2 => n19130, B1 => n25985, B2 => 
                           n19322, ZN => n25832);
   U1813 : AOI22_X1 port map( A1 => n18312, A2 => n19066, B1 => n25982, B2 => 
                           n19162, ZN => n25831);
   U1814 : AOI22_X1 port map( A1 => n25829, A2 => n19098, B1 => n18319, B2 => 
                           n19258, ZN => n25830);
   U1815 : NAND4_X1 port map( A1 => n25833, A2 => n25832, A3 => n25831, A4 => 
                           n25830, ZN => n25839);
   U1816 : AOI22_X1 port map( A1 => n18316, A2 => n18906, B1 => n25983, B2 => 
                           n19194, ZN => n25837);
   U1817 : AOI22_X1 port map( A1 => n18309, A2 => n18938, B1 => n25923, B2 => 
                           n19354, ZN => n25836);
   U1818 : AOI22_X1 port map( A1 => n25984, A2 => n19034, B1 => n25903, B2 => 
                           n19002, ZN => n25835);
   U1819 : AOI22_X1 port map( A1 => n18315, A2 => n19290, B1 => n18322, B2 => 
                           n19226, ZN => n25834);
   U1820 : NAND4_X1 port map( A1 => n25837, A2 => n25836, A3 => n25835, A4 => 
                           n25834, ZN => n25838);
   U1821 : NOR2_X1 port map( A1 => n25839, A2 => n25838, ZN => n25851);
   U1822 : AOI22_X1 port map( A1 => n18618, A2 => n26755, B1 => n18587, B2 => 
                           n25994, ZN => n25843);
   U1823 : AOI22_X1 port map( A1 => n18291, A2 => n18395, B1 => n18427, B2 => 
                           n25992, ZN => n25842);
   U1824 : AOI22_X1 port map( A1 => n18491, A2 => n25993, B1 => n18523, B2 => 
                           n25939, ZN => n25841);
   U1825 : AOI22_X1 port map( A1 => n18459, A2 => n26001, B1 => n18555, B2 => 
                           n25940, ZN => n25840);
   U1826 : NAND4_X1 port map( A1 => n25843, A2 => n25842, A3 => n25841, A4 => 
                           n25840, ZN => n25849);
   U1827 : AOI22_X1 port map( A1 => n18746, A2 => n25993, B1 => n18810, B2 => 
                           n25940, ZN => n25847);
   U1828 : AOI22_X1 port map( A1 => n18291, A2 => n18650, B1 => n19402, B2 => 
                           n18714, ZN => n25846);
   U1829 : AOI22_X1 port map( A1 => n18874, A2 => n26755, B1 => n18842, B2 => 
                           n25994, ZN => n25845);
   U1830 : AOI22_X1 port map( A1 => n18682, A2 => n25992, B1 => n18778, B2 => 
                           n25939, ZN => n25844);
   U1831 : NAND4_X1 port map( A1 => n25847, A2 => n25846, A3 => n25845, A4 => 
                           n25844, ZN => n25848);
   U1832 : AOI22_X1 port map( A1 => n26009, A2 => n25849, B1 => n26007, B2 => 
                           n25848, ZN => n25850);
   U1833 : OAI21_X1 port map( B1 => n26012, B2 => n25851, A => n25850, ZN => 
                           OUT2(6));
   U1834 : AOI22_X1 port map( A1 => n18324, A2 => n19035, B1 => n18319, B2 => 
                           n19259, ZN => n25855);
   U1835 : AOI22_X1 port map( A1 => n18316, A2 => n18907, B1 => n18313, B2 => 
                           n19323, ZN => n25854);
   U1836 : AOI22_X1 port map( A1 => n25903, A2 => n19003, B1 => n18323, B2 => 
                           n19355, ZN => n25853);
   U1837 : AOI22_X1 port map( A1 => n18318, A2 => n19195, B1 => n18321, B2 => 
                           n19387, ZN => n25852);
   U1838 : NAND4_X1 port map( A1 => n25855, A2 => n25854, A3 => n25853, A4 => 
                           n25852, ZN => n25861);
   U1839 : AOI22_X1 port map( A1 => n25949, A2 => n19291, B1 => n25982, B2 => 
                           n19163, ZN => n25859);
   U1840 : AOI22_X1 port map( A1 => n25975, A2 => n18939, B1 => n18322, B2 => 
                           n19227, ZN => n25858);
   U1841 : AOI22_X1 port map( A1 => n18310, A2 => n19099, B1 => n18320, B2 => 
                           n18971, ZN => n25857);
   U1842 : AOI22_X1 port map( A1 => n18312, A2 => n19067, B1 => n18317, B2 => 
                           n19131, ZN => n25856);
   U1843 : NAND4_X1 port map( A1 => n25859, A2 => n25858, A3 => n25857, A4 => 
                           n25856, ZN => n25860);
   U1844 : NOR2_X1 port map( A1 => n25861, A2 => n25860, ZN => n25874);
   U1845 : AOI22_X1 port map( A1 => n18428, A2 => n25992, B1 => n18588, B2 => 
                           n25994, ZN => n25865);
   U1846 : AOI22_X1 port map( A1 => n18492, A2 => n25993, B1 => n18556, B2 => 
                           n25940, ZN => n25864);
   U1847 : AOI22_X1 port map( A1 => n18396, A2 => n25961, B1 => n18524, B2 => 
                           n25939, ZN => n25863);
   U1848 : AOI22_X1 port map( A1 => n18460, A2 => n19402, B1 => n18619, B2 => 
                           n26000, ZN => n25862);
   U1849 : NAND4_X1 port map( A1 => n25865, A2 => n25864, A3 => n25863, A4 => 
                           n25862, ZN => n25872);
   U1850 : AOI22_X1 port map( A1 => n18683, A2 => n25992, B1 => n18811, B2 => 
                           n25940, ZN => n25870);
   U1851 : AOI22_X1 port map( A1 => n18875, A2 => n26755, B1 => n18843, B2 => 
                           n25994, ZN => n25869);
   U1852 : AOI22_X1 port map( A1 => n25961, A2 => n18651, B1 => n18747, B2 => 
                           n25866, ZN => n25868);
   U1853 : AOI22_X1 port map( A1 => n18715, A2 => n26001, B1 => n18779, B2 => 
                           n25939, ZN => n25867);
   U1854 : NAND4_X1 port map( A1 => n25870, A2 => n25869, A3 => n25868, A4 => 
                           n25867, ZN => n25871);
   U1855 : AOI22_X1 port map( A1 => n26009, A2 => n25872, B1 => n26007, B2 => 
                           n25871, ZN => n25873);
   U1856 : OAI21_X1 port map( B1 => n26012, B2 => n25874, A => n25873, ZN => 
                           OUT2(5));
   U1857 : AOI22_X1 port map( A1 => n25928, A2 => n19068, B1 => n25981, B2 => 
                           n19260, ZN => n25878);
   U1858 : AOI22_X1 port map( A1 => n18317, A2 => n19132, B1 => n25985, B2 => 
                           n19324, ZN => n25877);
   U1859 : AOI22_X1 port map( A1 => n18321, A2 => n19388, B1 => n18311, B2 => 
                           n19004, ZN => n25876);
   U1860 : AOI22_X1 port map( A1 => n18310, A2 => n19100, B1 => n18322, B2 => 
                           n19228, ZN => n25875);
   U1861 : NAND4_X1 port map( A1 => n25878, A2 => n25877, A3 => n25876, A4 => 
                           n25875, ZN => n25884);
   U1862 : AOI22_X1 port map( A1 => n18324, A2 => n19036, B1 => n18315, B2 => 
                           n19292, ZN => n25882);
   U1863 : AOI22_X1 port map( A1 => n25975, A2 => n18940, B1 => n18314, B2 => 
                           n19164, ZN => n25881);
   U1864 : AOI22_X1 port map( A1 => n18318, A2 => n19196, B1 => n25902, B2 => 
                           n18972, ZN => n25880);
   U1865 : AOI22_X1 port map( A1 => n25922, A2 => n18908, B1 => n25923, B2 => 
                           n19356, ZN => n25879);
   U1866 : NAND4_X1 port map( A1 => n25882, A2 => n25881, A3 => n25880, A4 => 
                           n25879, ZN => n25883);
   U1867 : NOR2_X1 port map( A1 => n25884, A2 => n25883, ZN => n25897);
   U1868 : AOI22_X1 port map( A1 => n18397, A2 => n25961, B1 => n18525, B2 => 
                           n25939, ZN => n25888);
   U1869 : AOI22_X1 port map( A1 => n18288, A2 => n18461, B1 => n18493, B2 => 
                           n26756, ZN => n25887);
   U1870 : AOI22_X1 port map( A1 => n18557, A2 => n26757, B1 => n18589, B2 => 
                           n26754, ZN => n25886);
   U1871 : AOI22_X1 port map( A1 => n18429, A2 => n25992, B1 => n18620, B2 => 
                           n25995, ZN => n25885);
   U1872 : NAND4_X1 port map( A1 => n25888, A2 => n25887, A3 => n25886, A4 => 
                           n25885, ZN => n25895);
   U1873 : AOI22_X1 port map( A1 => n18812, A2 => n25889, B1 => n18844, B2 => 
                           n25994, ZN => n25893);
   U1874 : AOI22_X1 port map( A1 => n18684, A2 => n25992, B1 => n18780, B2 => 
                           n25939, ZN => n25892);
   U1875 : AOI22_X1 port map( A1 => n26001, A2 => n18716, B1 => n18876, B2 => 
                           n25995, ZN => n25891);
   U1876 : AOI22_X1 port map( A1 => n18291, A2 => n18652, B1 => n18748, B2 => 
                           n25993, ZN => n25890);
   U1877 : NAND4_X1 port map( A1 => n25893, A2 => n25892, A3 => n25891, A4 => 
                           n25890, ZN => n25894);
   U1878 : AOI22_X1 port map( A1 => n26009, A2 => n25895, B1 => n26007, B2 => 
                           n25894, ZN => n25896);
   U1879 : OAI21_X1 port map( B1 => n26012, B2 => n25897, A => n25896, ZN => 
                           OUT2(4));
   U1880 : AOI22_X1 port map( A1 => n18310, A2 => n19101, B1 => n18323, B2 => 
                           n19357, ZN => n25901);
   U1881 : AOI22_X1 port map( A1 => n25950, A2 => n19133, B1 => n18319, B2 => 
                           n19261, ZN => n25900);
   U1882 : AOI22_X1 port map( A1 => n18315, A2 => n19293, B1 => n18314, B2 => 
                           n19165, ZN => n25899);
   U1883 : AOI22_X1 port map( A1 => n25928, A2 => n19069, B1 => n18321, B2 => 
                           n19389, ZN => n25898);
   U1884 : NAND4_X1 port map( A1 => n25901, A2 => n25900, A3 => n25899, A4 => 
                           n25898, ZN => n25909);
   U1885 : AOI22_X1 port map( A1 => n18309, A2 => n18941, B1 => n18318, B2 => 
                           n19197, ZN => n25907);
   U1886 : AOI22_X1 port map( A1 => n18324, A2 => n19037, B1 => n18322, B2 => 
                           n19229, ZN => n25906);
   U1887 : AOI22_X1 port map( A1 => n25922, A2 => n18909, B1 => n18313, B2 => 
                           n19325, ZN => n25905);
   U1888 : AOI22_X1 port map( A1 => n25903, A2 => n19005, B1 => n25902, B2 => 
                           n18973, ZN => n25904);
   U1889 : NAND4_X1 port map( A1 => n25907, A2 => n25906, A3 => n25905, A4 => 
                           n25904, ZN => n25908);
   U1890 : NOR2_X1 port map( A1 => n25909, A2 => n25908, ZN => n25921);
   U1891 : AOI22_X1 port map( A1 => n18291, A2 => n18398, B1 => n18430, B2 => 
                           n25992, ZN => n25913);
   U1892 : AOI22_X1 port map( A1 => n18494, A2 => n25993, B1 => n18526, B2 => 
                           n25939, ZN => n25912);
   U1893 : AOI22_X1 port map( A1 => n18462, A2 => n19402, B1 => n18590, B2 => 
                           n25994, ZN => n25911);
   U1894 : AOI22_X1 port map( A1 => n18621, A2 => n26000, B1 => n18558, B2 => 
                           n25940, ZN => n25910);
   U1895 : NAND4_X1 port map( A1 => n25913, A2 => n25912, A3 => n25911, A4 => 
                           n25910, ZN => n25919);
   U1896 : AOI22_X1 port map( A1 => n18291, A2 => n18653, B1 => n18749, B2 => 
                           n26756, ZN => n25917);
   U1897 : AOI22_X1 port map( A1 => n18717, A2 => n26001, B1 => n18845, B2 => 
                           n25994, ZN => n25916);
   U1898 : AOI22_X1 port map( A1 => n18685, A2 => n26758, B1 => n18877, B2 => 
                           n25995, ZN => n25915);
   U1899 : AOI22_X1 port map( A1 => n18813, A2 => n26757, B1 => n18781, B2 => 
                           n25939, ZN => n25914);
   U1900 : NAND4_X1 port map( A1 => n25917, A2 => n25916, A3 => n25915, A4 => 
                           n25914, ZN => n25918);
   U1901 : AOI22_X1 port map( A1 => n26009, A2 => n25919, B1 => n26007, B2 => 
                           n25918, ZN => n25920);
   U1902 : OAI21_X1 port map( B1 => n26012, B2 => n25921, A => n25920, ZN => 
                           OUT2(3));
   U1903 : AOI22_X1 port map( A1 => n25922, A2 => n18910, B1 => n25984, B2 => 
                           n19038, ZN => n25927);
   U1904 : AOI22_X1 port map( A1 => n18322, A2 => n19230, B1 => n18320, B2 => 
                           n18974, ZN => n25926);
   U1905 : AOI22_X1 port map( A1 => n18315, A2 => n19294, B1 => n18321, B2 => 
                           n19390, ZN => n25925);
   U1906 : AOI22_X1 port map( A1 => n25983, A2 => n19198, B1 => n25923, B2 => 
                           n19358, ZN => n25924);
   U1907 : NAND4_X1 port map( A1 => n25927, A2 => n25926, A3 => n25925, A4 => 
                           n25924, ZN => n25934);
   U1908 : AOI22_X1 port map( A1 => n18311, A2 => n19006, B1 => n18319, B2 => 
                           n19262, ZN => n25932);
   U1909 : AOI22_X1 port map( A1 => n25928, A2 => n19070, B1 => n18314, B2 => 
                           n19166, ZN => n25931);
   U1910 : AOI22_X1 port map( A1 => n18317, A2 => n19134, B1 => n18313, B2 => 
                           n19326, ZN => n25930);
   U1911 : AOI22_X1 port map( A1 => n25975, A2 => n18942, B1 => n18310, B2 => 
                           n19102, ZN => n25929);
   U1912 : NAND4_X1 port map( A1 => n25932, A2 => n25931, A3 => n25930, A4 => 
                           n25929, ZN => n25933);
   U1913 : NOR2_X1 port map( A1 => n25934, A2 => n25933, ZN => n25948);
   U1914 : AOI22_X1 port map( A1 => n18431, A2 => n25992, B1 => n18559, B2 => 
                           n25940, ZN => n25938);
   U1915 : AOI22_X1 port map( A1 => n18463, A2 => n19402, B1 => n18495, B2 => 
                           n26756, ZN => n25937);
   U1916 : AOI22_X1 port map( A1 => n18591, A2 => n26754, B1 => n18527, B2 => 
                           n25939, ZN => n25936);
   U1917 : AOI22_X1 port map( A1 => n18399, A2 => n18291, B1 => n18622, B2 => 
                           n25995, ZN => n25935);
   U1918 : NAND4_X1 port map( A1 => n25938, A2 => n25937, A3 => n25936, A4 => 
                           n25935, ZN => n25946);
   U1919 : AOI22_X1 port map( A1 => n25961, A2 => n18654, B1 => n18686, B2 => 
                           n25992, ZN => n25944);
   U1920 : AOI22_X1 port map( A1 => n18718, A2 => n18288, B1 => n18846, B2 => 
                           n25994, ZN => n25943);
   U1921 : AOI22_X1 port map( A1 => n18750, A2 => n25993, B1 => n18782, B2 => 
                           n25939, ZN => n25942);
   U1922 : AOI22_X1 port map( A1 => n18878, A2 => n26000, B1 => n18814, B2 => 
                           n25940, ZN => n25941);
   U1923 : NAND4_X1 port map( A1 => n25944, A2 => n25943, A3 => n25942, A4 => 
                           n25941, ZN => n25945);
   U1924 : AOI22_X1 port map( A1 => n26009, A2 => n25946, B1 => n26007, B2 => 
                           n25945, ZN => n25947);
   U1925 : OAI21_X1 port map( B1 => n26012, B2 => n25948, A => n25947, ZN => 
                           OUT2(2));
   U1926 : AOI22_X1 port map( A1 => n18312, A2 => n19071, B1 => n25949, B2 => 
                           n19295, ZN => n25954);
   U1927 : AOI22_X1 port map( A1 => n18324, A2 => n19039, B1 => n18319, B2 => 
                           n19263, ZN => n25953);
   U1928 : AOI22_X1 port map( A1 => n25950, A2 => n19135, B1 => n18313, B2 => 
                           n19327, ZN => n25952);
   U1929 : AOI22_X1 port map( A1 => n18321, A2 => n19391, B1 => n18310, B2 => 
                           n19103, ZN => n25951);
   U1930 : NAND4_X1 port map( A1 => n25954, A2 => n25953, A3 => n25952, A4 => 
                           n25951, ZN => n25960);
   U1931 : AOI22_X1 port map( A1 => n18309, A2 => n18943, B1 => n25976, B2 => 
                           n19231, ZN => n25958);
   U1932 : AOI22_X1 port map( A1 => n18314, A2 => n19167, B1 => n18320, B2 => 
                           n18975, ZN => n25957);
   U1933 : AOI22_X1 port map( A1 => n18316, A2 => n18911, B1 => n18323, B2 => 
                           n19359, ZN => n25956);
   U1934 : AOI22_X1 port map( A1 => n25983, A2 => n19199, B1 => n18311, B2 => 
                           n19007, ZN => n25955);
   U1935 : NAND4_X1 port map( A1 => n25958, A2 => n25957, A3 => n25956, A4 => 
                           n25955, ZN => n25959);
   U1936 : NOR2_X1 port map( A1 => n25960, A2 => n25959, ZN => n25973);
   U1937 : AOI22_X1 port map( A1 => n25961, A2 => n18400, B1 => n18432, B2 => 
                           n25992, ZN => n25965);
   U1938 : AOI22_X1 port map( A1 => n18592, A2 => n26754, B1 => n18528, B2 => 
                           n26759, ZN => n25964);
   U1939 : AOI22_X1 port map( A1 => n18496, A2 => n25993, B1 => n18560, B2 => 
                           n26757, ZN => n25963);
   U1940 : AOI22_X1 port map( A1 => n18464, A2 => n19402, B1 => n18623, B2 => 
                           n25995, ZN => n25962);
   U1941 : NAND4_X1 port map( A1 => n25965, A2 => n25964, A3 => n25963, A4 => 
                           n25962, ZN => n25971);
   U1942 : AOI22_X1 port map( A1 => n18751, A2 => n25993, B1 => n18815, B2 => 
                           n26757, ZN => n25969);
   U1943 : AOI22_X1 port map( A1 => n18288, A2 => n18719, B1 => n18291, B2 => 
                           n18655, ZN => n25968);
   U1944 : AOI22_X1 port map( A1 => n18687, A2 => n25992, B1 => n18847, B2 => 
                           n25994, ZN => n25967);
   U1945 : AOI22_X1 port map( A1 => n18879, A2 => n26000, B1 => n18783, B2 => 
                           n26759, ZN => n25966);
   U1946 : NAND4_X1 port map( A1 => n25969, A2 => n25968, A3 => n25967, A4 => 
                           n25966, ZN => n25970);
   U1947 : AOI22_X1 port map( A1 => n26009, A2 => n25971, B1 => n26007, B2 => 
                           n25970, ZN => n25972);
   U1948 : OAI21_X1 port map( B1 => n26012, B2 => n25973, A => n25972, ZN => 
                           OUT2(1));
   U1949 : AOI22_X1 port map( A1 => n25974, A2 => n19392, B1 => n18310, B2 => 
                           n19104, ZN => n25980);
   U1950 : AOI22_X1 port map( A1 => n18316, A2 => n18912, B1 => n25975, B2 => 
                           n18944, ZN => n25979);
   U1951 : AOI22_X1 port map( A1 => n18311, A2 => n19008, B1 => n25976, B2 => 
                           n19232, ZN => n25978);
   U1952 : AOI22_X1 port map( A1 => n18315, A2 => n19296, B1 => n18320, B2 => 
                           n18976, ZN => n25977);
   U1953 : NAND4_X1 port map( A1 => n25980, A2 => n25979, A3 => n25978, A4 => 
                           n25977, ZN => n25991);
   U1954 : AOI22_X1 port map( A1 => n25982, A2 => n19168, B1 => n25981, B2 => 
                           n19264, ZN => n25989);
   U1955 : AOI22_X1 port map( A1 => n25983, A2 => n19200, B1 => n18323, B2 => 
                           n19360, ZN => n25988);
   U1956 : AOI22_X1 port map( A1 => n18312, A2 => n19072, B1 => n25984, B2 => 
                           n19040, ZN => n25987);
   U1957 : AOI22_X1 port map( A1 => n18317, A2 => n19136, B1 => n25985, B2 => 
                           n19328, ZN => n25986);
   U1958 : NAND4_X1 port map( A1 => n25989, A2 => n25988, A3 => n25987, A4 => 
                           n25986, ZN => n25990);
   U1959 : NOR2_X1 port map( A1 => n25991, A2 => n25990, ZN => n26011);
   U1960 : AOI22_X1 port map( A1 => n18561, A2 => n26757, B1 => n18529, B2 => 
                           n26759, ZN => n25999);
   U1961 : AOI22_X1 port map( A1 => n18497, A2 => n25993, B1 => n18433, B2 => 
                           n25992, ZN => n25998);
   U1962 : AOI22_X1 port map( A1 => n18465, A2 => n18288, B1 => n18593, B2 => 
                           n25994, ZN => n25997);
   U1963 : AOI22_X1 port map( A1 => n18401, A2 => n18291, B1 => n18624, B2 => 
                           n25995, ZN => n25996);
   U1964 : NAND4_X1 port map( A1 => n25999, A2 => n25998, A3 => n25997, A4 => 
                           n25996, ZN => n26008);
   U1965 : AOI22_X1 port map( A1 => n18752, A2 => n26756, B1 => n18848, B2 => 
                           n26754, ZN => n26005);
   U1966 : AOI22_X1 port map( A1 => n18688, A2 => n26758, B1 => n18880, B2 => 
                           n26000, ZN => n26004);
   U1967 : AOI22_X1 port map( A1 => n26001, A2 => n18720, B1 => n19401, B2 => 
                           n18656, ZN => n26003);
   U1968 : AOI22_X1 port map( A1 => n18816, A2 => n26757, B1 => n18784, B2 => 
                           n26759, ZN => n26002);
   U1969 : NAND4_X1 port map( A1 => n26005, A2 => n26004, A3 => n26003, A4 => 
                           n26002, ZN => n26006);
   U1970 : AOI22_X1 port map( A1 => n26009, A2 => n26008, B1 => n26007, B2 => 
                           n26006, ZN => n26010);
   U1971 : OAI21_X1 port map( B1 => n26012, B2 => n26011, A => n26010, ZN => 
                           OUT2(0));
   U1972 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n26016)
                           ;
   U1973 : NOR2_X1 port map( A1 => n1518, A2 => n26016, ZN => n11132);
   U1974 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n26013);
   U1975 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => n26013, ZN => n25158);
   U1976 : INV_X1 port map( A => ADD_RD1(3), ZN => n26014);
   U1977 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n26014, ZN => n26015);
   U1978 : NOR2_X1 port map( A1 => n26015, A2 => n25158, ZN => n11154);
   U1979 : NOR2_X1 port map( A1 => n1518, A2 => n26015, ZN => n11136);
   U1980 : NOR2_X1 port map( A1 => n26016, A2 => n1519, ZN => n11153);
   U1981 : NOR2_X1 port map( A1 => n26015, A2 => n1517, ZN => n11139);
   U1982 : NOR2_X1 port map( A1 => n26015, A2 => n1516, ZN => n11152);
   U1983 : NOR2_X1 port map( A1 => n26015, A2 => n1514, ZN => n11141);
   U1984 : NOR2_X1 port map( A1 => n26015, A2 => n1519, ZN => n11151);
   U1985 : NOR2_X1 port map( A1 => n26016, A2 => n25158, ZN => n11137);
   U1986 : NOR2_X1 port map( A1 => n26016, A2 => n1516, ZN => n11150);
   U1987 : NOR2_X1 port map( A1 => n26015, A2 => n25157, ZN => n11138);
   U1988 : NOR2_X1 port map( A1 => n26016, A2 => n25157, ZN => n11149);
   U1989 : NOR2_X1 port map( A1 => n26015, A2 => n1515, ZN => n11133);
   U1990 : NOR2_X1 port map( A1 => n26016, A2 => n1514, ZN => n11140);
   U1991 : NOR2_X1 port map( A1 => n26016, A2 => n1517, ZN => n11142);
   U1992 : NOR2_X1 port map( A1 => n26016, A2 => n1515, ZN => n11143);
   U1993 : CLKBUF_X1 port map( A => n18299, Z => n26695);
   U1994 : CLKBUF_X1 port map( A => n18294, Z => n26726);
   U1995 : AOI22_X1 port map( A1 => n19361, A2 => n26695, B1 => n19297, B2 => 
                           n26726, ZN => n26020);
   U1996 : AOI22_X1 port map( A1 => n18913, A2 => n18296, B1 => n19073, B2 => 
                           n18298, ZN => n26019);
   U1997 : CLKBUF_X1 port map( A => n18302, Z => n26667);
   U1998 : AOI22_X1 port map( A1 => n18977, A2 => n26667, B1 => n19233, B2 => 
                           n18295, ZN => n26018);
   U1999 : CLKBUF_X1 port map( A => n18304, Z => n26666);
   U2000 : AOI22_X1 port map( A1 => n19041, A2 => n26666, B1 => n19105, B2 => 
                           n18303, ZN => n26017);
   U2001 : NAND4_X1 port map( A1 => n26020, A2 => n26019, A3 => n26018, A4 => 
                           n26017, ZN => n26026);
   U2002 : AOI22_X1 port map( A1 => n19137, A2 => n18308, B1 => n19201, B2 => 
                           n18305, ZN => n26024);
   U2003 : AOI22_X1 port map( A1 => n19169, A2 => n18293, B1 => n19329, B2 => 
                           n18297, ZN => n26023);
   U2004 : AOI22_X1 port map( A1 => n19009, A2 => n18307, B1 => n18945, B2 => 
                           n18301, ZN => n26022);
   U2005 : AOI22_X1 port map( A1 => n18881, A2 => n18306, B1 => n19265, B2 => 
                           n18300, ZN => n26021);
   U2006 : NAND4_X1 port map( A1 => n26024, A2 => n26023, A3 => n26022, A4 => 
                           n26021, ZN => n26025);
   U2007 : NOR2_X1 port map( A1 => n26026, A2 => n26025, ZN => n26038);
   U2008 : NOR3_X1 port map( A1 => n18369, A2 => n20464, A3 => n26689, ZN => 
                           n26478);
   U2009 : CLKBUF_X1 port map( A => n26478, Z => n26523);
   U2010 : CLKBUF_X1 port map( A => n18364, Z => n26737);
   U2011 : AOI22_X1 port map( A1 => n18530, A2 => n18367, B1 => n18466, B2 => 
                           n26737, ZN => n26030);
   U2012 : AOI22_X1 port map( A1 => n18434, A2 => n19399, B1 => n18371, B2 => 
                           n19400, ZN => n26029);
   U2013 : INV_X1 port map( A => n25153, ZN => n26742);
   U2014 : CLKBUF_X1 port map( A => n18363, Z => n26680);
   U2015 : AOI22_X1 port map( A1 => n18498, A2 => n26742, B1 => n18402, B2 => 
                           n26680, ZN => n26028);
   U2016 : INV_X1 port map( A => n25152, ZN => n26736);
   U2017 : AOI22_X1 port map( A1 => n18562, A2 => n26736, B1 => n18594, B2 => 
                           n18368, ZN => n26027);
   U2018 : NAND4_X1 port map( A1 => n26030, A2 => n26029, A3 => n26028, A4 => 
                           n26027, ZN => n26036);
   U2019 : NOR3_X1 port map( A1 => n20464, A2 => n20430, A3 => n26689, ZN => 
                           n26256);
   U2020 : CLKBUF_X1 port map( A => n26742, Z => n26674);
   U2021 : AOI22_X1 port map( A1 => n18753, A2 => n26674, B1 => n18689, B2 => 
                           n18290, ZN => n26034);
   U2022 : AOI22_X1 port map( A1 => n18785, A2 => n18367, B1 => n18849, B2 => 
                           n19398, ZN => n26033);
   U2023 : AOI22_X1 port map( A1 => n18817, A2 => n26761, B1 => n18657, B2 => 
                           n18363, ZN => n26032);
   U2024 : AOI22_X1 port map( A1 => n18721, A2 => n19397, B1 => n18625, B2 => 
                           n18292, ZN => n26031);
   U2025 : NAND4_X1 port map( A1 => n26034, A2 => n26033, A3 => n26032, A4 => 
                           n26031, ZN => n26035);
   U2026 : AOI22_X1 port map( A1 => n26523, A2 => n26036, B1 => n26256, B2 => 
                           n26035, ZN => n26037);
   U2027 : OAI21_X1 port map( B1 => n26689, B2 => n26038, A => n26037, ZN => 
                           OUT1(31));
   U2028 : AOI22_X1 port map( A1 => n18978, A2 => n18302, B1 => n18946, B2 => 
                           n18301, ZN => n26042);
   U2029 : AOI22_X1 port map( A1 => n18914, A2 => n18296, B1 => n19298, B2 => 
                           n18294, ZN => n26041);
   U2030 : AOI22_X1 port map( A1 => n19074, A2 => n18298, B1 => n19170, B2 => 
                           n18293, ZN => n26040);
   U2031 : CLKBUF_X1 port map( A => n18307, Z => n26725);
   U2032 : AOI22_X1 port map( A1 => n19010, A2 => n26725, B1 => n19042, B2 => 
                           n26666, ZN => n26039);
   U2033 : NAND4_X1 port map( A1 => n26042, A2 => n26041, A3 => n26040, A4 => 
                           n26039, ZN => n26048);
   U2034 : AOI22_X1 port map( A1 => n19266, A2 => n18300, B1 => n19234, B2 => 
                           n18295, ZN => n26046);
   U2035 : AOI22_X1 port map( A1 => n19330, A2 => n18297, B1 => n19202, B2 => 
                           n18305, ZN => n26045);
   U2036 : CLKBUF_X1 port map( A => n18303, Z => n26637);
   U2037 : AOI22_X1 port map( A1 => n19362, A2 => n18299, B1 => n19106, B2 => 
                           n26637, ZN => n26044);
   U2038 : AOI22_X1 port map( A1 => n19138, A2 => n18308, B1 => n18882, B2 => 
                           n18306, ZN => n26043);
   U2039 : NAND4_X1 port map( A1 => n26046, A2 => n26045, A3 => n26044, A4 => 
                           n26043, ZN => n26047);
   U2040 : NOR2_X1 port map( A1 => n26048, A2 => n26047, ZN => n26060);
   U2041 : AOI22_X1 port map( A1 => n18435, A2 => n19399, B1 => n18467, B2 => 
                           n18364, ZN => n26052);
   U2042 : AOI22_X1 port map( A1 => n18403, A2 => n19396, B1 => n18563, B2 => 
                           n26736, ZN => n26051);
   U2043 : CLKBUF_X1 port map( A => n18367, Z => n26624);
   U2044 : AOI22_X1 port map( A1 => n18531, A2 => n26624, B1 => n18499, B2 => 
                           n26760, ZN => n26050);
   U2045 : CLKBUF_X1 port map( A => n18292, Z => n26703);
   U2046 : AOI22_X1 port map( A1 => n18595, A2 => n18368, B1 => n18372, B2 => 
                           n26703, ZN => n26049);
   U2047 : NAND4_X1 port map( A1 => n26052, A2 => n26051, A3 => n26050, A4 => 
                           n26049, ZN => n26058);
   U2048 : CLKBUF_X1 port map( A => n26256, Z => n26748);
   U2049 : AOI22_X1 port map( A1 => n18754, A2 => n26742, B1 => n18850, B2 => 
                           n18368, ZN => n26056);
   U2050 : AOI22_X1 port map( A1 => n18818, A2 => n26736, B1 => n18722, B2 => 
                           n26737, ZN => n26055);
   U2051 : AOI22_X1 port map( A1 => n18658, A2 => n26680, B1 => n18626, B2 => 
                           n18292, ZN => n26054);
   U2052 : AOI22_X1 port map( A1 => n18690, A2 => n18290, B1 => n18786, B2 => 
                           n26624, ZN => n26053);
   U2053 : NAND4_X1 port map( A1 => n26056, A2 => n26055, A3 => n26054, A4 => 
                           n26053, ZN => n26057);
   U2054 : AOI22_X1 port map( A1 => n26523, A2 => n26058, B1 => n26748, B2 => 
                           n26057, ZN => n26059);
   U2055 : OAI21_X1 port map( B1 => n26689, B2 => n26060, A => n26059, ZN => 
                           OUT1(30));
   U2056 : AOI22_X1 port map( A1 => n19363, A2 => n18299, B1 => n19299, B2 => 
                           n18294, ZN => n26064);
   U2057 : AOI22_X1 port map( A1 => n18979, A2 => n26667, B1 => n19235, B2 => 
                           n18295, ZN => n26063);
   U2058 : CLKBUF_X1 port map( A => n18305, Z => n26719);
   U2059 : CLKBUF_X1 port map( A => n18308, Z => n26694);
   U2060 : AOI22_X1 port map( A1 => n19203, A2 => n26719, B1 => n19139, B2 => 
                           n26694, ZN => n26062);
   U2061 : AOI22_X1 port map( A1 => n19043, A2 => n18304, B1 => n19011, B2 => 
                           n18307, ZN => n26061);
   U2062 : NAND4_X1 port map( A1 => n26064, A2 => n26063, A3 => n26062, A4 => 
                           n26061, ZN => n26070);
   U2063 : AOI22_X1 port map( A1 => n19267, A2 => n18300, B1 => n19331, B2 => 
                           n18297, ZN => n26068);
   U2064 : AOI22_X1 port map( A1 => n19171, A2 => n18293, B1 => n19107, B2 => 
                           n18303, ZN => n26067);
   U2065 : CLKBUF_X1 port map( A => n18306, Z => n26696);
   U2066 : AOI22_X1 port map( A1 => n19075, A2 => n18298, B1 => n18883, B2 => 
                           n26696, ZN => n26066);
   U2067 : AOI22_X1 port map( A1 => n18915, A2 => n18296, B1 => n18947, B2 => 
                           n18301, ZN => n26065);
   U2068 : NAND4_X1 port map( A1 => n26068, A2 => n26067, A3 => n26066, A4 => 
                           n26065, ZN => n26069);
   U2069 : NOR2_X1 port map( A1 => n26070, A2 => n26069, ZN => n26082);
   U2070 : AOI22_X1 port map( A1 => n18468, A2 => n18364, B1 => n18436, B2 => 
                           n19399, ZN => n26074);
   U2071 : AOI22_X1 port map( A1 => n18596, A2 => n19398, B1 => n18532, B2 => 
                           n18367, ZN => n26073);
   U2072 : AOI22_X1 port map( A1 => n18500, A2 => n26742, B1 => n18373, B2 => 
                           n19400, ZN => n26072);
   U2073 : AOI22_X1 port map( A1 => n18564, A2 => n26761, B1 => n18404, B2 => 
                           n18363, ZN => n26071);
   U2074 : NAND4_X1 port map( A1 => n26074, A2 => n26073, A3 => n26072, A4 => 
                           n26071, ZN => n26080);
   U2075 : CLKBUF_X1 port map( A => n18290, Z => n26734);
   U2076 : AOI22_X1 port map( A1 => n18851, A2 => n18368, B1 => n18691, B2 => 
                           n26734, ZN => n26078);
   U2077 : AOI22_X1 port map( A1 => n18787, A2 => n26624, B1 => n18627, B2 => 
                           n18292, ZN => n26077);
   U2078 : AOI22_X1 port map( A1 => n18723, A2 => n19397, B1 => n18659, B2 => 
                           n26680, ZN => n26076);
   U2079 : AOI22_X1 port map( A1 => n18819, A2 => n26761, B1 => n18755, B2 => 
                           n26760, ZN => n26075);
   U2080 : NAND4_X1 port map( A1 => n26078, A2 => n26077, A3 => n26076, A4 => 
                           n26075, ZN => n26079);
   U2081 : AOI22_X1 port map( A1 => n26523, A2 => n26080, B1 => n26256, B2 => 
                           n26079, ZN => n26081);
   U2082 : OAI21_X1 port map( B1 => n26689, B2 => n26082, A => n26081, ZN => 
                           OUT1(29));
   U2083 : AOI22_X1 port map( A1 => n19108, A2 => n18303, B1 => n19364, B2 => 
                           n26695, ZN => n26086);
   U2084 : AOI22_X1 port map( A1 => n18916, A2 => n18296, B1 => n19204, B2 => 
                           n18305, ZN => n26085);
   U2085 : AOI22_X1 port map( A1 => n19268, A2 => n18300, B1 => n19172, B2 => 
                           n18293, ZN => n26084);
   U2086 : CLKBUF_X1 port map( A => n18297, Z => n26720);
   U2087 : AOI22_X1 port map( A1 => n19236, A2 => n18295, B1 => n19332, B2 => 
                           n26720, ZN => n26083);
   U2088 : NAND4_X1 port map( A1 => n26086, A2 => n26085, A3 => n26084, A4 => 
                           n26083, ZN => n26092);
   U2089 : AOI22_X1 port map( A1 => n19140, A2 => n18308, B1 => n19076, B2 => 
                           n18298, ZN => n26090);
   U2090 : AOI22_X1 port map( A1 => n19044, A2 => n26666, B1 => n18980, B2 => 
                           n18302, ZN => n26089);
   U2091 : AOI22_X1 port map( A1 => n18948, A2 => n18301, B1 => n18884, B2 => 
                           n18306, ZN => n26088);
   U2092 : AOI22_X1 port map( A1 => n19300, A2 => n26726, B1 => n19012, B2 => 
                           n18307, ZN => n26087);
   U2093 : NAND4_X1 port map( A1 => n26090, A2 => n26089, A3 => n26088, A4 => 
                           n26087, ZN => n26091);
   U2094 : NOR2_X1 port map( A1 => n26092, A2 => n26091, ZN => n26104);
   U2095 : AOI22_X1 port map( A1 => n18405, A2 => n26680, B1 => n18501, B2 => 
                           n26760, ZN => n26096);
   U2096 : AOI22_X1 port map( A1 => n18437, A2 => n19399, B1 => n18374, B2 => 
                           n26703, ZN => n26095);
   U2097 : AOI22_X1 port map( A1 => n18597, A2 => n19398, B1 => n18469, B2 => 
                           n18364, ZN => n26094);
   U2098 : AOI22_X1 port map( A1 => n18565, A2 => n26761, B1 => n18533, B2 => 
                           n19395, ZN => n26093);
   U2099 : NAND4_X1 port map( A1 => n26096, A2 => n26095, A3 => n26094, A4 => 
                           n26093, ZN => n26102);
   U2100 : AOI22_X1 port map( A1 => n18692, A2 => n26734, B1 => n18660, B2 => 
                           n19396, ZN => n26100);
   U2101 : CLKBUF_X1 port map( A => n18368, Z => n26735);
   U2102 : AOI22_X1 port map( A1 => n18852, A2 => n26735, B1 => n18788, B2 => 
                           n18367, ZN => n26099);
   U2103 : AOI22_X1 port map( A1 => n18628, A2 => n26703, B1 => n18756, B2 => 
                           n26760, ZN => n26098);
   U2104 : CLKBUF_X1 port map( A => n26736, Z => n26675);
   U2105 : AOI22_X1 port map( A1 => n18724, A2 => n18364, B1 => n18820, B2 => 
                           n26675, ZN => n26097);
   U2106 : NAND4_X1 port map( A1 => n26100, A2 => n26099, A3 => n26098, A4 => 
                           n26097, ZN => n26101);
   U2107 : AOI22_X1 port map( A1 => n26523, A2 => n26102, B1 => n26748, B2 => 
                           n26101, ZN => n26103);
   U2108 : OAI21_X1 port map( B1 => n26689, B2 => n26104, A => n26103, ZN => 
                           OUT1(28));
   U2109 : AOI22_X1 port map( A1 => n19013, A2 => n26725, B1 => n19173, B2 => 
                           n18293, ZN => n26108);
   U2110 : AOI22_X1 port map( A1 => n18885, A2 => n18306, B1 => n19045, B2 => 
                           n18304, ZN => n26107);
   U2111 : AOI22_X1 port map( A1 => n19205, A2 => n26719, B1 => n19333, B2 => 
                           n18297, ZN => n26106);
   U2112 : CLKBUF_X1 port map( A => n18301, Z => n26716);
   U2113 : AOI22_X1 port map( A1 => n18917, A2 => n18296, B1 => n18949, B2 => 
                           n26716, ZN => n26105);
   U2114 : NAND4_X1 port map( A1 => n26108, A2 => n26107, A3 => n26106, A4 => 
                           n26105, ZN => n26114);
   U2115 : AOI22_X1 port map( A1 => n19237, A2 => n18295, B1 => n19109, B2 => 
                           n18303, ZN => n26112);
   U2116 : AOI22_X1 port map( A1 => n19141, A2 => n26694, B1 => n19301, B2 => 
                           n26726, ZN => n26111);
   U2117 : AOI22_X1 port map( A1 => n19365, A2 => n18299, B1 => n18981, B2 => 
                           n26667, ZN => n26110);
   U2118 : CLKBUF_X1 port map( A => n18298, Z => n26718);
   U2119 : CLKBUF_X1 port map( A => n18300, Z => n26665);
   U2120 : AOI22_X1 port map( A1 => n19077, A2 => n26718, B1 => n19269, B2 => 
                           n26665, ZN => n26109);
   U2121 : NAND4_X1 port map( A1 => n26112, A2 => n26111, A3 => n26110, A4 => 
                           n26109, ZN => n26113);
   U2122 : NOR2_X1 port map( A1 => n26114, A2 => n26113, ZN => n26126);
   U2123 : AOI22_X1 port map( A1 => n18566, A2 => n26736, B1 => n18375, B2 => 
                           n18292, ZN => n26118);
   U2124 : AOI22_X1 port map( A1 => n18470, A2 => n26737, B1 => n18598, B2 => 
                           n19398, ZN => n26117);
   U2125 : AOI22_X1 port map( A1 => n18534, A2 => n26624, B1 => n18502, B2 => 
                           n26760, ZN => n26116);
   U2126 : AOI22_X1 port map( A1 => n18406, A2 => n18363, B1 => n18438, B2 => 
                           n19399, ZN => n26115);
   U2127 : NAND4_X1 port map( A1 => n26118, A2 => n26117, A3 => n26116, A4 => 
                           n26115, ZN => n26124);
   U2128 : AOI22_X1 port map( A1 => n18821, A2 => n26761, B1 => n18853, B2 => 
                           n26735, ZN => n26122);
   U2129 : AOI22_X1 port map( A1 => n18629, A2 => n19400, B1 => n18757, B2 => 
                           n26674, ZN => n26121);
   U2130 : AOI22_X1 port map( A1 => n18693, A2 => n18290, B1 => n18661, B2 => 
                           n18363, ZN => n26120);
   U2131 : AOI22_X1 port map( A1 => n18789, A2 => n18367, B1 => n18725, B2 => 
                           n26737, ZN => n26119);
   U2132 : NAND4_X1 port map( A1 => n26122, A2 => n26121, A3 => n26120, A4 => 
                           n26119, ZN => n26123);
   U2133 : AOI22_X1 port map( A1 => n26523, A2 => n26124, B1 => n26256, B2 => 
                           n26123, ZN => n26125);
   U2134 : OAI21_X1 port map( B1 => n26689, B2 => n26126, A => n26125, ZN => 
                           OUT1(27));
   U2135 : AOI22_X1 port map( A1 => n18982, A2 => n18302, B1 => n18918, B2 => 
                           n18296, ZN => n26130);
   U2136 : CLKBUF_X1 port map( A => n18293, Z => n26717);
   U2137 : AOI22_X1 port map( A1 => n19174, A2 => n26717, B1 => n19014, B2 => 
                           n18307, ZN => n26129);
   U2138 : AOI22_X1 port map( A1 => n19206, A2 => n26719, B1 => n19142, B2 => 
                           n18308, ZN => n26128);
   U2139 : AOI22_X1 port map( A1 => n19078, A2 => n18298, B1 => n19334, B2 => 
                           n26720, ZN => n26127);
   U2140 : NAND4_X1 port map( A1 => n26130, A2 => n26129, A3 => n26128, A4 => 
                           n26127, ZN => n26136);
   U2141 : AOI22_X1 port map( A1 => n18886, A2 => n18306, B1 => n18950, B2 => 
                           n18301, ZN => n26134);
   U2142 : AOI22_X1 port map( A1 => n19302, A2 => n18294, B1 => n19270, B2 => 
                           n18300, ZN => n26133);
   U2143 : AOI22_X1 port map( A1 => n19110, A2 => n18303, B1 => n19366, B2 => 
                           n26695, ZN => n26132);
   U2144 : CLKBUF_X1 port map( A => n18295, Z => n26727);
   U2145 : AOI22_X1 port map( A1 => n19046, A2 => n18304, B1 => n19238, B2 => 
                           n26727, ZN => n26131);
   U2146 : NAND4_X1 port map( A1 => n26134, A2 => n26133, A3 => n26132, A4 => 
                           n26131, ZN => n26135);
   U2147 : NOR2_X1 port map( A1 => n26136, A2 => n26135, ZN => n26148);
   U2148 : AOI22_X1 port map( A1 => n18407, A2 => n26680, B1 => n18471, B2 => 
                           n26737, ZN => n26140);
   U2149 : AOI22_X1 port map( A1 => n18503, A2 => n26742, B1 => n18535, B2 => 
                           n26624, ZN => n26139);
   U2150 : AOI22_X1 port map( A1 => n18599, A2 => n26735, B1 => n18567, B2 => 
                           n26675, ZN => n26138);
   U2151 : AOI22_X1 port map( A1 => n18376, A2 => n26703, B1 => n18439, B2 => 
                           n26734, ZN => n26137);
   U2152 : NAND4_X1 port map( A1 => n26140, A2 => n26139, A3 => n26138, A4 => 
                           n26137, ZN => n26146);
   U2153 : AOI22_X1 port map( A1 => n18758, A2 => n26742, B1 => n18726, B2 => 
                           n19397, ZN => n26144);
   U2154 : AOI22_X1 port map( A1 => n18822, A2 => n26761, B1 => n18854, B2 => 
                           n18368, ZN => n26143);
   U2155 : AOI22_X1 port map( A1 => n18662, A2 => n26680, B1 => n18630, B2 => 
                           n26703, ZN => n26142);
   U2156 : AOI22_X1 port map( A1 => n18694, A2 => n19399, B1 => n18790, B2 => 
                           n19395, ZN => n26141);
   U2157 : NAND4_X1 port map( A1 => n26144, A2 => n26143, A3 => n26142, A4 => 
                           n26141, ZN => n26145);
   U2158 : AOI22_X1 port map( A1 => n26523, A2 => n26146, B1 => n26748, B2 => 
                           n26145, ZN => n26147);
   U2159 : OAI21_X1 port map( B1 => n26689, B2 => n26148, A => n26147, ZN => 
                           OUT1(26));
   U2160 : AOI22_X1 port map( A1 => n19143, A2 => n18308, B1 => n19335, B2 => 
                           n18297, ZN => n26152);
   U2161 : CLKBUF_X1 port map( A => n18296, Z => n26638);
   U2162 : AOI22_X1 port map( A1 => n18919, A2 => n26638, B1 => n19111, B2 => 
                           n26637, ZN => n26151);
   U2163 : AOI22_X1 port map( A1 => n18951, A2 => n18301, B1 => n19367, B2 => 
                           n26695, ZN => n26150);
   U2164 : AOI22_X1 port map( A1 => n19207, A2 => n18305, B1 => n19175, B2 => 
                           n26717, ZN => n26149);
   U2165 : NAND4_X1 port map( A1 => n26152, A2 => n26151, A3 => n26150, A4 => 
                           n26149, ZN => n26158);
   U2166 : AOI22_X1 port map( A1 => n19271, A2 => n26665, B1 => n19047, B2 => 
                           n18304, ZN => n26156);
   U2167 : AOI22_X1 port map( A1 => n18983, A2 => n18302, B1 => n18887, B2 => 
                           n26696, ZN => n26155);
   U2168 : AOI22_X1 port map( A1 => n19303, A2 => n18294, B1 => n19239, B2 => 
                           n26727, ZN => n26154);
   U2169 : AOI22_X1 port map( A1 => n19015, A2 => n18307, B1 => n19079, B2 => 
                           n26718, ZN => n26153);
   U2170 : NAND4_X1 port map( A1 => n26156, A2 => n26155, A3 => n26154, A4 => 
                           n26153, ZN => n26157);
   U2171 : NOR2_X1 port map( A1 => n26158, A2 => n26157, ZN => n26170);
   U2172 : AOI22_X1 port map( A1 => n18568, A2 => n26761, B1 => n18377, B2 => 
                           n18292, ZN => n26162);
   U2173 : AOI22_X1 port map( A1 => n18504, A2 => n26674, B1 => n18472, B2 => 
                           n19397, ZN => n26161);
   U2174 : AOI22_X1 port map( A1 => n18440, A2 => n26734, B1 => n18408, B2 => 
                           n18363, ZN => n26160);
   U2175 : AOI22_X1 port map( A1 => n18536, A2 => n18367, B1 => n18600, B2 => 
                           n19398, ZN => n26159);
   U2176 : NAND4_X1 port map( A1 => n26162, A2 => n26161, A3 => n26160, A4 => 
                           n26159, ZN => n26168);
   U2177 : AOI22_X1 port map( A1 => n18855, A2 => n18368, B1 => n18823, B2 => 
                           n26675, ZN => n26166);
   U2178 : AOI22_X1 port map( A1 => n18727, A2 => n26737, B1 => n18631, B2 => 
                           n19400, ZN => n26165);
   U2179 : AOI22_X1 port map( A1 => n18759, A2 => n26674, B1 => n18663, B2 => 
                           n19396, ZN => n26164);
   U2180 : AOI22_X1 port map( A1 => n18695, A2 => n19399, B1 => n18791, B2 => 
                           n26624, ZN => n26163);
   U2181 : NAND4_X1 port map( A1 => n26166, A2 => n26165, A3 => n26164, A4 => 
                           n26163, ZN => n26167);
   U2182 : AOI22_X1 port map( A1 => n26523, A2 => n26168, B1 => n26748, B2 => 
                           n26167, ZN => n26169);
   U2183 : OAI21_X1 port map( B1 => n26689, B2 => n26170, A => n26169, ZN => 
                           OUT1(25));
   U2184 : AOI22_X1 port map( A1 => n19304, A2 => n18294, B1 => n19048, B2 => 
                           n26666, ZN => n26174);
   U2185 : AOI22_X1 port map( A1 => n19240, A2 => n18295, B1 => n19272, B2 => 
                           n18300, ZN => n26173);
   U2186 : AOI22_X1 port map( A1 => n19176, A2 => n18293, B1 => n18888, B2 => 
                           n18306, ZN => n26172);
   U2187 : AOI22_X1 port map( A1 => n19368, A2 => n26695, B1 => n19016, B2 => 
                           n26725, ZN => n26171);
   U2188 : NAND4_X1 port map( A1 => n26174, A2 => n26173, A3 => n26172, A4 => 
                           n26171, ZN => n26180);
   U2189 : AOI22_X1 port map( A1 => n19112, A2 => n18303, B1 => n19336, B2 => 
                           n26720, ZN => n26178);
   U2190 : AOI22_X1 port map( A1 => n19144, A2 => n18308, B1 => n19208, B2 => 
                           n26719, ZN => n26177);
   U2191 : AOI22_X1 port map( A1 => n19080, A2 => n26718, B1 => n18952, B2 => 
                           n26716, ZN => n26176);
   U2192 : AOI22_X1 port map( A1 => n18984, A2 => n18302, B1 => n18920, B2 => 
                           n26638, ZN => n26175);
   U2193 : NAND4_X1 port map( A1 => n26178, A2 => n26177, A3 => n26176, A4 => 
                           n26175, ZN => n26179);
   U2194 : NOR2_X1 port map( A1 => n26180, A2 => n26179, ZN => n26192);
   U2195 : AOI22_X1 port map( A1 => n18505, A2 => n26674, B1 => n18601, B2 => 
                           n18368, ZN => n26184);
   U2196 : AOI22_X1 port map( A1 => n18441, A2 => n26734, B1 => n18409, B2 => 
                           n19396, ZN => n26183);
   U2197 : AOI22_X1 port map( A1 => n18473, A2 => n18364, B1 => n18569, B2 => 
                           n26736, ZN => n26182);
   U2198 : AOI22_X1 port map( A1 => n19394, A2 => n26703, B1 => n18537, B2 => 
                           n18367, ZN => n26181);
   U2199 : NAND4_X1 port map( A1 => n26184, A2 => n26183, A3 => n26182, A4 => 
                           n26181, ZN => n26190);
   U2200 : AOI22_X1 port map( A1 => n18760, A2 => n26760, B1 => n18824, B2 => 
                           n26736, ZN => n26188);
   U2201 : AOI22_X1 port map( A1 => n18792, A2 => n26624, B1 => n18856, B2 => 
                           n26735, ZN => n26187);
   U2202 : AOI22_X1 port map( A1 => n18696, A2 => n18290, B1 => n18632, B2 => 
                           n26703, ZN => n26186);
   U2203 : AOI22_X1 port map( A1 => n18728, A2 => n19397, B1 => n18664, B2 => 
                           n26680, ZN => n26185);
   U2204 : NAND4_X1 port map( A1 => n26188, A2 => n26187, A3 => n26186, A4 => 
                           n26185, ZN => n26189);
   U2205 : AOI22_X1 port map( A1 => n26523, A2 => n26190, B1 => n26256, B2 => 
                           n26189, ZN => n26191);
   U2206 : OAI21_X1 port map( B1 => n26689, B2 => n26192, A => n26191, ZN => 
                           OUT1(24));
   U2207 : AOI22_X1 port map( A1 => n19145, A2 => n18308, B1 => n19017, B2 => 
                           n18307, ZN => n26196);
   U2208 : AOI22_X1 port map( A1 => n19081, A2 => n18298, B1 => n19209, B2 => 
                           n18305, ZN => n26195);
   U2209 : AOI22_X1 port map( A1 => n18889, A2 => n26696, B1 => n18953, B2 => 
                           n18301, ZN => n26194);
   U2210 : AOI22_X1 port map( A1 => n18985, A2 => n26667, B1 => n19305, B2 => 
                           n18294, ZN => n26193);
   U2211 : NAND4_X1 port map( A1 => n26196, A2 => n26195, A3 => n26194, A4 => 
                           n26193, ZN => n26202);
   U2212 : AOI22_X1 port map( A1 => n19337, A2 => n26720, B1 => n19049, B2 => 
                           n18304, ZN => n26200);
   U2213 : AOI22_X1 port map( A1 => n19241, A2 => n26727, B1 => n18921, B2 => 
                           n18296, ZN => n26199);
   U2214 : AOI22_X1 port map( A1 => n19177, A2 => n18293, B1 => n19113, B2 => 
                           n26637, ZN => n26198);
   U2215 : AOI22_X1 port map( A1 => n19369, A2 => n26695, B1 => n19273, B2 => 
                           n18300, ZN => n26197);
   U2216 : NAND4_X1 port map( A1 => n26200, A2 => n26199, A3 => n26198, A4 => 
                           n26197, ZN => n26201);
   U2217 : NOR2_X1 port map( A1 => n26202, A2 => n26201, ZN => n26214);
   U2218 : AOI22_X1 port map( A1 => n18410, A2 => n19396, B1 => n18506, B2 => 
                           n26674, ZN => n26206);
   U2219 : AOI22_X1 port map( A1 => n18378, A2 => n19400, B1 => n18538, B2 => 
                           n19395, ZN => n26205);
   U2220 : AOI22_X1 port map( A1 => n18570, A2 => n26761, B1 => n18442, B2 => 
                           n19399, ZN => n26204);
   U2221 : AOI22_X1 port map( A1 => n18474, A2 => n26737, B1 => n18602, B2 => 
                           n19398, ZN => n26203);
   U2222 : NAND4_X1 port map( A1 => n26206, A2 => n26205, A3 => n26204, A4 => 
                           n26203, ZN => n26212);
   U2223 : AOI22_X1 port map( A1 => n18665, A2 => n19396, B1 => n18793, B2 => 
                           n18367, ZN => n26210);
   U2224 : AOI22_X1 port map( A1 => n18825, A2 => n26761, B1 => n18729, B2 => 
                           n19397, ZN => n26209);
   U2225 : AOI22_X1 port map( A1 => n18761, A2 => n26760, B1 => n18697, B2 => 
                           n26734, ZN => n26208);
   U2226 : AOI22_X1 port map( A1 => n18857, A2 => n26735, B1 => n18633, B2 => 
                           n19400, ZN => n26207);
   U2227 : NAND4_X1 port map( A1 => n26210, A2 => n26209, A3 => n26208, A4 => 
                           n26207, ZN => n26211);
   U2228 : AOI22_X1 port map( A1 => n26523, A2 => n26212, B1 => n26256, B2 => 
                           n26211, ZN => n26213);
   U2229 : OAI21_X1 port map( B1 => n26753, B2 => n26214, A => n26213, ZN => 
                           OUT1(23));
   U2230 : AOI22_X1 port map( A1 => n19370, A2 => n26695, B1 => n19178, B2 => 
                           n18293, ZN => n26218);
   U2231 : AOI22_X1 port map( A1 => n19018, A2 => n18307, B1 => n18890, B2 => 
                           n26696, ZN => n26217);
   U2232 : AOI22_X1 port map( A1 => n19338, A2 => n18297, B1 => n19114, B2 => 
                           n26637, ZN => n26216);
   U2233 : AOI22_X1 port map( A1 => n19210, A2 => n18305, B1 => n18922, B2 => 
                           n18296, ZN => n26215);
   U2234 : NAND4_X1 port map( A1 => n26218, A2 => n26217, A3 => n26216, A4 => 
                           n26215, ZN => n26224);
   U2235 : AOI22_X1 port map( A1 => n19274, A2 => n18300, B1 => n18954, B2 => 
                           n26716, ZN => n26222);
   U2236 : AOI22_X1 port map( A1 => n19306, A2 => n26726, B1 => n19082, B2 => 
                           n18298, ZN => n26221);
   U2237 : AOI22_X1 port map( A1 => n18986, A2 => n26667, B1 => n19050, B2 => 
                           n26666, ZN => n26220);
   U2238 : AOI22_X1 port map( A1 => n19242, A2 => n18295, B1 => n19146, B2 => 
                           n26694, ZN => n26219);
   U2239 : NAND4_X1 port map( A1 => n26222, A2 => n26221, A3 => n26220, A4 => 
                           n26219, ZN => n26223);
   U2240 : NOR2_X1 port map( A1 => n26224, A2 => n26223, ZN => n26236);
   U2241 : AOI22_X1 port map( A1 => n18475, A2 => n18364, B1 => n18411, B2 => 
                           n18363, ZN => n26228);
   U2242 : AOI22_X1 port map( A1 => n18603, A2 => n18368, B1 => n18443, B2 => 
                           n19399, ZN => n26227);
   U2243 : AOI22_X1 port map( A1 => n18539, A2 => n26624, B1 => n18571, B2 => 
                           n26675, ZN => n26226);
   U2244 : AOI22_X1 port map( A1 => n18507, A2 => n26760, B1 => n18379, B2 => 
                           n18292, ZN => n26225);
   U2245 : NAND4_X1 port map( A1 => n26228, A2 => n26227, A3 => n26226, A4 => 
                           n26225, ZN => n26234);
   U2246 : AOI22_X1 port map( A1 => n18762, A2 => n26760, B1 => n18730, B2 => 
                           n18364, ZN => n26232);
   U2247 : AOI22_X1 port map( A1 => n18634, A2 => n19400, B1 => n18858, B2 => 
                           n18368, ZN => n26231);
   U2248 : AOI22_X1 port map( A1 => n18826, A2 => n26761, B1 => n18794, B2 => 
                           n18367, ZN => n26230);
   U2249 : AOI22_X1 port map( A1 => n18698, A2 => n19399, B1 => n18666, B2 => 
                           n19396, ZN => n26229);
   U2250 : NAND4_X1 port map( A1 => n26232, A2 => n26231, A3 => n26230, A4 => 
                           n26229, ZN => n26233);
   U2251 : AOI22_X1 port map( A1 => n26523, A2 => n26234, B1 => n26256, B2 => 
                           n26233, ZN => n26235);
   U2252 : OAI21_X1 port map( B1 => n26753, B2 => n26236, A => n26235, ZN => 
                           OUT1(22));
   U2253 : AOI22_X1 port map( A1 => n19051, A2 => n18304, B1 => n19019, B2 => 
                           n26725, ZN => n26240);
   U2254 : AOI22_X1 port map( A1 => n19211, A2 => n18305, B1 => n19179, B2 => 
                           n18293, ZN => n26239);
   U2255 : AOI22_X1 port map( A1 => n19371, A2 => n18299, B1 => n18923, B2 => 
                           n18296, ZN => n26238);
   U2256 : AOI22_X1 port map( A1 => n19339, A2 => n18297, B1 => n18891, B2 => 
                           n18306, ZN => n26237);
   U2257 : NAND4_X1 port map( A1 => n26240, A2 => n26239, A3 => n26238, A4 => 
                           n26237, ZN => n26246);
   U2258 : AOI22_X1 port map( A1 => n19147, A2 => n26694, B1 => n19115, B2 => 
                           n18303, ZN => n26244);
   U2259 : AOI22_X1 port map( A1 => n19083, A2 => n26718, B1 => n19275, B2 => 
                           n26665, ZN => n26243);
   U2260 : AOI22_X1 port map( A1 => n19307, A2 => n26726, B1 => n19243, B2 => 
                           n26727, ZN => n26242);
   U2261 : AOI22_X1 port map( A1 => n18987, A2 => n18302, B1 => n18955, B2 => 
                           n18301, ZN => n26241);
   U2262 : NAND4_X1 port map( A1 => n26244, A2 => n26243, A3 => n26242, A4 => 
                           n26241, ZN => n26245);
   U2263 : NOR2_X1 port map( A1 => n26246, A2 => n26245, ZN => n26259);
   U2264 : AOI22_X1 port map( A1 => n18540, A2 => n18367, B1 => n18380, B2 => 
                           n26703, ZN => n26250);
   U2265 : AOI22_X1 port map( A1 => n18476, A2 => n19397, B1 => n18444, B2 => 
                           n18290, ZN => n26249);
   U2266 : AOI22_X1 port map( A1 => n18572, A2 => n26761, B1 => n18508, B2 => 
                           n26674, ZN => n26248);
   U2267 : AOI22_X1 port map( A1 => n18604, A2 => n19398, B1 => n18412, B2 => 
                           n18363, ZN => n26247);
   U2268 : NAND4_X1 port map( A1 => n26250, A2 => n26249, A3 => n26248, A4 => 
                           n26247, ZN => n26257);
   U2269 : AOI22_X1 port map( A1 => n18699, A2 => n19399, B1 => n18667, B2 => 
                           n26680, ZN => n26254);
   U2270 : AOI22_X1 port map( A1 => n18795, A2 => n18367, B1 => n18763, B2 => 
                           n26674, ZN => n26253);
   U2271 : AOI22_X1 port map( A1 => n18635, A2 => n19400, B1 => n18859, B2 => 
                           n19398, ZN => n26252);
   U2272 : AOI22_X1 port map( A1 => n18827, A2 => n26761, B1 => n18731, B2 => 
                           n19397, ZN => n26251);
   U2273 : NAND4_X1 port map( A1 => n26254, A2 => n26253, A3 => n26252, A4 => 
                           n26251, ZN => n26255);
   U2274 : AOI22_X1 port map( A1 => n26523, A2 => n26257, B1 => n26256, B2 => 
                           n26255, ZN => n26258);
   U2275 : OAI21_X1 port map( B1 => n26753, B2 => n26259, A => n26258, ZN => 
                           OUT1(21));
   U2276 : AOI22_X1 port map( A1 => n18892, A2 => n26696, B1 => n19084, B2 => 
                           n26718, ZN => n26263);
   U2277 : AOI22_X1 port map( A1 => n19020, A2 => n18307, B1 => n19116, B2 => 
                           n18303, ZN => n26262);
   U2278 : AOI22_X1 port map( A1 => n19052, A2 => n18304, B1 => n19148, B2 => 
                           n26694, ZN => n26261);
   U2279 : AOI22_X1 port map( A1 => n19308, A2 => n18294, B1 => n18988, B2 => 
                           n26667, ZN => n26260);
   U2280 : NAND4_X1 port map( A1 => n26263, A2 => n26262, A3 => n26261, A4 => 
                           n26260, ZN => n26269);
   U2281 : AOI22_X1 port map( A1 => n19180, A2 => n18293, B1 => n19212, B2 => 
                           n26719, ZN => n26267);
   U2282 : AOI22_X1 port map( A1 => n19340, A2 => n26720, B1 => n18956, B2 => 
                           n18301, ZN => n26266);
   U2283 : AOI22_X1 port map( A1 => n19372, A2 => n18299, B1 => n19244, B2 => 
                           n18295, ZN => n26265);
   U2284 : AOI22_X1 port map( A1 => n18924, A2 => n26638, B1 => n19276, B2 => 
                           n26665, ZN => n26264);
   U2285 : NAND4_X1 port map( A1 => n26267, A2 => n26266, A3 => n26265, A4 => 
                           n26264, ZN => n26268);
   U2286 : NOR2_X1 port map( A1 => n26269, A2 => n26268, ZN => n26281);
   U2287 : AOI22_X1 port map( A1 => n18605, A2 => n18368, B1 => n18509, B2 => 
                           n26674, ZN => n26273);
   U2288 : AOI22_X1 port map( A1 => n18541, A2 => n26624, B1 => n18573, B2 => 
                           n26736, ZN => n26272);
   U2289 : AOI22_X1 port map( A1 => n18445, A2 => n18290, B1 => n18381, B2 => 
                           n18292, ZN => n26271);
   U2290 : AOI22_X1 port map( A1 => n18413, A2 => n18363, B1 => n18477, B2 => 
                           n18364, ZN => n26270);
   U2291 : NAND4_X1 port map( A1 => n26273, A2 => n26272, A3 => n26271, A4 => 
                           n26270, ZN => n26279);
   U2292 : AOI22_X1 port map( A1 => n18732, A2 => n26737, B1 => n18764, B2 => 
                           n26674, ZN => n26277);
   U2293 : AOI22_X1 port map( A1 => n18668, A2 => n26680, B1 => n18796, B2 => 
                           n26624, ZN => n26276);
   U2294 : AOI22_X1 port map( A1 => n18828, A2 => n26761, B1 => n18636, B2 => 
                           n26703, ZN => n26275);
   U2295 : AOI22_X1 port map( A1 => n18700, A2 => n18290, B1 => n18860, B2 => 
                           n18368, ZN => n26274);
   U2296 : NAND4_X1 port map( A1 => n26277, A2 => n26276, A3 => n26275, A4 => 
                           n26274, ZN => n26278);
   U2297 : AOI22_X1 port map( A1 => n26523, A2 => n26279, B1 => n26748, B2 => 
                           n26278, ZN => n26280);
   U2298 : OAI21_X1 port map( B1 => n26753, B2 => n26281, A => n26280, ZN => 
                           OUT1(20));
   U2299 : AOI22_X1 port map( A1 => n19021, A2 => n26725, B1 => n18925, B2 => 
                           n26638, ZN => n26285);
   U2300 : AOI22_X1 port map( A1 => n19213, A2 => n26719, B1 => n19277, B2 => 
                           n18300, ZN => n26284);
   U2301 : AOI22_X1 port map( A1 => n19181, A2 => n26717, B1 => n19053, B2 => 
                           n18304, ZN => n26283);
   U2302 : AOI22_X1 port map( A1 => n18893, A2 => n18306, B1 => n19149, B2 => 
                           n18308, ZN => n26282);
   U2303 : NAND4_X1 port map( A1 => n26285, A2 => n26284, A3 => n26283, A4 => 
                           n26282, ZN => n26291);
   U2304 : AOI22_X1 port map( A1 => n19085, A2 => n18298, B1 => n19373, B2 => 
                           n18299, ZN => n26289);
   U2305 : AOI22_X1 port map( A1 => n18989, A2 => n26667, B1 => n19245, B2 => 
                           n18295, ZN => n26288);
   U2306 : AOI22_X1 port map( A1 => n19117, A2 => n18303, B1 => n19309, B2 => 
                           n18294, ZN => n26287);
   U2307 : AOI22_X1 port map( A1 => n19341, A2 => n18297, B1 => n18957, B2 => 
                           n18301, ZN => n26286);
   U2308 : NAND4_X1 port map( A1 => n26289, A2 => n26288, A3 => n26287, A4 => 
                           n26286, ZN => n26290);
   U2309 : NOR2_X1 port map( A1 => n26291, A2 => n26290, ZN => n26303);
   U2310 : AOI22_X1 port map( A1 => n18414, A2 => n26680, B1 => n18510, B2 => 
                           n26674, ZN => n26295);
   U2311 : AOI22_X1 port map( A1 => n18542, A2 => n26624, B1 => n18446, B2 => 
                           n26734, ZN => n26294);
   U2312 : AOI22_X1 port map( A1 => n18382, A2 => n18292, B1 => n18606, B2 => 
                           n26735, ZN => n26293);
   U2313 : AOI22_X1 port map( A1 => n18574, A2 => n26761, B1 => n18478, B2 => 
                           n19397, ZN => n26292);
   U2314 : NAND4_X1 port map( A1 => n26295, A2 => n26294, A3 => n26293, A4 => 
                           n26292, ZN => n26301);
   U2315 : AOI22_X1 port map( A1 => n18637, A2 => n19400, B1 => n18733, B2 => 
                           n18364, ZN => n26299);
   U2316 : AOI22_X1 port map( A1 => n18765, A2 => n26742, B1 => n18829, B2 => 
                           n26736, ZN => n26298);
   U2317 : AOI22_X1 port map( A1 => n18797, A2 => n18367, B1 => n18861, B2 => 
                           n18368, ZN => n26297);
   U2318 : AOI22_X1 port map( A1 => n18669, A2 => n18363, B1 => n18701, B2 => 
                           n18290, ZN => n26296);
   U2319 : NAND4_X1 port map( A1 => n26299, A2 => n26298, A3 => n26297, A4 => 
                           n26296, ZN => n26300);
   U2320 : AOI22_X1 port map( A1 => n26523, A2 => n26301, B1 => n26748, B2 => 
                           n26300, ZN => n26302);
   U2321 : OAI21_X1 port map( B1 => n26753, B2 => n26303, A => n26302, ZN => 
                           OUT1(19));
   U2322 : AOI22_X1 port map( A1 => n18926, A2 => n26638, B1 => n19118, B2 => 
                           n18303, ZN => n26307);
   U2323 : AOI22_X1 port map( A1 => n18894, A2 => n18306, B1 => n19310, B2 => 
                           n18294, ZN => n26306);
   U2324 : AOI22_X1 port map( A1 => n18958, A2 => n26716, B1 => n19054, B2 => 
                           n26666, ZN => n26305);
   U2325 : AOI22_X1 port map( A1 => n19022, A2 => n18307, B1 => n19214, B2 => 
                           n18305, ZN => n26304);
   U2326 : NAND4_X1 port map( A1 => n26307, A2 => n26306, A3 => n26305, A4 => 
                           n26304, ZN => n26313);
   U2327 : AOI22_X1 port map( A1 => n19374, A2 => n26695, B1 => n19342, B2 => 
                           n18297, ZN => n26311);
   U2328 : AOI22_X1 port map( A1 => n19246, A2 => n26727, B1 => n19086, B2 => 
                           n18298, ZN => n26310);
   U2329 : AOI22_X1 port map( A1 => n19182, A2 => n26717, B1 => n19278, B2 => 
                           n18300, ZN => n26309);
   U2330 : AOI22_X1 port map( A1 => n19150, A2 => n26694, B1 => n18990, B2 => 
                           n18302, ZN => n26308);
   U2331 : NAND4_X1 port map( A1 => n26311, A2 => n26310, A3 => n26309, A4 => 
                           n26308, ZN => n26312);
   U2332 : NOR2_X1 port map( A1 => n26313, A2 => n26312, ZN => n26325);
   U2333 : AOI22_X1 port map( A1 => n18511, A2 => n26760, B1 => n18575, B2 => 
                           n26736, ZN => n26317);
   U2334 : AOI22_X1 port map( A1 => n18415, A2 => n19396, B1 => n18447, B2 => 
                           n26734, ZN => n26316);
   U2335 : AOI22_X1 port map( A1 => n18479, A2 => n19397, B1 => n18543, B2 => 
                           n19395, ZN => n26315);
   U2336 : AOI22_X1 port map( A1 => n18607, A2 => n26735, B1 => n18383, B2 => 
                           n18292, ZN => n26314);
   U2337 : NAND4_X1 port map( A1 => n26317, A2 => n26316, A3 => n26315, A4 => 
                           n26314, ZN => n26323);
   U2338 : AOI22_X1 port map( A1 => n18638, A2 => n18292, B1 => n18670, B2 => 
                           n18363, ZN => n26321);
   U2339 : AOI22_X1 port map( A1 => n18830, A2 => n26761, B1 => n18734, B2 => 
                           n26737, ZN => n26320);
   U2340 : AOI22_X1 port map( A1 => n18862, A2 => n19398, B1 => n18798, B2 => 
                           n26624, ZN => n26319);
   U2341 : AOI22_X1 port map( A1 => n18766, A2 => n26760, B1 => n18702, B2 => 
                           n19399, ZN => n26318);
   U2342 : NAND4_X1 port map( A1 => n26321, A2 => n26320, A3 => n26319, A4 => 
                           n26318, ZN => n26322);
   U2343 : AOI22_X1 port map( A1 => n26523, A2 => n26323, B1 => n26748, B2 => 
                           n26322, ZN => n26324);
   U2344 : OAI21_X1 port map( B1 => n26753, B2 => n26325, A => n26324, ZN => 
                           OUT1(18));
   U2345 : AOI22_X1 port map( A1 => n19151, A2 => n18308, B1 => n19375, B2 => 
                           n18299, ZN => n26329);
   U2346 : AOI22_X1 port map( A1 => n19183, A2 => n18293, B1 => n19279, B2 => 
                           n18300, ZN => n26328);
   U2347 : AOI22_X1 port map( A1 => n19215, A2 => n18305, B1 => n19311, B2 => 
                           n26726, ZN => n26327);
   U2348 : AOI22_X1 port map( A1 => n19055, A2 => n18304, B1 => n19087, B2 => 
                           n26718, ZN => n26326);
   U2349 : NAND4_X1 port map( A1 => n26329, A2 => n26328, A3 => n26327, A4 => 
                           n26326, ZN => n26335);
   U2350 : AOI22_X1 port map( A1 => n19247, A2 => n18295, B1 => n19343, B2 => 
                           n18297, ZN => n26333);
   U2351 : AOI22_X1 port map( A1 => n18959, A2 => n26716, B1 => n18895, B2 => 
                           n26696, ZN => n26332);
   U2352 : AOI22_X1 port map( A1 => n18991, A2 => n18302, B1 => n19119, B2 => 
                           n26637, ZN => n26331);
   U2353 : AOI22_X1 port map( A1 => n18927, A2 => n18296, B1 => n19023, B2 => 
                           n18307, ZN => n26330);
   U2354 : NAND4_X1 port map( A1 => n26333, A2 => n26332, A3 => n26331, A4 => 
                           n26330, ZN => n26334);
   U2355 : NOR2_X1 port map( A1 => n26335, A2 => n26334, ZN => n26347);
   U2356 : AOI22_X1 port map( A1 => n18384, A2 => n18292, B1 => n18448, B2 => 
                           n18290, ZN => n26339);
   U2357 : AOI22_X1 port map( A1 => n18416, A2 => n19396, B1 => n18512, B2 => 
                           n26674, ZN => n26338);
   U2358 : AOI22_X1 port map( A1 => n18544, A2 => n18367, B1 => n18576, B2 => 
                           n26736, ZN => n26337);
   U2359 : AOI22_X1 port map( A1 => n19393, A2 => n19398, B1 => n18480, B2 => 
                           n18364, ZN => n26336);
   U2360 : NAND4_X1 port map( A1 => n26339, A2 => n26338, A3 => n26337, A4 => 
                           n26336, ZN => n26345);
   U2361 : AOI22_X1 port map( A1 => n18735, A2 => n18364, B1 => n18767, B2 => 
                           n26674, ZN => n26343);
   U2362 : AOI22_X1 port map( A1 => n18831, A2 => n26761, B1 => n18703, B2 => 
                           n19399, ZN => n26342);
   U2363 : AOI22_X1 port map( A1 => n18799, A2 => n19395, B1 => n18639, B2 => 
                           n18292, ZN => n26341);
   U2364 : AOI22_X1 port map( A1 => n18671, A2 => n19396, B1 => n18863, B2 => 
                           n18368, ZN => n26340);
   U2365 : NAND4_X1 port map( A1 => n26343, A2 => n26342, A3 => n26341, A4 => 
                           n26340, ZN => n26344);
   U2366 : AOI22_X1 port map( A1 => n26523, A2 => n26345, B1 => n26748, B2 => 
                           n26344, ZN => n26346);
   U2367 : OAI21_X1 port map( B1 => n26753, B2 => n26347, A => n26346, ZN => 
                           OUT1(17));
   U2368 : AOI22_X1 port map( A1 => n18960, A2 => n26716, B1 => n19024, B2 => 
                           n26725, ZN => n26351);
   U2369 : AOI22_X1 port map( A1 => n19344, A2 => n26720, B1 => n19152, B2 => 
                           n18308, ZN => n26350);
   U2370 : AOI22_X1 port map( A1 => n18896, A2 => n18306, B1 => n19280, B2 => 
                           n26665, ZN => n26349);
   U2371 : AOI22_X1 port map( A1 => n19312, A2 => n18294, B1 => n19216, B2 => 
                           n26719, ZN => n26348);
   U2372 : NAND4_X1 port map( A1 => n26351, A2 => n26350, A3 => n26349, A4 => 
                           n26348, ZN => n26357);
   U2373 : AOI22_X1 port map( A1 => n19248, A2 => n26727, B1 => n18992, B2 => 
                           n18302, ZN => n26355);
   U2374 : AOI22_X1 port map( A1 => n19120, A2 => n18303, B1 => n19056, B2 => 
                           n18304, ZN => n26354);
   U2375 : AOI22_X1 port map( A1 => n19184, A2 => n18293, B1 => n18928, B2 => 
                           n26638, ZN => n26353);
   U2376 : AOI22_X1 port map( A1 => n19376, A2 => n18299, B1 => n19088, B2 => 
                           n18298, ZN => n26352);
   U2377 : NAND4_X1 port map( A1 => n26355, A2 => n26354, A3 => n26353, A4 => 
                           n26352, ZN => n26356);
   U2378 : NOR2_X1 port map( A1 => n26357, A2 => n26356, ZN => n26369);
   U2379 : CLKBUF_X1 port map( A => n26478, Z => n26750);
   U2380 : AOI22_X1 port map( A1 => n18545, A2 => n19395, B1 => n18385, B2 => 
                           n19400, ZN => n26361);
   U2381 : AOI22_X1 port map( A1 => n18577, A2 => n26761, B1 => n18417, B2 => 
                           n18363, ZN => n26360);
   U2382 : AOI22_X1 port map( A1 => n18608, A2 => n18368, B1 => n18513, B2 => 
                           n26674, ZN => n26359);
   U2383 : AOI22_X1 port map( A1 => n18449, A2 => n19399, B1 => n18481, B2 => 
                           n19397, ZN => n26358);
   U2384 : NAND4_X1 port map( A1 => n26361, A2 => n26360, A3 => n26359, A4 => 
                           n26358, ZN => n26367);
   U2385 : AOI22_X1 port map( A1 => n18736, A2 => n18364, B1 => n18672, B2 => 
                           n19396, ZN => n26365);
   U2386 : AOI22_X1 port map( A1 => n18640, A2 => n18292, B1 => n18800, B2 => 
                           n18367, ZN => n26364);
   U2387 : AOI22_X1 port map( A1 => n18768, A2 => n26760, B1 => n18704, B2 => 
                           n18290, ZN => n26363);
   U2388 : AOI22_X1 port map( A1 => n18864, A2 => n18368, B1 => n18832, B2 => 
                           n26675, ZN => n26362);
   U2389 : NAND4_X1 port map( A1 => n26365, A2 => n26364, A3 => n26363, A4 => 
                           n26362, ZN => n26366);
   U2390 : AOI22_X1 port map( A1 => n26750, A2 => n26367, B1 => n26748, B2 => 
                           n26366, ZN => n26368);
   U2391 : OAI21_X1 port map( B1 => n26753, B2 => n26369, A => n26368, ZN => 
                           OUT1(16));
   U2392 : AOI22_X1 port map( A1 => n19057, A2 => n26666, B1 => n18993, B2 => 
                           n18302, ZN => n26373);
   U2393 : AOI22_X1 port map( A1 => n19217, A2 => n18305, B1 => n18929, B2 => 
                           n18296, ZN => n26372);
   U2394 : AOI22_X1 port map( A1 => n19025, A2 => n18307, B1 => n19281, B2 => 
                           n18300, ZN => n26371);
   U2395 : AOI22_X1 port map( A1 => n19377, A2 => n18299, B1 => n19089, B2 => 
                           n18298, ZN => n26370);
   U2396 : NAND4_X1 port map( A1 => n26373, A2 => n26372, A3 => n26371, A4 => 
                           n26370, ZN => n26379);
   U2397 : AOI22_X1 port map( A1 => n19313, A2 => n18294, B1 => n18961, B2 => 
                           n18301, ZN => n26377);
   U2398 : AOI22_X1 port map( A1 => n19185, A2 => n18293, B1 => n19121, B2 => 
                           n18303, ZN => n26376);
   U2399 : AOI22_X1 port map( A1 => n19345, A2 => n18297, B1 => n19153, B2 => 
                           n18308, ZN => n26375);
   U2400 : AOI22_X1 port map( A1 => n19249, A2 => n26727, B1 => n18897, B2 => 
                           n18306, ZN => n26374);
   U2401 : NAND4_X1 port map( A1 => n26377, A2 => n26376, A3 => n26375, A4 => 
                           n26374, ZN => n26378);
   U2402 : NOR2_X1 port map( A1 => n26379, A2 => n26378, ZN => n26391);
   U2403 : AOI22_X1 port map( A1 => n18546, A2 => n18367, B1 => n18609, B2 => 
                           n26735, ZN => n26383);
   U2404 : AOI22_X1 port map( A1 => n18418, A2 => n26680, B1 => n18386, B2 => 
                           n26703, ZN => n26382);
   U2405 : AOI22_X1 port map( A1 => n18450, A2 => n26734, B1 => n18482, B2 => 
                           n26737, ZN => n26381);
   U2406 : AOI22_X1 port map( A1 => n18514, A2 => n26742, B1 => n18578, B2 => 
                           n26675, ZN => n26380);
   U2407 : NAND4_X1 port map( A1 => n26383, A2 => n26382, A3 => n26381, A4 => 
                           n26380, ZN => n26389);
   U2408 : AOI22_X1 port map( A1 => n18769, A2 => n26742, B1 => n18641, B2 => 
                           n18292, ZN => n26387);
   U2409 : AOI22_X1 port map( A1 => n18833, A2 => n26761, B1 => n18865, B2 => 
                           n18368, ZN => n26386);
   U2410 : AOI22_X1 port map( A1 => n18673, A2 => n26680, B1 => n18801, B2 => 
                           n18367, ZN => n26385);
   U2411 : AOI22_X1 port map( A1 => n18737, A2 => n19397, B1 => n18705, B2 => 
                           n19399, ZN => n26384);
   U2412 : NAND4_X1 port map( A1 => n26387, A2 => n26386, A3 => n26385, A4 => 
                           n26384, ZN => n26388);
   U2413 : AOI22_X1 port map( A1 => n26478, A2 => n26389, B1 => n26748, B2 => 
                           n26388, ZN => n26390);
   U2414 : OAI21_X1 port map( B1 => n26753, B2 => n26391, A => n26390, ZN => 
                           OUT1(15));
   U2415 : AOI22_X1 port map( A1 => n19026, A2 => n18307, B1 => n19186, B2 => 
                           n18293, ZN => n26395);
   U2416 : AOI22_X1 port map( A1 => n19314, A2 => n26726, B1 => n19346, B2 => 
                           n18297, ZN => n26394);
   U2417 : AOI22_X1 port map( A1 => n19122, A2 => n26637, B1 => n18994, B2 => 
                           n26667, ZN => n26393);
   U2418 : AOI22_X1 port map( A1 => n19218, A2 => n18305, B1 => n19378, B2 => 
                           n18299, ZN => n26392);
   U2419 : NAND4_X1 port map( A1 => n26395, A2 => n26394, A3 => n26393, A4 => 
                           n26392, ZN => n26401);
   U2420 : AOI22_X1 port map( A1 => n18962, A2 => n18301, B1 => n19154, B2 => 
                           n26694, ZN => n26399);
   U2421 : AOI22_X1 port map( A1 => n18930, A2 => n26638, B1 => n19058, B2 => 
                           n26666, ZN => n26398);
   U2422 : AOI22_X1 port map( A1 => n19250, A2 => n26727, B1 => n19282, B2 => 
                           n26665, ZN => n26397);
   U2423 : AOI22_X1 port map( A1 => n19090, A2 => n26718, B1 => n18898, B2 => 
                           n18306, ZN => n26396);
   U2424 : NAND4_X1 port map( A1 => n26399, A2 => n26398, A3 => n26397, A4 => 
                           n26396, ZN => n26400);
   U2425 : NOR2_X1 port map( A1 => n26401, A2 => n26400, ZN => n26413);
   U2426 : AOI22_X1 port map( A1 => n18515, A2 => n26760, B1 => n18387, B2 => 
                           n26703, ZN => n26405);
   U2427 : AOI22_X1 port map( A1 => n18483, A2 => n26737, B1 => n18419, B2 => 
                           n26680, ZN => n26404);
   U2428 : AOI22_X1 port map( A1 => n18579, A2 => n26761, B1 => n18610, B2 => 
                           n26735, ZN => n26403);
   U2429 : AOI22_X1 port map( A1 => n18451, A2 => n18290, B1 => n18547, B2 => 
                           n18367, ZN => n26402);
   U2430 : NAND4_X1 port map( A1 => n26405, A2 => n26404, A3 => n26403, A4 => 
                           n26402, ZN => n26411);
   U2431 : AOI22_X1 port map( A1 => n18706, A2 => n18290, B1 => n18642, B2 => 
                           n18292, ZN => n26409);
   U2432 : AOI22_X1 port map( A1 => n18770, A2 => n26760, B1 => n18802, B2 => 
                           n26624, ZN => n26408);
   U2433 : AOI22_X1 port map( A1 => n18674, A2 => n26680, B1 => n18834, B2 => 
                           n26736, ZN => n26407);
   U2434 : AOI22_X1 port map( A1 => n18738, A2 => n26737, B1 => n18866, B2 => 
                           n26735, ZN => n26406);
   U2435 : NAND4_X1 port map( A1 => n26409, A2 => n26408, A3 => n26407, A4 => 
                           n26406, ZN => n26410);
   U2436 : AOI22_X1 port map( A1 => n26523, A2 => n26411, B1 => n26748, B2 => 
                           n26410, ZN => n26412);
   U2437 : OAI21_X1 port map( B1 => n26753, B2 => n26413, A => n26412, ZN => 
                           OUT1(14));
   U2438 : AOI22_X1 port map( A1 => n19059, A2 => n18304, B1 => n19315, B2 => 
                           n26726, ZN => n26417);
   U2439 : AOI22_X1 port map( A1 => n19091, A2 => n18298, B1 => n18899, B2 => 
                           n18306, ZN => n26416);
   U2440 : AOI22_X1 port map( A1 => n18995, A2 => n26667, B1 => n19155, B2 => 
                           n18308, ZN => n26415);
   U2441 : AOI22_X1 port map( A1 => n19283, A2 => n26665, B1 => n18931, B2 => 
                           n18296, ZN => n26414);
   U2442 : NAND4_X1 port map( A1 => n26417, A2 => n26416, A3 => n26415, A4 => 
                           n26414, ZN => n26423);
   U2443 : AOI22_X1 port map( A1 => n19187, A2 => n26717, B1 => n19027, B2 => 
                           n18307, ZN => n26421);
   U2444 : AOI22_X1 port map( A1 => n19379, A2 => n18299, B1 => n19251, B2 => 
                           n18295, ZN => n26420);
   U2445 : AOI22_X1 port map( A1 => n19347, A2 => n26720, B1 => n19219, B2 => 
                           n18305, ZN => n26419);
   U2446 : AOI22_X1 port map( A1 => n18963, A2 => n18301, B1 => n19123, B2 => 
                           n18303, ZN => n26418);
   U2447 : NAND4_X1 port map( A1 => n26421, A2 => n26420, A3 => n26419, A4 => 
                           n26418, ZN => n26422);
   U2448 : NOR2_X1 port map( A1 => n26423, A2 => n26422, ZN => n26435);
   U2449 : AOI22_X1 port map( A1 => n18452, A2 => n19399, B1 => n18484, B2 => 
                           n18364, ZN => n26427);
   U2450 : AOI22_X1 port map( A1 => n18580, A2 => n26761, B1 => n18516, B2 => 
                           n26674, ZN => n26426);
   U2451 : AOI22_X1 port map( A1 => n18388, A2 => n19400, B1 => n18611, B2 => 
                           n19398, ZN => n26425);
   U2452 : AOI22_X1 port map( A1 => n18548, A2 => n26624, B1 => n18420, B2 => 
                           n18363, ZN => n26424);
   U2453 : NAND4_X1 port map( A1 => n26427, A2 => n26426, A3 => n26425, A4 => 
                           n26424, ZN => n26433);
   U2454 : AOI22_X1 port map( A1 => n18771, A2 => n26760, B1 => n18643, B2 => 
                           n26703, ZN => n26431);
   U2455 : AOI22_X1 port map( A1 => n18835, A2 => n26761, B1 => n18707, B2 => 
                           n18290, ZN => n26430);
   U2456 : AOI22_X1 port map( A1 => n18739, A2 => n26737, B1 => n18675, B2 => 
                           n26680, ZN => n26429);
   U2457 : AOI22_X1 port map( A1 => n18803, A2 => n19395, B1 => n18867, B2 => 
                           n19398, ZN => n26428);
   U2458 : NAND4_X1 port map( A1 => n26431, A2 => n26430, A3 => n26429, A4 => 
                           n26428, ZN => n26432);
   U2459 : AOI22_X1 port map( A1 => n26750, A2 => n26433, B1 => n26748, B2 => 
                           n26432, ZN => n26434);
   U2460 : OAI21_X1 port map( B1 => n26753, B2 => n26435, A => n26434, ZN => 
                           OUT1(13));
   U2461 : AOI22_X1 port map( A1 => n18964, A2 => n18301, B1 => n19060, B2 => 
                           n18304, ZN => n26439);
   U2462 : AOI22_X1 port map( A1 => n19220, A2 => n26719, B1 => n18996, B2 => 
                           n18302, ZN => n26438);
   U2463 : AOI22_X1 port map( A1 => n19380, A2 => n26695, B1 => n19284, B2 => 
                           n18300, ZN => n26437);
   U2464 : AOI22_X1 port map( A1 => n19316, A2 => n18294, B1 => n18932, B2 => 
                           n18296, ZN => n26436);
   U2465 : NAND4_X1 port map( A1 => n26439, A2 => n26438, A3 => n26437, A4 => 
                           n26436, ZN => n26445);
   U2466 : AOI22_X1 port map( A1 => n19156, A2 => n18308, B1 => n18900, B2 => 
                           n18306, ZN => n26443);
   U2467 : AOI22_X1 port map( A1 => n19348, A2 => n18297, B1 => n19092, B2 => 
                           n18298, ZN => n26442);
   U2468 : AOI22_X1 port map( A1 => n19028, A2 => n26725, B1 => n19124, B2 => 
                           n18303, ZN => n26441);
   U2469 : AOI22_X1 port map( A1 => n19188, A2 => n18293, B1 => n19252, B2 => 
                           n18295, ZN => n26440);
   U2470 : NAND4_X1 port map( A1 => n26443, A2 => n26442, A3 => n26441, A4 => 
                           n26440, ZN => n26444);
   U2471 : NOR2_X1 port map( A1 => n26445, A2 => n26444, ZN => n26457);
   U2472 : AOI22_X1 port map( A1 => n18517, A2 => n26760, B1 => n18549, B2 => 
                           n26624, ZN => n26449);
   U2473 : AOI22_X1 port map( A1 => n18421, A2 => n26680, B1 => n18453, B2 => 
                           n26734, ZN => n26448);
   U2474 : AOI22_X1 port map( A1 => n18389, A2 => n26703, B1 => n18612, B2 => 
                           n18368, ZN => n26447);
   U2475 : AOI22_X1 port map( A1 => n18581, A2 => n26761, B1 => n18485, B2 => 
                           n19397, ZN => n26446);
   U2476 : NAND4_X1 port map( A1 => n26449, A2 => n26448, A3 => n26447, A4 => 
                           n26446, ZN => n26455);
   U2477 : AOI22_X1 port map( A1 => n18708, A2 => n18290, B1 => n18676, B2 => 
                           n26680, ZN => n26453);
   U2478 : AOI22_X1 port map( A1 => n18644, A2 => n19400, B1 => n18772, B2 => 
                           n26674, ZN => n26452);
   U2479 : AOI22_X1 port map( A1 => n18836, A2 => n26761, B1 => n18868, B2 => 
                           n19398, ZN => n26451);
   U2480 : AOI22_X1 port map( A1 => n18740, A2 => n18364, B1 => n18804, B2 => 
                           n18367, ZN => n26450);
   U2481 : NAND4_X1 port map( A1 => n26453, A2 => n26452, A3 => n26451, A4 => 
                           n26450, ZN => n26454);
   U2482 : AOI22_X1 port map( A1 => n26523, A2 => n26455, B1 => n26748, B2 => 
                           n26454, ZN => n26456);
   U2483 : OAI21_X1 port map( B1 => n26753, B2 => n26457, A => n26456, ZN => 
                           OUT1(12));
   U2484 : AOI22_X1 port map( A1 => n18901, A2 => n26696, B1 => n19349, B2 => 
                           n18297, ZN => n26461);
   U2485 : AOI22_X1 port map( A1 => n19157, A2 => n18308, B1 => n18997, B2 => 
                           n18302, ZN => n26460);
   U2486 : AOI22_X1 port map( A1 => n19125, A2 => n26637, B1 => n19093, B2 => 
                           n18298, ZN => n26459);
   U2487 : AOI22_X1 port map( A1 => n19061, A2 => n26666, B1 => n19253, B2 => 
                           n18295, ZN => n26458);
   U2488 : NAND4_X1 port map( A1 => n26461, A2 => n26460, A3 => n26459, A4 => 
                           n26458, ZN => n26467);
   U2489 : AOI22_X1 port map( A1 => n19285, A2 => n26665, B1 => n19381, B2 => 
                           n18299, ZN => n26465);
   U2490 : AOI22_X1 port map( A1 => n19029, A2 => n26725, B1 => n18965, B2 => 
                           n26716, ZN => n26464);
   U2491 : AOI22_X1 port map( A1 => n19189, A2 => n18293, B1 => n18933, B2 => 
                           n26638, ZN => n26463);
   U2492 : AOI22_X1 port map( A1 => n19221, A2 => n26719, B1 => n19317, B2 => 
                           n18294, ZN => n26462);
   U2493 : NAND4_X1 port map( A1 => n26465, A2 => n26464, A3 => n26463, A4 => 
                           n26462, ZN => n26466);
   U2494 : NOR2_X1 port map( A1 => n26467, A2 => n26466, ZN => n26480);
   U2495 : AOI22_X1 port map( A1 => n18486, A2 => n18364, B1 => n18454, B2 => 
                           n26734, ZN => n26471);
   U2496 : AOI22_X1 port map( A1 => n18518, A2 => n26760, B1 => n18582, B2 => 
                           n26736, ZN => n26470);
   U2497 : AOI22_X1 port map( A1 => n18550, A2 => n18367, B1 => n18422, B2 => 
                           n19396, ZN => n26469);
   U2498 : AOI22_X1 port map( A1 => n18613, A2 => n26735, B1 => n18390, B2 => 
                           n18292, ZN => n26468);
   U2499 : NAND4_X1 port map( A1 => n26471, A2 => n26470, A3 => n26469, A4 => 
                           n26468, ZN => n26477);
   U2500 : AOI22_X1 port map( A1 => n18869, A2 => n26735, B1 => n18645, B2 => 
                           n18292, ZN => n26475);
   U2501 : AOI22_X1 port map( A1 => n18773, A2 => n26760, B1 => n18741, B2 => 
                           n19397, ZN => n26474);
   U2502 : AOI22_X1 port map( A1 => n18837, A2 => n26736, B1 => n18805, B2 => 
                           n19395, ZN => n26473);
   U2503 : AOI22_X1 port map( A1 => n18677, A2 => n19396, B1 => n18709, B2 => 
                           n18290, ZN => n26472);
   U2504 : NAND4_X1 port map( A1 => n26475, A2 => n26474, A3 => n26473, A4 => 
                           n26472, ZN => n26476);
   U2505 : AOI22_X1 port map( A1 => n26478, A2 => n26477, B1 => n26748, B2 => 
                           n26476, ZN => n26479);
   U2506 : OAI21_X1 port map( B1 => n26753, B2 => n26480, A => n26479, ZN => 
                           OUT1(11));
   U2507 : AOI22_X1 port map( A1 => n19286, A2 => n26665, B1 => n18998, B2 => 
                           n18302, ZN => n26484);
   U2508 : AOI22_X1 port map( A1 => n19318, A2 => n18294, B1 => n19254, B2 => 
                           n18295, ZN => n26483);
   U2509 : AOI22_X1 port map( A1 => n19158, A2 => n26694, B1 => n19350, B2 => 
                           n26720, ZN => n26482);
   U2510 : AOI22_X1 port map( A1 => n19222, A2 => n18305, B1 => n19094, B2 => 
                           n26718, ZN => n26481);
   U2511 : NAND4_X1 port map( A1 => n26484, A2 => n26483, A3 => n26482, A4 => 
                           n26481, ZN => n26490);
   U2512 : AOI22_X1 port map( A1 => n19382, A2 => n26695, B1 => n19126, B2 => 
                           n26637, ZN => n26488);
   U2513 : AOI22_X1 port map( A1 => n19062, A2 => n18304, B1 => n18902, B2 => 
                           n26696, ZN => n26487);
   U2514 : AOI22_X1 port map( A1 => n19190, A2 => n26717, B1 => n18966, B2 => 
                           n18301, ZN => n26486);
   U2515 : AOI22_X1 port map( A1 => n18934, A2 => n26638, B1 => n19030, B2 => 
                           n18307, ZN => n26485);
   U2516 : NAND4_X1 port map( A1 => n26488, A2 => n26487, A3 => n26486, A4 => 
                           n26485, ZN => n26489);
   U2517 : NOR2_X1 port map( A1 => n26490, A2 => n26489, ZN => n26502);
   U2518 : AOI22_X1 port map( A1 => n18487, A2 => n18364, B1 => n18423, B2 => 
                           n18363, ZN => n26494);
   U2519 : AOI22_X1 port map( A1 => n18519, A2 => n26760, B1 => n18391, B2 => 
                           n18292, ZN => n26493);
   U2520 : AOI22_X1 port map( A1 => n18455, A2 => n26734, B1 => n18583, B2 => 
                           n26675, ZN => n26492);
   U2521 : AOI22_X1 port map( A1 => n18551, A2 => n19395, B1 => n18614, B2 => 
                           n26735, ZN => n26491);
   U2522 : NAND4_X1 port map( A1 => n26494, A2 => n26493, A3 => n26492, A4 => 
                           n26491, ZN => n26500);
   U2523 : AOI22_X1 port map( A1 => n18774, A2 => n26760, B1 => n18870, B2 => 
                           n26735, ZN => n26498);
   U2524 : AOI22_X1 port map( A1 => n18710, A2 => n26734, B1 => n18742, B2 => 
                           n26737, ZN => n26497);
   U2525 : AOI22_X1 port map( A1 => n18838, A2 => n26675, B1 => n18678, B2 => 
                           n18363, ZN => n26496);
   U2526 : AOI22_X1 port map( A1 => n18806, A2 => n18367, B1 => n18646, B2 => 
                           n18292, ZN => n26495);
   U2527 : NAND4_X1 port map( A1 => n26498, A2 => n26497, A3 => n26496, A4 => 
                           n26495, ZN => n26499);
   U2528 : AOI22_X1 port map( A1 => n26523, A2 => n26500, B1 => n26748, B2 => 
                           n26499, ZN => n26501);
   U2529 : OAI21_X1 port map( B1 => n26689, B2 => n26502, A => n26501, ZN => 
                           OUT1(10));
   U2530 : AOI22_X1 port map( A1 => n19191, A2 => n26717, B1 => n18935, B2 => 
                           n18296, ZN => n26506);
   U2531 : AOI22_X1 port map( A1 => n19287, A2 => n18300, B1 => n18967, B2 => 
                           n26716, ZN => n26505);
   U2532 : AOI22_X1 port map( A1 => n18999, A2 => n18302, B1 => n19031, B2 => 
                           n18307, ZN => n26504);
   U2533 : AOI22_X1 port map( A1 => n18903, A2 => n18306, B1 => n19063, B2 => 
                           n18304, ZN => n26503);
   U2534 : NAND4_X1 port map( A1 => n26506, A2 => n26505, A3 => n26504, A4 => 
                           n26503, ZN => n26512);
   U2535 : AOI22_X1 port map( A1 => n19095, A2 => n18298, B1 => n19319, B2 => 
                           n18294, ZN => n26510);
   U2536 : AOI22_X1 port map( A1 => n19383, A2 => n18299, B1 => n19127, B2 => 
                           n26637, ZN => n26509);
   U2537 : AOI22_X1 port map( A1 => n19159, A2 => n18308, B1 => n19255, B2 => 
                           n26727, ZN => n26508);
   U2538 : AOI22_X1 port map( A1 => n19351, A2 => n18297, B1 => n19223, B2 => 
                           n18305, ZN => n26507);
   U2539 : NAND4_X1 port map( A1 => n26510, A2 => n26509, A3 => n26508, A4 => 
                           n26507, ZN => n26511);
   U2540 : NOR2_X1 port map( A1 => n26512, A2 => n26511, ZN => n26525);
   U2541 : AOI22_X1 port map( A1 => n18456, A2 => n18290, B1 => n18552, B2 => 
                           n18367, ZN => n26516);
   U2542 : AOI22_X1 port map( A1 => n18615, A2 => n18368, B1 => n18424, B2 => 
                           n19396, ZN => n26515);
   U2543 : AOI22_X1 port map( A1 => n18488, A2 => n19397, B1 => n18584, B2 => 
                           n26736, ZN => n26514);
   U2544 : AOI22_X1 port map( A1 => n18520, A2 => n26760, B1 => n18392, B2 => 
                           n26703, ZN => n26513);
   U2545 : NAND4_X1 port map( A1 => n26516, A2 => n26515, A3 => n26514, A4 => 
                           n26513, ZN => n26522);
   U2546 : AOI22_X1 port map( A1 => n18711, A2 => n18290, B1 => n18807, B2 => 
                           n26624, ZN => n26520);
   U2547 : AOI22_X1 port map( A1 => n18679, A2 => n18363, B1 => n18775, B2 => 
                           n26742, ZN => n26519);
   U2548 : AOI22_X1 port map( A1 => n18743, A2 => n26737, B1 => n18647, B2 => 
                           n18292, ZN => n26518);
   U2549 : AOI22_X1 port map( A1 => n18871, A2 => n19398, B1 => n18839, B2 => 
                           n26736, ZN => n26517);
   U2550 : NAND4_X1 port map( A1 => n26520, A2 => n26519, A3 => n26518, A4 => 
                           n26517, ZN => n26521);
   U2551 : AOI22_X1 port map( A1 => n26523, A2 => n26522, B1 => n26748, B2 => 
                           n26521, ZN => n26524);
   U2552 : OAI21_X1 port map( B1 => n26753, B2 => n26525, A => n26524, ZN => 
                           OUT1(9));
   U2553 : AOI22_X1 port map( A1 => n19352, A2 => n18297, B1 => n19224, B2 => 
                           n18305, ZN => n26529);
   U2554 : AOI22_X1 port map( A1 => n18936, A2 => n18296, B1 => n18904, B2 => 
                           n18306, ZN => n26528);
   U2555 : AOI22_X1 port map( A1 => n19000, A2 => n18302, B1 => n19288, B2 => 
                           n26665, ZN => n26527);
   U2556 : AOI22_X1 port map( A1 => n19128, A2 => n26637, B1 => n19160, B2 => 
                           n18308, ZN => n26526);
   U2557 : NAND4_X1 port map( A1 => n26529, A2 => n26528, A3 => n26527, A4 => 
                           n26526, ZN => n26535);
   U2558 : AOI22_X1 port map( A1 => n19032, A2 => n18307, B1 => n19064, B2 => 
                           n18304, ZN => n26533);
   U2559 : AOI22_X1 port map( A1 => n19192, A2 => n26717, B1 => n19256, B2 => 
                           n26727, ZN => n26532);
   U2560 : AOI22_X1 port map( A1 => n18968, A2 => n26716, B1 => n19320, B2 => 
                           n18294, ZN => n26531);
   U2561 : AOI22_X1 port map( A1 => n19384, A2 => n18299, B1 => n19096, B2 => 
                           n18298, ZN => n26530);
   U2562 : NAND4_X1 port map( A1 => n26533, A2 => n26532, A3 => n26531, A4 => 
                           n26530, ZN => n26534);
   U2563 : NOR2_X1 port map( A1 => n26535, A2 => n26534, ZN => n26547);
   U2564 : AOI22_X1 port map( A1 => n18553, A2 => n26624, B1 => n18521, B2 => 
                           n26742, ZN => n26539);
   U2565 : AOI22_X1 port map( A1 => n18425, A2 => n19396, B1 => n18489, B2 => 
                           n18364, ZN => n26538);
   U2566 : AOI22_X1 port map( A1 => n18457, A2 => n18290, B1 => n18393, B2 => 
                           n26703, ZN => n26537);
   U2567 : AOI22_X1 port map( A1 => n18616, A2 => n26735, B1 => n18585, B2 => 
                           n26675, ZN => n26536);
   U2568 : NAND4_X1 port map( A1 => n26539, A2 => n26538, A3 => n26537, A4 => 
                           n26536, ZN => n26545);
   U2569 : AOI22_X1 port map( A1 => n18712, A2 => n26734, B1 => n18648, B2 => 
                           n18292, ZN => n26543);
   U2570 : AOI22_X1 port map( A1 => n18744, A2 => n18364, B1 => n18872, B2 => 
                           n18368, ZN => n26542);
   U2571 : AOI22_X1 port map( A1 => n18808, A2 => n19395, B1 => n18776, B2 => 
                           n26742, ZN => n26541);
   U2572 : AOI22_X1 port map( A1 => n18840, A2 => n26736, B1 => n18680, B2 => 
                           n26680, ZN => n26540);
   U2573 : NAND4_X1 port map( A1 => n26543, A2 => n26542, A3 => n26541, A4 => 
                           n26540, ZN => n26544);
   U2574 : AOI22_X1 port map( A1 => n26750, A2 => n26545, B1 => n26748, B2 => 
                           n26544, ZN => n26546);
   U2575 : OAI21_X1 port map( B1 => n26753, B2 => n26547, A => n26546, ZN => 
                           OUT1(8));
   U2576 : AOI22_X1 port map( A1 => n19065, A2 => n26666, B1 => n19289, B2 => 
                           n26665, ZN => n26551);
   U2577 : AOI22_X1 port map( A1 => n19097, A2 => n18298, B1 => n19321, B2 => 
                           n26726, ZN => n26550);
   U2578 : AOI22_X1 port map( A1 => n18969, A2 => n18301, B1 => n19001, B2 => 
                           n26667, ZN => n26549);
   U2579 : AOI22_X1 port map( A1 => n19033, A2 => n18307, B1 => n19353, B2 => 
                           n18297, ZN => n26548);
   U2580 : NAND4_X1 port map( A1 => n26551, A2 => n26550, A3 => n26549, A4 => 
                           n26548, ZN => n26557);
   U2581 : AOI22_X1 port map( A1 => n19161, A2 => n18308, B1 => n19129, B2 => 
                           n18303, ZN => n26555);
   U2582 : AOI22_X1 port map( A1 => n19385, A2 => n18299, B1 => n19257, B2 => 
                           n26727, ZN => n26554);
   U2583 : AOI22_X1 port map( A1 => n19193, A2 => n18293, B1 => n19225, B2 => 
                           n18305, ZN => n26553);
   U2584 : AOI22_X1 port map( A1 => n18937, A2 => n18296, B1 => n18905, B2 => 
                           n26696, ZN => n26552);
   U2585 : NAND4_X1 port map( A1 => n26555, A2 => n26554, A3 => n26553, A4 => 
                           n26552, ZN => n26556);
   U2586 : NOR2_X1 port map( A1 => n26557, A2 => n26556, ZN => n26569);
   U2587 : AOI22_X1 port map( A1 => n18554, A2 => n26624, B1 => n18458, B2 => 
                           n26734, ZN => n26561);
   U2588 : AOI22_X1 port map( A1 => n18522, A2 => n26760, B1 => n18490, B2 => 
                           n19397, ZN => n26560);
   U2589 : AOI22_X1 port map( A1 => n18426, A2 => n18363, B1 => n18617, B2 => 
                           n19398, ZN => n26559);
   U2590 : AOI22_X1 port map( A1 => n18394, A2 => n18292, B1 => n18586, B2 => 
                           n26675, ZN => n26558);
   U2591 : NAND4_X1 port map( A1 => n26561, A2 => n26560, A3 => n26559, A4 => 
                           n26558, ZN => n26567);
   U2592 : AOI22_X1 port map( A1 => n18745, A2 => n18364, B1 => n18713, B2 => 
                           n18290, ZN => n26565);
   U2593 : AOI22_X1 port map( A1 => n18681, A2 => n19396, B1 => n18873, B2 => 
                           n19398, ZN => n26564);
   U2594 : AOI22_X1 port map( A1 => n18649, A2 => n26703, B1 => n18809, B2 => 
                           n19395, ZN => n26563);
   U2595 : AOI22_X1 port map( A1 => n18841, A2 => n26736, B1 => n18777, B2 => 
                           n26742, ZN => n26562);
   U2596 : NAND4_X1 port map( A1 => n26565, A2 => n26564, A3 => n26563, A4 => 
                           n26562, ZN => n26566);
   U2597 : AOI22_X1 port map( A1 => n26750, A2 => n26567, B1 => n26748, B2 => 
                           n26566, ZN => n26568);
   U2598 : OAI21_X1 port map( B1 => n26753, B2 => n26569, A => n26568, ZN => 
                           OUT1(7));
   U2599 : AOI22_X1 port map( A1 => n19194, A2 => n18293, B1 => n19322, B2 => 
                           n18294, ZN => n26573);
   U2600 : AOI22_X1 port map( A1 => n19386, A2 => n26695, B1 => n19258, B2 => 
                           n18295, ZN => n26572);
   U2601 : AOI22_X1 port map( A1 => n18938, A2 => n18296, B1 => n19290, B2 => 
                           n18300, ZN => n26571);
   U2602 : AOI22_X1 port map( A1 => n19226, A2 => n18305, B1 => n19130, B2 => 
                           n18303, ZN => n26570);
   U2603 : NAND4_X1 port map( A1 => n26573, A2 => n26572, A3 => n26571, A4 => 
                           n26570, ZN => n26579);
   U2604 : AOI22_X1 port map( A1 => n18970, A2 => n18301, B1 => n19098, B2 => 
                           n26718, ZN => n26577);
   U2605 : AOI22_X1 port map( A1 => n19034, A2 => n18307, B1 => n19162, B2 => 
                           n18308, ZN => n26576);
   U2606 : AOI22_X1 port map( A1 => n19354, A2 => n18297, B1 => n19066, B2 => 
                           n18304, ZN => n26575);
   U2607 : AOI22_X1 port map( A1 => n18906, A2 => n18306, B1 => n19002, B2 => 
                           n26667, ZN => n26574);
   U2608 : NAND4_X1 port map( A1 => n26577, A2 => n26576, A3 => n26575, A4 => 
                           n26574, ZN => n26578);
   U2609 : NOR2_X1 port map( A1 => n26579, A2 => n26578, ZN => n26591);
   U2610 : AOI22_X1 port map( A1 => n18587, A2 => n26736, B1 => n18523, B2 => 
                           n26742, ZN => n26583);
   U2611 : AOI22_X1 port map( A1 => n18427, A2 => n26680, B1 => n18459, B2 => 
                           n19399, ZN => n26582);
   U2612 : AOI22_X1 port map( A1 => n18618, A2 => n26735, B1 => n18395, B2 => 
                           n26703, ZN => n26581);
   U2613 : AOI22_X1 port map( A1 => n18491, A2 => n18364, B1 => n18555, B2 => 
                           n19395, ZN => n26580);
   U2614 : NAND4_X1 port map( A1 => n26583, A2 => n26582, A3 => n26581, A4 => 
                           n26580, ZN => n26589);
   U2615 : AOI22_X1 port map( A1 => n18714, A2 => n18290, B1 => n18874, B2 => 
                           n18368, ZN => n26587);
   U2616 : AOI22_X1 port map( A1 => n18650, A2 => n26703, B1 => n18842, B2 => 
                           n26675, ZN => n26586);
   U2617 : AOI22_X1 port map( A1 => n18746, A2 => n26737, B1 => n18682, B2 => 
                           n18363, ZN => n26585);
   U2618 : AOI22_X1 port map( A1 => n18810, A2 => n26624, B1 => n18778, B2 => 
                           n26742, ZN => n26584);
   U2619 : NAND4_X1 port map( A1 => n26587, A2 => n26586, A3 => n26585, A4 => 
                           n26584, ZN => n26588);
   U2620 : AOI22_X1 port map( A1 => n26750, A2 => n26589, B1 => n26748, B2 => 
                           n26588, ZN => n26590);
   U2621 : OAI21_X1 port map( B1 => n26753, B2 => n26591, A => n26590, ZN => 
                           OUT1(6));
   U2622 : AOI22_X1 port map( A1 => n19387, A2 => n18299, B1 => n19355, B2 => 
                           n26720, ZN => n26595);
   U2623 : AOI22_X1 port map( A1 => n19163, A2 => n18308, B1 => n18907, B2 => 
                           n18306, ZN => n26594);
   U2624 : AOI22_X1 port map( A1 => n18971, A2 => n18301, B1 => n19035, B2 => 
                           n26725, ZN => n26593);
   U2625 : AOI22_X1 port map( A1 => n19227, A2 => n18305, B1 => n19259, B2 => 
                           n18295, ZN => n26592);
   U2626 : NAND4_X1 port map( A1 => n26595, A2 => n26594, A3 => n26593, A4 => 
                           n26592, ZN => n26601);
   U2627 : AOI22_X1 port map( A1 => n19131, A2 => n18303, B1 => n19099, B2 => 
                           n18298, ZN => n26599);
   U2628 : AOI22_X1 port map( A1 => n18939, A2 => n26638, B1 => n19323, B2 => 
                           n18294, ZN => n26598);
   U2629 : AOI22_X1 port map( A1 => n19067, A2 => n18304, B1 => n19003, B2 => 
                           n18302, ZN => n26597);
   U2630 : AOI22_X1 port map( A1 => n19291, A2 => n18300, B1 => n19195, B2 => 
                           n26717, ZN => n26596);
   U2631 : NAND4_X1 port map( A1 => n26599, A2 => n26598, A3 => n26597, A4 => 
                           n26596, ZN => n26600);
   U2632 : NOR2_X1 port map( A1 => n26601, A2 => n26600, ZN => n26613);
   U2633 : AOI22_X1 port map( A1 => n18428, A2 => n19396, B1 => n18588, B2 => 
                           n26675, ZN => n26605);
   U2634 : AOI22_X1 port map( A1 => n18556, A2 => n18367, B1 => n18396, B2 => 
                           n26703, ZN => n26604);
   U2635 : AOI22_X1 port map( A1 => n18492, A2 => n26737, B1 => n18524, B2 => 
                           n26742, ZN => n26603);
   U2636 : AOI22_X1 port map( A1 => n18460, A2 => n18290, B1 => n18619, B2 => 
                           n19398, ZN => n26602);
   U2637 : NAND4_X1 port map( A1 => n26605, A2 => n26604, A3 => n26603, A4 => 
                           n26602, ZN => n26611);
   U2638 : AOI22_X1 port map( A1 => n18811, A2 => n19395, B1 => n18875, B2 => 
                           n26735, ZN => n26609);
   U2639 : AOI22_X1 port map( A1 => n18651, A2 => n19400, B1 => n18715, B2 => 
                           n26734, ZN => n26608);
   U2640 : AOI22_X1 port map( A1 => n18843, A2 => n26761, B1 => n18779, B2 => 
                           n26742, ZN => n26607);
   U2641 : AOI22_X1 port map( A1 => n18683, A2 => n18363, B1 => n18747, B2 => 
                           n18364, ZN => n26606);
   U2642 : NAND4_X1 port map( A1 => n26609, A2 => n26608, A3 => n26607, A4 => 
                           n26606, ZN => n26610);
   U2643 : AOI22_X1 port map( A1 => n26750, A2 => n26611, B1 => n26748, B2 => 
                           n26610, ZN => n26612);
   U2644 : OAI21_X1 port map( B1 => n26689, B2 => n26613, A => n26612, ZN => 
                           OUT1(5));
   U2645 : AOI22_X1 port map( A1 => n19100, A2 => n18298, B1 => n19004, B2 => 
                           n18302, ZN => n26617);
   U2646 : AOI22_X1 port map( A1 => n19164, A2 => n26694, B1 => n19228, B2 => 
                           n26719, ZN => n26616);
   U2647 : AOI22_X1 port map( A1 => n19356, A2 => n26720, B1 => n19324, B2 => 
                           n18294, ZN => n26615);
   U2648 : AOI22_X1 port map( A1 => n18972, A2 => n26716, B1 => n19388, B2 => 
                           n18299, ZN => n26614);
   U2649 : NAND4_X1 port map( A1 => n26617, A2 => n26616, A3 => n26615, A4 => 
                           n26614, ZN => n26623);
   U2650 : AOI22_X1 port map( A1 => n18940, A2 => n26638, B1 => n19292, B2 => 
                           n18300, ZN => n26621);
   U2651 : AOI22_X1 port map( A1 => n18908, A2 => n18306, B1 => n19132, B2 => 
                           n26637, ZN => n26620);
   U2652 : AOI22_X1 port map( A1 => n19036, A2 => n26725, B1 => n19196, B2 => 
                           n26717, ZN => n26619);
   U2653 : AOI22_X1 port map( A1 => n19068, A2 => n18304, B1 => n19260, B2 => 
                           n18295, ZN => n26618);
   U2654 : NAND4_X1 port map( A1 => n26621, A2 => n26620, A3 => n26619, A4 => 
                           n26618, ZN => n26622);
   U2655 : NOR2_X1 port map( A1 => n26623, A2 => n26622, ZN => n26636);
   U2656 : AOI22_X1 port map( A1 => n18589, A2 => n26736, B1 => n18557, B2 => 
                           n26624, ZN => n26628);
   U2657 : AOI22_X1 port map( A1 => n18397, A2 => n19400, B1 => n18493, B2 => 
                           n26737, ZN => n26627);
   U2658 : AOI22_X1 port map( A1 => n18525, A2 => n26760, B1 => n18461, B2 => 
                           n26734, ZN => n26626);
   U2659 : AOI22_X1 port map( A1 => n18429, A2 => n18363, B1 => n18620, B2 => 
                           n18368, ZN => n26625);
   U2660 : NAND4_X1 port map( A1 => n26628, A2 => n26627, A3 => n26626, A4 => 
                           n26625, ZN => n26634);
   U2661 : AOI22_X1 port map( A1 => n18812, A2 => n19395, B1 => n18652, B2 => 
                           n19400, ZN => n26632);
   U2662 : AOI22_X1 port map( A1 => n18876, A2 => n19398, B1 => n18748, B2 => 
                           n18364, ZN => n26631);
   U2663 : AOI22_X1 port map( A1 => n18780, A2 => n26760, B1 => n18716, B2 => 
                           n18290, ZN => n26630);
   U2664 : AOI22_X1 port map( A1 => n18844, A2 => n26736, B1 => n18684, B2 => 
                           n19396, ZN => n26629);
   U2665 : NAND4_X1 port map( A1 => n26632, A2 => n26631, A3 => n26630, A4 => 
                           n26629, ZN => n26633);
   U2666 : AOI22_X1 port map( A1 => n26750, A2 => n26634, B1 => n26748, B2 => 
                           n26633, ZN => n26635);
   U2667 : OAI21_X1 port map( B1 => n26753, B2 => n26636, A => n26635, ZN => 
                           OUT1(4));
   U2668 : AOI22_X1 port map( A1 => n19325, A2 => n18294, B1 => n19357, B2 => 
                           n18297, ZN => n26642);
   U2669 : AOI22_X1 port map( A1 => n19037, A2 => n18307, B1 => n19005, B2 => 
                           n18302, ZN => n26641);
   U2670 : AOI22_X1 port map( A1 => n18973, A2 => n26716, B1 => n19133, B2 => 
                           n26637, ZN => n26640);
   U2671 : AOI22_X1 port map( A1 => n18941, A2 => n26638, B1 => n19197, B2 => 
                           n18293, ZN => n26639);
   U2672 : NAND4_X1 port map( A1 => n26642, A2 => n26641, A3 => n26640, A4 => 
                           n26639, ZN => n26648);
   U2673 : AOI22_X1 port map( A1 => n19229, A2 => n26719, B1 => n18909, B2 => 
                           n26696, ZN => n26646);
   U2674 : AOI22_X1 port map( A1 => n19101, A2 => n26718, B1 => n19293, B2 => 
                           n18300, ZN => n26645);
   U2675 : AOI22_X1 port map( A1 => n19261, A2 => n18295, B1 => n19069, B2 => 
                           n26666, ZN => n26644);
   U2676 : AOI22_X1 port map( A1 => n19389, A2 => n18299, B1 => n19165, B2 => 
                           n26694, ZN => n26643);
   U2677 : NAND4_X1 port map( A1 => n26646, A2 => n26645, A3 => n26644, A4 => 
                           n26643, ZN => n26647);
   U2678 : NOR2_X1 port map( A1 => n26648, A2 => n26647, ZN => n26660);
   U2679 : AOI22_X1 port map( A1 => n18621, A2 => n18368, B1 => n18558, B2 => 
                           n19395, ZN => n26652);
   U2680 : AOI22_X1 port map( A1 => n18398, A2 => n19400, B1 => n18590, B2 => 
                           n26675, ZN => n26651);
   U2681 : AOI22_X1 port map( A1 => n18430, A2 => n26680, B1 => n18462, B2 => 
                           n19399, ZN => n26650);
   U2682 : AOI22_X1 port map( A1 => n18494, A2 => n19397, B1 => n18526, B2 => 
                           n26742, ZN => n26649);
   U2683 : NAND4_X1 port map( A1 => n26652, A2 => n26651, A3 => n26650, A4 => 
                           n26649, ZN => n26658);
   U2684 : AOI22_X1 port map( A1 => n18845, A2 => n26736, B1 => n18877, B2 => 
                           n18368, ZN => n26656);
   U2685 : AOI22_X1 port map( A1 => n18717, A2 => n18290, B1 => n18813, B2 => 
                           n18367, ZN => n26655);
   U2686 : AOI22_X1 port map( A1 => n18653, A2 => n19400, B1 => n18749, B2 => 
                           n26737, ZN => n26654);
   U2687 : AOI22_X1 port map( A1 => n18685, A2 => n18363, B1 => n18781, B2 => 
                           n26742, ZN => n26653);
   U2688 : NAND4_X1 port map( A1 => n26656, A2 => n26655, A3 => n26654, A4 => 
                           n26653, ZN => n26657);
   U2689 : AOI22_X1 port map( A1 => n26750, A2 => n26658, B1 => n26748, B2 => 
                           n26657, ZN => n26659);
   U2690 : OAI21_X1 port map( B1 => n26753, B2 => n26660, A => n26659, ZN => 
                           OUT1(3));
   U2691 : AOI22_X1 port map( A1 => n18942, A2 => n18296, B1 => n19230, B2 => 
                           n18305, ZN => n26664);
   U2692 : AOI22_X1 port map( A1 => n19262, A2 => n18295, B1 => n18974, B2 => 
                           n18301, ZN => n26663);
   U2693 : AOI22_X1 port map( A1 => n19198, A2 => n18293, B1 => n19390, B2 => 
                           n18299, ZN => n26662);
   U2694 : AOI22_X1 port map( A1 => n18910, A2 => n26696, B1 => n19358, B2 => 
                           n26720, ZN => n26661);
   U2695 : NAND4_X1 port map( A1 => n26664, A2 => n26663, A3 => n26662, A4 => 
                           n26661, ZN => n26673);
   U2696 : AOI22_X1 port map( A1 => n19326, A2 => n26726, B1 => n19294, B2 => 
                           n26665, ZN => n26671);
   U2697 : AOI22_X1 port map( A1 => n19070, A2 => n26666, B1 => n19038, B2 => 
                           n26725, ZN => n26670);
   U2698 : AOI22_X1 port map( A1 => n19166, A2 => n26694, B1 => n19006, B2 => 
                           n26667, ZN => n26669);
   U2699 : AOI22_X1 port map( A1 => n19102, A2 => n18298, B1 => n19134, B2 => 
                           n18303, ZN => n26668);
   U2700 : NAND4_X1 port map( A1 => n26671, A2 => n26670, A3 => n26669, A4 => 
                           n26668, ZN => n26672);
   U2701 : NOR2_X1 port map( A1 => n26673, A2 => n26672, ZN => n26688);
   U2702 : AOI22_X1 port map( A1 => n18463, A2 => n26734, B1 => n18622, B2 => 
                           n26735, ZN => n26679);
   U2703 : AOI22_X1 port map( A1 => n18527, A2 => n26674, B1 => n18399, B2 => 
                           n18292, ZN => n26678);
   U2704 : AOI22_X1 port map( A1 => n18559, A2 => n18367, B1 => n18591, B2 => 
                           n26675, ZN => n26677);
   U2705 : AOI22_X1 port map( A1 => n18431, A2 => n18363, B1 => n18495, B2 => 
                           n18364, ZN => n26676);
   U2706 : NAND4_X1 port map( A1 => n26679, A2 => n26678, A3 => n26677, A4 => 
                           n26676, ZN => n26686);
   U2707 : AOI22_X1 port map( A1 => n18654, A2 => n19400, B1 => n18718, B2 => 
                           n26734, ZN => n26684);
   U2708 : AOI22_X1 port map( A1 => n18750, A2 => n18364, B1 => n18782, B2 => 
                           n26742, ZN => n26683);
   U2709 : AOI22_X1 port map( A1 => n18878, A2 => n26735, B1 => n18814, B2 => 
                           n19395, ZN => n26682);
   U2710 : AOI22_X1 port map( A1 => n18686, A2 => n26680, B1 => n18846, B2 => 
                           n26736, ZN => n26681);
   U2711 : NAND4_X1 port map( A1 => n26684, A2 => n26683, A3 => n26682, A4 => 
                           n26681, ZN => n26685);
   U2712 : AOI22_X1 port map( A1 => n26750, A2 => n26686, B1 => n26748, B2 => 
                           n26685, ZN => n26687);
   U2713 : OAI21_X1 port map( B1 => n26689, B2 => n26688, A => n26687, ZN => 
                           OUT1(2));
   U2714 : AOI22_X1 port map( A1 => n18975, A2 => n18301, B1 => n19039, B2 => 
                           n18307, ZN => n26693);
   U2715 : AOI22_X1 port map( A1 => n19231, A2 => n18305, B1 => n19199, B2 => 
                           n26717, ZN => n26692);
   U2716 : AOI22_X1 port map( A1 => n19359, A2 => n18297, B1 => n19103, B2 => 
                           n26718, ZN => n26691);
   U2717 : AOI22_X1 port map( A1 => n19007, A2 => n18302, B1 => n19327, B2 => 
                           n26726, ZN => n26690);
   U2718 : NAND4_X1 port map( A1 => n26693, A2 => n26692, A3 => n26691, A4 => 
                           n26690, ZN => n26702);
   U2719 : AOI22_X1 port map( A1 => n19167, A2 => n26694, B1 => n19263, B2 => 
                           n18295, ZN => n26700);
   U2720 : AOI22_X1 port map( A1 => n19071, A2 => n18304, B1 => n19135, B2 => 
                           n18303, ZN => n26699);
   U2721 : AOI22_X1 port map( A1 => n18943, A2 => n18296, B1 => n19391, B2 => 
                           n26695, ZN => n26698);
   U2722 : AOI22_X1 port map( A1 => n18911, A2 => n26696, B1 => n19295, B2 => 
                           n18300, ZN => n26697);
   U2723 : NAND4_X1 port map( A1 => n26700, A2 => n26699, A3 => n26698, A4 => 
                           n26697, ZN => n26701);
   U2724 : NOR2_X1 port map( A1 => n26702, A2 => n26701, ZN => n26715);
   U2725 : AOI22_X1 port map( A1 => n18400, A2 => n26703, B1 => n18623, B2 => 
                           n18368, ZN => n26707);
   U2726 : AOI22_X1 port map( A1 => n18496, A2 => n19397, B1 => n18560, B2 => 
                           n19395, ZN => n26706);
   U2727 : AOI22_X1 port map( A1 => n18528, A2 => n26742, B1 => n18464, B2 => 
                           n19399, ZN => n26705);
   U2728 : AOI22_X1 port map( A1 => n18432, A2 => n18363, B1 => n18592, B2 => 
                           n26736, ZN => n26704);
   U2729 : NAND4_X1 port map( A1 => n26707, A2 => n26706, A3 => n26705, A4 => 
                           n26704, ZN => n26713);
   U2730 : AOI22_X1 port map( A1 => n18815, A2 => n19395, B1 => n18719, B2 => 
                           n26734, ZN => n26711);
   U2731 : AOI22_X1 port map( A1 => n18655, A2 => n18292, B1 => n18783, B2 => 
                           n26760, ZN => n26710);
   U2732 : AOI22_X1 port map( A1 => n18751, A2 => n26737, B1 => n18687, B2 => 
                           n19396, ZN => n26709);
   U2733 : AOI22_X1 port map( A1 => n18847, A2 => n26736, B1 => n18879, B2 => 
                           n18368, ZN => n26708);
   U2734 : NAND4_X1 port map( A1 => n26711, A2 => n26710, A3 => n26709, A4 => 
                           n26708, ZN => n26712);
   U2735 : AOI22_X1 port map( A1 => n26750, A2 => n26713, B1 => n26748, B2 => 
                           n26712, ZN => n26714);
   U2736 : OAI21_X1 port map( B1 => n26753, B2 => n26715, A => n26714, ZN => 
                           OUT1(1));
   U2737 : AOI22_X1 port map( A1 => n18912, A2 => n18306, B1 => n18944, B2 => 
                           n18296, ZN => n26724);
   U2738 : AOI22_X1 port map( A1 => n19200, A2 => n26717, B1 => n18976, B2 => 
                           n26716, ZN => n26723);
   U2739 : AOI22_X1 port map( A1 => n19104, A2 => n26718, B1 => n19296, B2 => 
                           n18300, ZN => n26722);
   U2740 : AOI22_X1 port map( A1 => n19360, A2 => n26720, B1 => n19232, B2 => 
                           n26719, ZN => n26721);
   U2741 : NAND4_X1 port map( A1 => n26724, A2 => n26723, A3 => n26722, A4 => 
                           n26721, ZN => n26733);
   U2742 : AOI22_X1 port map( A1 => n19168, A2 => n18308, B1 => n19040, B2 => 
                           n26725, ZN => n26731);
   U2743 : AOI22_X1 port map( A1 => n19264, A2 => n26727, B1 => n19328, B2 => 
                           n26726, ZN => n26730);
   U2744 : AOI22_X1 port map( A1 => n19136, A2 => n18303, B1 => n19072, B2 => 
                           n18304, ZN => n26729);
   U2745 : AOI22_X1 port map( A1 => n19392, A2 => n18299, B1 => n19008, B2 => 
                           n18302, ZN => n26728);
   U2746 : NAND4_X1 port map( A1 => n26731, A2 => n26730, A3 => n26729, A4 => 
                           n26728, ZN => n26732);
   U2747 : NOR2_X1 port map( A1 => n26733, A2 => n26732, ZN => n26752);
   U2748 : AOI22_X1 port map( A1 => n18529, A2 => n26742, B1 => n18465, B2 => 
                           n26734, ZN => n26741);
   U2749 : AOI22_X1 port map( A1 => n18561, A2 => n19395, B1 => n18433, B2 => 
                           n18363, ZN => n26740);
   U2750 : AOI22_X1 port map( A1 => n18593, A2 => n26736, B1 => n18624, B2 => 
                           n26735, ZN => n26739);
   U2751 : AOI22_X1 port map( A1 => n18497, A2 => n26737, B1 => n18401, B2 => 
                           n19400, ZN => n26738);
   U2752 : NAND4_X1 port map( A1 => n26741, A2 => n26740, A3 => n26739, A4 => 
                           n26738, ZN => n26749);
   U2753 : AOI22_X1 port map( A1 => n18688, A2 => n18363, B1 => n18784, B2 => 
                           n26742, ZN => n26746);
   U2754 : AOI22_X1 port map( A1 => n18752, A2 => n19397, B1 => n18656, B2 => 
                           n18292, ZN => n26745);
   U2755 : AOI22_X1 port map( A1 => n18880, A2 => n19398, B1 => n18720, B2 => 
                           n18290, ZN => n26744);
   U2756 : AOI22_X1 port map( A1 => n18848, A2 => n26761, B1 => n18816, B2 => 
                           n19395, ZN => n26743);
   U2757 : NAND4_X1 port map( A1 => n26746, A2 => n26745, A3 => n26744, A4 => 
                           n26743, ZN => n26747);
   U2758 : AOI22_X1 port map( A1 => n26750, A2 => n26749, B1 => n26748, B2 => 
                           n26747, ZN => n26751);
   U2759 : OAI21_X1 port map( B1 => n26753, B2 => n26752, A => n26751, ZN => 
                           OUT1(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, 
      DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, 
      DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, 
      DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, 
      DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, 
      DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, 
      DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, 
      DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, 
      DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, 
      DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_17_port, curr_instruction_to_cu_i_16_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n151, cu_i_n135, 
      cu_i_N279, cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, 
      cu_i_N273, cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, 
      cu_i_cmd_alu_op_type_0_port, cu_i_cmd_alu_op_type_1_port, 
      cu_i_cmd_alu_op_type_2_port, cu_i_cmd_alu_op_type_3_port, 
      cu_i_cmd_word_3_port, cu_i_cmd_word_6_port, cu_i_cmd_word_8_port, 
      datapath_i_alu_output_val_i_0_port, datapath_i_alu_output_val_i_1_port, 
      datapath_i_alu_output_val_i_2_port, datapath_i_alu_output_val_i_3_port, 
      datapath_i_alu_output_val_i_4_port, datapath_i_alu_output_val_i_5_port, 
      datapath_i_alu_output_val_i_6_port, datapath_i_alu_output_val_i_7_port, 
      datapath_i_alu_output_val_i_8_port, datapath_i_alu_output_val_i_9_port, 
      datapath_i_alu_output_val_i_10_port, datapath_i_alu_output_val_i_11_port,
      datapath_i_alu_output_val_i_12_port, datapath_i_alu_output_val_i_13_port,
      datapath_i_alu_output_val_i_14_port, datapath_i_alu_output_val_i_15_port,
      datapath_i_alu_output_val_i_16_port, datapath_i_alu_output_val_i_17_port,
      datapath_i_alu_output_val_i_18_port, datapath_i_alu_output_val_i_19_port,
      datapath_i_alu_output_val_i_20_port, datapath_i_alu_output_val_i_21_port,
      datapath_i_alu_output_val_i_22_port, datapath_i_alu_output_val_i_23_port,
      datapath_i_alu_output_val_i_24_port, datapath_i_alu_output_val_i_25_port,
      datapath_i_alu_output_val_i_26_port, datapath_i_alu_output_val_i_27_port,
      datapath_i_alu_output_val_i_28_port, datapath_i_alu_output_val_i_29_port,
      datapath_i_alu_output_val_i_30_port, datapath_i_alu_output_val_i_31_port,
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_decode_stage_dp_n44, datapath_i_decode_stage_dp_n43, 
      datapath_i_decode_stage_dp_n42, datapath_i_decode_stage_dp_n41, 
      datapath_i_decode_stage_dp_n40, datapath_i_decode_stage_dp_n39, 
      datapath_i_decode_stage_dp_n38, datapath_i_decode_stage_dp_n37, 
      datapath_i_decode_stage_dp_n36, datapath_i_decode_stage_dp_n35, 
      datapath_i_decode_stage_dp_n34, datapath_i_decode_stage_dp_n33, 
      datapath_i_decode_stage_dp_n32, datapath_i_decode_stage_dp_n31, 
      datapath_i_decode_stage_dp_n30, datapath_i_decode_stage_dp_n29, 
      datapath_i_decode_stage_dp_n28, datapath_i_decode_stage_dp_n27, 
      datapath_i_decode_stage_dp_n26, datapath_i_decode_stage_dp_n25, 
      datapath_i_decode_stage_dp_n24, datapath_i_decode_stage_dp_n23, 
      datapath_i_decode_stage_dp_n22, datapath_i_decode_stage_dp_n21, 
      datapath_i_decode_stage_dp_n20, datapath_i_decode_stage_dp_n19, 
      datapath_i_decode_stage_dp_n18, datapath_i_decode_stage_dp_n17, 
      datapath_i_decode_stage_dp_n16, datapath_i_decode_stage_dp_n15, 
      datapath_i_decode_stage_dp_n14, datapath_i_decode_stage_dp_n13, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, n301, n302, n464, n474, n477, 
      n492, n1302, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1323, n1324, n1325, n1328, n1330, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1350, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1385, n3627, n1388, n3628, n1390, n1393, 
      n1394, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1404, n1405, 
      n1411, n1412, n1413, n1414, n1415, n1422, n1423, n1424, n1425, n1427, 
      n1916, n1429, n1431, n1433, n1435, n1437, n1439, n1441, n1443, n1445, 
      n1447, n1449, n1453, n1458, n1460, n1475, n1477, n1497, n1498, n1500, 
      n1505, n1507, n1510, n1512, n1513, n1518, n1521, n1524, n1527, n1530, 
      n1533, n1536, n1539, n1542, n1545, n1548, n1551, n1554, n1557, n1560, 
      n1563, n1566, n1569, n1572, n1575, n1578, n1581, n1584, n1587, n1590, 
      n1593, n1596, n1599, n1602, n1605, n1608, n1611, n1613, n1614, n1615, 
      n1617, n1619, n1621, n1623, n1625, n1627, n1629, n1631, n1633, n1635, 
      n1637, n1639, n1641, n1643, n1645, n1647, n1649, n1651, n1653, n1655, 
      n1657, n1659, n1661, n1663, n1665, n1667, n1669, n1671, n1673, n1727, 
      n1728, n1758, n1760, n1779, n3629, n1801, n1802, n2299, n2350, n2358, 
      n2359, n2363, n2398, n2416, n2478, n2483, n2485, n2486, n2530, n2547, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
      n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, 
      n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
      n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, 
      n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, 
      n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, 
      n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3158, 
      n3159, n3160, n3161, n3162, IRAM_ADDRESS_1_port, n3164, 
      IRAM_ADDRESS_0_port, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
      n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, 
      n3265, n3266, n3268, n3269, n3271, n3272, n3273, n3275, n3276, n3277, 
      n3278, n3279, n3280, n3281, n3282, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
      n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, 
      n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
      n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, 
      n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, 
      n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, 
      n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, 
      n3510, n3511, n3512, n3513, IRAM_ADDRESS_7_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_9_port, IRAM_ADDRESS_11_port, IRAM_ADDRESS_13_port, 
      IRAM_ADDRESS_15_port, IRAM_ADDRESS_17_port, IRAM_ADDRESS_19_port, 
      IRAM_ADDRESS_21_port, IRAM_ADDRESS_23_port, IRAM_ADDRESS_25_port, 
      IRAM_ADDRESS_27_port, IRAM_ADDRESS_29_port, n3527, n3528, n3529, n3530, 
      n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, 
      n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, 
      n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, 
      IRAM_ADDRESS_6_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3593, n3692, 
      n3596, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, 
      n3643, n3644, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
      n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
      n3664, n3665, n3666, n3667, n3668, n3670, n3671, n3672, n3673, n3674, 
      n3675, n3676, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, 
      n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, 
      n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, 
      n3885, n3886, n3887, n3888, n3889, n3890, n4033, n4034, n4035, n4036, 
      n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
      n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, 
      n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_30_port, n4078, 
      n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, 
      n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
      n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
      n4130, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, 
      n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, 
      n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, 
      n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, 
      n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, 
      n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, 
      n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, 
      n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, 
      n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, 
      n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, 
      n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, 
      n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, 
      n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, 
      n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, 
      n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, 
      n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, 
      n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, 
      n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, 
      n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, 
      n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, 
      n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, 
      n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, 
      n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, 
      n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, 
      n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, 
      n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, 
      n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, 
      n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, 
      n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, 
      n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, 
      n4431, n4432, n4433, n4434, n4435, n_3818, n_3819, n_3820, n_3821, n_3822
      , n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831,
      n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, 
      n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, 
      n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, 
      n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, 
      n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, 
      n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, 
      n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, 
      n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, 
      n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, 
      n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, 
      n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, 
      n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, 
      n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, 
      n_3949, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, 
      n_3958, n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, 
      n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, 
      n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, 
      n_3985, n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, 
      n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, 
      n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, 
      n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, 
      n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, 
      n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, 
      n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, 
      n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, 
      n_4057, n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, 
      n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, 
      n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, 
      n_4084, n_4085, n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, 
      n_4093, n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, 
      n_4102, n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, 
      n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, 
      n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, 
      n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, 
      n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, 
      n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, 
      n_4156, n_4157, n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, 
      n_4165, n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, 
      n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, 
      n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, 
      n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, 
      n_4201, n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, 
      n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, 
      n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, 
      n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, 
      n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, 
      n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, 
      n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, 
      n_4264, n_4265, n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, 
      n_4273, n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, 
      n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, 
      n_4291, n_4292, n_4293, n_4294, n_4295 : std_logic;

begin
   IRAM_ADDRESS <= ( n3692, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => n1513);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => n1512);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_n151);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => n1510);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n4426, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n4430, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n4430, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n4430, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n4430, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n4430, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n4430, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n4430, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n4430, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n4430, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n4430, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n4430, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n3543, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n3543, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n3543, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n3543, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n3543, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n4430, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n4426, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n4426, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n4426, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n4426, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n4426, Z 
                           => DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n4426, Z 
                           => DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n4426, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n4426, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n4426, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n4426, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n4426, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n4426, Z 
                           => DRAM_ADDRESS_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n301, D => n3237, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n4435, D => n3538, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n4435, D => n3537, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n4435, D => n3236, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n301, D => n3238, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n301, D => n3536, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n301, D => n3198, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n301, D => n3199, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n301, D => n3200, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n301, D => n3201, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n301, D => n3202, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n301, D => n3227, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n4435, D => n3231, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n4435, D => n3535, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n4435, D => n3233, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n301, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n301, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n301, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n301, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n301, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n4435, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n301, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n4432, D => n3237, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n4432, D => n3538, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n4057, D => n3537, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n4057, D => n3236, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n4057, D => n3238, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n4057, D => n3536, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n4057, D => n3198, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n4057, D => n3199, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n4057, D => n3200, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n4057, D => n3201, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n4057, D => n3202, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n4057, D => n3227, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n4057, D => n3231, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n4057, D => n3535, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n4057, D => n3233, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n4057, D => n3229, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n4057, D => n3228, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n4432, D => n3232, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n4057, D => n3534, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n4432, D => n3234, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n4057, D => n3230, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n4432, D => n3203, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n4432, D => n3204, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n4057, D => n3205, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n4432, D => n3206, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n4057, D => n3207, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n4432, D => n3207, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n4057, D => n3207, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n4432, D => n3207, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n4057, D => n3207, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n4432, D => n3207, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n4057, D => n3207, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   clk_r_REG6817_S5 : DFFR_X1 port map( D => n1801, CK => CLK, RN => RST, Q => 
                           n_3818, QN => n3593);
   clk_r_REG6665_S5 : DFFR_X1 port map( D => n4046, CK => CLK, RN => RST, Q => 
                           n_3819, QN => n4416);
   clk_r_REG6711_S3 : DFFR_X1 port map( D => n4045, CK => CLK, RN => RST, Q => 
                           DRAM_READNOTWRITE, QN => n_3820);
   clk_r_REG6702_S3 : DFFR_X1 port map( D => n4056, CK => CLK, RN => RST, Q => 
                           n3590, QN => n_3821);
   clk_r_REG6659_S2 : DFFR_X1 port map( D => n3635, CK => CLK, RN => RST, Q => 
                           n3589, QN => n_3822);
   clk_r_REG6655_S1 : DFFR_X1 port map( D => n4053, CK => CLK, RN => RST, Q => 
                           n3588, QN => n4428);
   clk_r_REG6738_S4 : DFFR_X1 port map( D => n3587, CK => CLK, RN => RST, Q => 
                           n3586, QN => n_3823);
   clk_r_REG6734_S3 : DFFR_X1 port map( D => n4037, CK => CLK, RN => RST, Q => 
                           n3585, QN => n_3824);
   clk_r_REG6735_S4 : DFFR_X1 port map( D => n3585, CK => CLK, RN => RST, Q => 
                           n3584, QN => n_3825);
   clk_r_REG6732_S3 : DFFR_X1 port map( D => n4036, CK => CLK, RN => RST, Q => 
                           n3583, QN => n_3826);
   clk_r_REG6733_S4 : DFFR_X1 port map( D => n3583, CK => CLK, RN => RST, Q => 
                           n3582, QN => n_3827);
   clk_r_REG6728_S3 : DFFR_X1 port map( D => n4035, CK => CLK, RN => RST, Q => 
                           n3581, QN => n_3828);
   clk_r_REG6729_S4 : DFFR_X1 port map( D => n3581, CK => CLK, RN => RST, Q => 
                           n3580, QN => n_3829);
   clk_r_REG6726_S3 : DFFR_X1 port map( D => n4034, CK => CLK, RN => RST, Q => 
                           n3579, QN => n_3830);
   clk_r_REG6727_S4 : DFFR_X1 port map( D => n3579, CK => CLK, RN => RST, Q => 
                           n3578, QN => n_3831);
   clk_r_REG6660_S3 : DFFR_X1 port map( D => n4435, CK => CLK, RN => RST, Q => 
                           n3577, QN => n_3832);
   clk_r_REG5002_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_2_port, QN => 
                           n_3833);
   clk_r_REG4856_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_3834);
   clk_r_REG4580_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, CK => 
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_3835);
   clk_r_REG4704_S8 : DFFR_X1 port map( D => n1453, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_6_port, QN => n_3836);
   clk_r_REG4248_S12 : DFFR_X1 port map( D => n1449, CK => CLK, RN => RST, Q =>
                           n_3837, QN => n3655);
   clk_r_REG4010_S15 : DFFR_X1 port map( D => n1447, CK => CLK, RN => RST, Q =>
                           n_3838, QN => n3667);
   clk_r_REG4015_S5 : DFFR_X1 port map( D => n1445, CK => CLK, RN => RST, Q => 
                           n_3839, QN => n3666);
   clk_r_REG4021_S5 : DFFR_X1 port map( D => n1443, CK => CLK, RN => RST, Q => 
                           n_3840, QN => n3668);
   clk_r_REG4027_S12 : DFFR_X1 port map( D => n1441, CK => CLK, RN => RST, Q =>
                           n_3841, QN => n3665);
   clk_r_REG4033_S12 : DFFR_X1 port map( D => n1439, CK => CLK, RN => RST, Q =>
                           n_3842, QN => n3661);
   clk_r_REG4039_S6 : DFFR_X1 port map( D => n1437, CK => CLK, RN => RST, Q => 
                           n_3843, QN => n3656);
   clk_r_REG4583_S5 : DFFR_X1 port map( D => n1435, CK => CLK, RN => RST, Q => 
                           n_3844, QN => n3657);
   clk_r_REG4589_S12 : DFFR_X1 port map( D => n1433, CK => CLK, RN => RST, Q =>
                           n_3845, QN => n3660);
   clk_r_REG4595_S6 : DFFR_X1 port map( D => n1431, CK => CLK, RN => RST, Q => 
                           n_3846, QN => n3663);
   clk_r_REG4601_S12 : DFFR_X1 port map( D => n1429, CK => CLK, RN => RST, Q =>
                           n_3847, QN => n3662);
   clk_r_REG4609_S6 : DFFR_X1 port map( D => n1427, CK => CLK, RN => RST, Q => 
                           n_3848, QN => n3659);
   clk_r_REG6772_S5 : DFFS_X1 port map( D => n1507, CK => CLK, SN => RST, Q => 
                           n3559, QN => n_3849);
   clk_r_REG6777_S3 : DFFS_X1 port map( D => n1802, CK => CLK, SN => RST, Q => 
                           n3558, QN => n_3850);
   clk_r_REG5926_S4 : DFFR_X1 port map( D => n3646, CK => CLK, RN => RST, Q => 
                           n3557, QN => n4419);
   clk_r_REG4661_S17 : DFFR_X1 port map( D => n3652, CK => CLK, RN => RST, Q =>
                           n3556, QN => n_3851);
   clk_r_REG6818_S5 : DFFR_X1 port map( D => n1801, CK => CLK, RN => RST, Q => 
                           n3555, QN => n_3852);
   clk_r_REG5932_S5 : DFFR_X1 port map( D => n3554, CK => CLK, RN => RST, Q => 
                           n3553, QN => n_3853);
   clk_r_REG6788_S5 : DFFS_X1 port map( D => n4047, CK => CLK, SN => RST, Q => 
                           n3552, QN => n_3854);
   clk_r_REG3642_S3 : DFFS_X1 port map( D => n4040, CK => CLK, SN => RST, Q => 
                           n_3855, QN => n3646);
   clk_r_REG4619_S16 : DFFS_X1 port map( D => n4097, CK => CLK, SN => RST, Q =>
                           n3550, QN => n_3856);
   clk_r_REG4620_S17 : DFFS_X1 port map( D => n3550, CK => CLK, SN => RST, Q =>
                           n3549, QN => n_3857);
   clk_r_REG4853_S6 : DFFS_X1 port map( D => n3673, CK => CLK, SN => RST, Q => 
                           n3548, QN => n_3858);
   clk_r_REG4854_S7 : DFFS_X1 port map( D => n3548, CK => CLK, SN => RST, Q => 
                           n3547, QN => n_3859);
   clk_r_REG4999_S6 : DFFS_X1 port map( D => n3672, CK => CLK, SN => RST, Q => 
                           n3546, QN => n_3860);
   clk_r_REG5000_S7 : DFFS_X1 port map( D => n3546, CK => CLK, SN => RST, Q => 
                           n3545, QN => n_3861);
   clk_r_REG6909_S1 : DFFR_X1 port map( D => n4052, CK => CLK, RN => RST, Q => 
                           n3544, QN => n_3862);
   clk_r_REG6707_S3 : DFFS_X1 port map( D => n1760, CK => CLK, SN => RST, Q => 
                           n3543, QN => n_3863);
   clk_r_REG5656_S6 : DFFS_X1 port map( D => n3671, CK => CLK, SN => RST, Q => 
                           n3542, QN => n_3864);
   clk_r_REG5657_S7 : DFFS_X1 port map( D => n3542, CK => CLK, SN => RST, Q => 
                           n3541, QN => n_3865);
   clk_r_REG5924_S6 : DFFS_X1 port map( D => n3676, CK => CLK, SN => RST, Q => 
                           n3540, QN => n_3866);
   clk_r_REG5925_S7 : DFFS_X1 port map( D => n3540, CK => CLK, SN => RST, Q => 
                           n3539, QN => n_3867);
   clk_r_REG6873_S6 : DFFR_X1 port map( D => n4050, CK => CLK, RN => RST, Q => 
                           n3538, QN => n_3868);
   clk_r_REG6871_S6 : DFFR_X1 port map( D => n4051, CK => CLK, RN => RST, Q => 
                           n3537, QN => n_3869);
   clk_r_REG6875_S6 : DFFR_X1 port map( D => n4049, CK => CLK, RN => RST, Q => 
                           n3536, QN => n_3870);
   clk_r_REG6816_S6 : DFFR_X1 port map( D => n4112, CK => CLK, RN => RST, Q => 
                           n3535, QN => n_3871);
   clk_r_REG6815_S6 : DFFR_X1 port map( D => n4113, CK => CLK, RN => RST, Q => 
                           n3534, QN => n_3872);
   clk_r_REG6865_S6 : DFFR_X1 port map( D => n4064, CK => CLK, RN => RST, Q => 
                           n3533, QN => n_3873);
   clk_r_REG6869_S6 : DFFR_X1 port map( D => n4058, CK => CLK, RN => RST, Q => 
                           n3532, QN => n_3874);
   clk_r_REG6868_S6 : DFFR_X1 port map( D => n4061, CK => CLK, RN => RST, Q => 
                           n3531, QN => n_3875);
   clk_r_REG6860_S6 : DFFR_X1 port map( D => n4065, CK => CLK, RN => RST, Q => 
                           n3530, QN => n_3876);
   clk_r_REG6866_S6 : DFFR_X1 port map( D => n4062, CK => CLK, RN => RST, Q => 
                           n3529, QN => n_3877);
   clk_r_REG6910_S1 : DFFR_X1 port map( D => n4063, CK => CLK, RN => RST, Q => 
                           n3528, QN => n_3878);
   clk_r_REG6779_S4 : DFFS_X1 port map( D => n4041, CK => CLK, SN => RST, Q => 
                           n3527, QN => n_3879);
   clk_r_REG4605_S6 : DFFR_X1 port map( D => n4078, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_29_port, QN => n_3880);
   clk_r_REG4599_S6 : DFFR_X1 port map( D => n4079, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_27_port, QN => n_3881);
   clk_r_REG4593_S5 : DFFR_X1 port map( D => n4080, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_25_port, QN => n_3882);
   clk_r_REG4587_S5 : DFFR_X1 port map( D => n4081, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_23_port, QN => n_3883);
   clk_r_REG4043_S5 : DFFR_X1 port map( D => n4086, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_21_port, QN => n_3884);
   clk_r_REG4037_S5 : DFFR_X1 port map( D => n4085, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_19_port, QN => n_3885);
   clk_r_REG4031_S6 : DFFR_X1 port map( D => n4084, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_17_port, QN => n_3886);
   clk_r_REG4025_S5 : DFFR_X1 port map( D => n4082, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_15_port, QN => n_3887);
   clk_r_REG4019_S5 : DFFR_X1 port map( D => n4083, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_13_port, QN => n_3888);
   clk_r_REG4013_S5 : DFFR_X1 port map( D => n4114, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_11_port, QN => n_3889);
   clk_r_REG4242_S5 : DFFR_X1 port map( D => n4115, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_9_port, QN => n_3890);
   clk_r_REG5916_S5 : DFFR_X1 port map( D => n4117, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_5_port, QN => n_3891);
   clk_r_REG4232_S5 : DFFR_X1 port map( D => n4116, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_7_port, QN => n_3892);
   clk_r_REG4621_S16 : DFFS_X1 port map( D => n4096, CK => CLK, SN => RST, Q =>
                           n3513, QN => n_3893);
   clk_r_REG4622_S17 : DFFS_X1 port map( D => n3513, CK => CLK, SN => RST, Q =>
                           n3512, QN => n_3894);
   clk_r_REG4627_S16 : DFFS_X1 port map( D => n4111, CK => CLK, SN => RST, Q =>
                           n3511, QN => n_3895);
   clk_r_REG4628_S17 : DFFS_X1 port map( D => n3511, CK => CLK, SN => RST, Q =>
                           n3510, QN => n_3896);
   clk_r_REG4636_S16 : DFFS_X1 port map( D => n4104, CK => CLK, SN => RST, Q =>
                           n3509, QN => n_3897);
   clk_r_REG4637_S17 : DFFS_X1 port map( D => n3509, CK => CLK, SN => RST, Q =>
                           n3508, QN => n_3898);
   clk_r_REG4642_S16 : DFFS_X1 port map( D => n4103, CK => CLK, SN => RST, Q =>
                           n3507, QN => n_3899);
   clk_r_REG4643_S17 : DFFS_X1 port map( D => n3507, CK => CLK, SN => RST, Q =>
                           n3506, QN => n_3900);
   clk_r_REG4648_S16 : DFFS_X1 port map( D => n4098, CK => CLK, SN => RST, Q =>
                           n3505, QN => n_3901);
   clk_r_REG4649_S17 : DFFS_X1 port map( D => n3505, CK => CLK, SN => RST, Q =>
                           n3504, QN => n_3902);
   clk_r_REG4655_S16 : DFFS_X1 port map( D => n4105, CK => CLK, SN => RST, Q =>
                           n3503, QN => n_3903);
   clk_r_REG4656_S17 : DFFS_X1 port map( D => n3503, CK => CLK, SN => RST, Q =>
                           n3502, QN => n_3904);
   clk_r_REG4663_S16 : DFFS_X1 port map( D => n4099, CK => CLK, SN => RST, Q =>
                           n3501, QN => n_3905);
   clk_r_REG4664_S17 : DFFS_X1 port map( D => n3501, CK => CLK, SN => RST, Q =>
                           n3500, QN => n_3906);
   clk_r_REG4672_S16 : DFFS_X1 port map( D => n4102, CK => CLK, SN => RST, Q =>
                           n3499, QN => n_3907);
   clk_r_REG4673_S17 : DFFS_X1 port map( D => n3499, CK => CLK, SN => RST, Q =>
                           n3498, QN => n_3908);
   clk_r_REG4681_S16 : DFFS_X1 port map( D => n4106, CK => CLK, SN => RST, Q =>
                           n3497, QN => n_3909);
   clk_r_REG4682_S17 : DFFS_X1 port map( D => n3497, CK => CLK, SN => RST, Q =>
                           n3496, QN => n_3910);
   clk_r_REG4690_S16 : DFFS_X1 port map( D => n4100, CK => CLK, SN => RST, Q =>
                           n3495, QN => n_3911);
   clk_r_REG4691_S17 : DFFS_X1 port map( D => n3495, CK => CLK, SN => RST, Q =>
                           n3494, QN => n_3912);
   clk_r_REG4702_S10 : DFFS_X1 port map( D => n4107, CK => CLK, SN => RST, Q =>
                           n3493, QN => n_3913);
   clk_r_REG4703_S11 : DFFS_X1 port map( D => n3493, CK => CLK, SN => RST, Q =>
                           n3492, QN => n_3914);
   clk_r_REG4254_S6 : DFFS_X1 port map( D => n4109, CK => CLK, SN => RST, Q => 
                           n3491, QN => n_3915);
   clk_r_REG4255_S7 : DFFS_X1 port map( D => n3491, CK => CLK, SN => RST, Q => 
                           n3490, QN => n_3916);
   clk_r_REG3647_S6 : DFFS_X1 port map( D => n3675, CK => CLK, SN => RST, Q => 
                           n3489, QN => n_3917);
   clk_r_REG3648_S7 : DFFS_X1 port map( D => n3489, CK => CLK, SN => RST, Q => 
                           n3488, QN => n_3918);
   clk_r_REG4569_S6 : DFFS_X1 port map( D => n3644, CK => CLK, SN => RST, Q => 
                           n3487, QN => n_3919);
   clk_r_REG4570_S7 : DFFS_X1 port map( D => n3487, CK => CLK, SN => RST, Q => 
                           n3486, QN => n_3920);
   clk_r_REG4624_S16 : DFFS_X1 port map( D => n4119, CK => CLK, SN => RST, Q =>
                           n3485, QN => n3647);
   clk_r_REG4625_S17 : DFFR_X1 port map( D => n3647, CK => CLK, RN => RST, Q =>
                           n_3921, QN => n3484);
   clk_r_REG4632_S16 : DFFS_X1 port map( D => n4120, CK => CLK, SN => RST, Q =>
                           n3483, QN => n3648);
   clk_r_REG4633_S17 : DFFR_X1 port map( D => n3648, CK => CLK, RN => RST, Q =>
                           n_3922, QN => n3482);
   clk_r_REG4639_S16 : DFFS_X1 port map( D => n4121, CK => CLK, SN => RST, Q =>
                           n3481, QN => n3649);
   clk_r_REG4640_S17 : DFFR_X1 port map( D => n3649, CK => CLK, RN => RST, Q =>
                           n_3923, QN => n3480);
   clk_r_REG4645_S16 : DFFS_X1 port map( D => n4122, CK => CLK, SN => RST, Q =>
                           n3479, QN => n3650);
   clk_r_REG4646_S17 : DFFR_X1 port map( D => n3650, CK => CLK, RN => RST, Q =>
                           n_3924, QN => n3478);
   clk_r_REG4651_S16 : DFFS_X1 port map( D => n4123, CK => CLK, SN => RST, Q =>
                           n3477, QN => n3651);
   clk_r_REG4652_S17 : DFFR_X1 port map( D => n3651, CK => CLK, RN => RST, Q =>
                           n_3925, QN => n3476);
   clk_r_REG4659_S16 : DFFS_X1 port map( D => n4124, CK => CLK, SN => RST, Q =>
                           n3475, QN => n3652);
   clk_r_REG4660_S17 : DFFR_X1 port map( D => n3652, CK => CLK, RN => RST, Q =>
                           n_3926, QN => n3474);
   clk_r_REG6783_S1 : DFFS_X1 port map( D => n4048, CK => CLK, SN => RST, Q => 
                           n3473, QN => n_3927);
   clk_r_REG4667_S16 : DFFS_X1 port map( D => n4125, CK => CLK, SN => RST, Q =>
                           n3472, QN => n3653);
   clk_r_REG4668_S17 : DFFR_X1 port map( D => n3653, CK => CLK, RN => RST, Q =>
                           n_3928, QN => n3471);
   clk_r_REG4678_S16 : DFFS_X1 port map( D => n4126, CK => CLK, SN => RST, Q =>
                           n3470, QN => n3632);
   clk_r_REG4679_S17 : DFFR_X1 port map( D => n3632, CK => CLK, RN => RST, Q =>
                           n_3929, QN => n3469);
   clk_r_REG4684_S16 : DFFS_X1 port map( D => n4127, CK => CLK, SN => RST, Q =>
                           n3468, QN => n3633);
   clk_r_REG4685_S17 : DFFR_X1 port map( D => n3633, CK => CLK, RN => RST, Q =>
                           n_3930, QN => n3467);
   clk_r_REG4696_S16 : DFFS_X1 port map( D => n4128, CK => CLK, SN => RST, Q =>
                           n3466, QN => n3634);
   clk_r_REG4697_S17 : DFFR_X1 port map( D => n3634, CK => CLK, RN => RST, Q =>
                           n_3931, QN => n3465);
   clk_r_REG4244_S6 : DFFS_X1 port map( D => n4118, CK => CLK, SN => RST, Q => 
                           n3464, QN => n3636);
   clk_r_REG4245_S7 : DFFR_X1 port map( D => n3636, CK => CLK, RN => RST, Q => 
                           n_3932, QN => n3463);
   clk_r_REG4572_S6 : DFFS_X1 port map( D => n3674, CK => CLK, SN => RST, Q => 
                           n3462, QN => n3637);
   clk_r_REG4573_S7 : DFFR_X1 port map( D => n3637, CK => CLK, RN => RST, Q => 
                           n_3933, QN => n3461);
   clk_r_REG4235_S6 : DFFS_X1 port map( D => n4130, CK => CLK, SN => RST, Q => 
                           n3460, QN => n3640);
   clk_r_REG4236_S7 : DFFR_X1 port map( D => n3640, CK => CLK, RN => RST, Q => 
                           n_3934, QN => n3459);
   clk_r_REG6907_S1 : DFFR_X1 port map( D => n4054, CK => CLK, RN => RST, Q => 
                           n3458, QN => n_3935);
   clk_r_REG3645_S4 : DFFR_X1 port map( D => n3654, CK => CLK, RN => RST, Q => 
                           n3457, QN => n_3936);
   clk_r_REG6876_S5 : DFFS_X1 port map( D => n4047, CK => CLK, SN => RST, Q => 
                           n3456, QN => n_3937);
   clk_r_REG4574_S7 : DFFR_X1 port map( D => n3637, CK => CLK, RN => RST, Q => 
                           n3455, QN => n_3938);
   clk_r_REG4237_S7 : DFFR_X1 port map( D => n3640, CK => CLK, RN => RST, Q => 
                           n3454, QN => n_3939);
   clk_r_REG4246_S7 : DFFR_X1 port map( D => n3636, CK => CLK, RN => RST, Q => 
                           n3453, QN => n_3940);
   clk_r_REG4698_S17 : DFFR_X1 port map( D => n3634, CK => CLK, RN => RST, Q =>
                           n3452, QN => n_3941);
   clk_r_REG4686_S17 : DFFR_X1 port map( D => n3633, CK => CLK, RN => RST, Q =>
                           n3451, QN => n_3942);
   clk_r_REG4680_S17 : DFFR_X1 port map( D => n3632, CK => CLK, RN => RST, Q =>
                           n3450, QN => n_3943);
   clk_r_REG4669_S17 : DFFR_X1 port map( D => n3653, CK => CLK, RN => RST, Q =>
                           n3449, QN => n_3944);
   clk_r_REG4653_S17 : DFFR_X1 port map( D => n3651, CK => CLK, RN => RST, Q =>
                           n3448, QN => n_3945);
   clk_r_REG4647_S17 : DFFR_X1 port map( D => n3650, CK => CLK, RN => RST, Q =>
                           n3447, QN => n_3946);
   clk_r_REG4641_S17 : DFFR_X1 port map( D => n3649, CK => CLK, RN => RST, Q =>
                           n3446, QN => n_3947);
   clk_r_REG4634_S17 : DFFR_X1 port map( D => n3648, CK => CLK, RN => RST, Q =>
                           n3445, QN => n_3948);
   clk_r_REG4626_S17 : DFFR_X1 port map( D => n3647, CK => CLK, RN => RST, Q =>
                           n3444, QN => n_3949);
   clk_r_REG5917_S4 : DFFR_X1 port map( D => n3654, CK => CLK, RN => RST, Q => 
                           n3443, QN => n_3950);
   clk_r_REG6708_S3 : DFFR_X1 port map( D => n4044, CK => CLK, RN => RST, Q => 
                           DRAM_ENABLE, QN => n_3951);
   clk_r_REG6195_S3 : DFFR_X1 port map( D => n3441, CK => CLK, RN => RST, Q => 
                           n3440, QN => n_3952);
   clk_r_REG6258_S2 : DFF_X1 port map( D => n1671, CK => CLK, Q => n3439, QN =>
                           n_3953);
   clk_r_REG6259_S3 : DFFR_X1 port map( D => n3439, CK => CLK, RN => RST, Q => 
                           n3438, QN => n_3954);
   clk_r_REG3639_S2 : DFF_X1 port map( D => n1669, CK => CLK, Q => n3437, QN =>
                           n_3955);
   clk_r_REG5934_S3 : DFFR_X1 port map( D => n3437, CK => CLK, RN => RST, Q => 
                           n3436, QN => n_3956);
   clk_r_REG3685_S2 : DFF_X1 port map( D => n1667, CK => CLK, Q => n3435, QN =>
                           n_3957);
   clk_r_REG3686_S3 : DFFR_X1 port map( D => n3435, CK => CLK, RN => RST, Q => 
                           n3434, QN => n_3958);
   clk_r_REG6323_S2 : DFF_X1 port map( D => n1665, CK => CLK, Q => n3433, QN =>
                           n_3959);
   clk_r_REG6324_S3 : DFFR_X1 port map( D => n3433, CK => CLK, RN => RST, Q => 
                           n3432, QN => n_3960);
   clk_r_REG6387_S2 : DFF_X1 port map( D => n1663, CK => CLK, Q => n3431, QN =>
                           n_3961);
   clk_r_REG6388_S3 : DFFR_X1 port map( D => n3431, CK => CLK, RN => RST, Q => 
                           n3430, QN => n_3962);
   clk_r_REG3776_S2 : DFF_X1 port map( D => n1661, CK => CLK, Q => n3429, QN =>
                           n_3963);
   clk_r_REG3777_S3 : DFFR_X1 port map( D => n3429, CK => CLK, RN => RST, Q => 
                           n3428, QN => n_3964);
   clk_r_REG6452_S2 : DFF_X1 port map( D => n1659, CK => CLK, Q => n3427, QN =>
                           n_3965);
   clk_r_REG6453_S3 : DFFR_X1 port map( D => n3427, CK => CLK, RN => RST, Q => 
                           n3426, QN => n_3966);
   clk_r_REG3707_S2 : DFF_X1 port map( D => n1657, CK => CLK, Q => n3425, QN =>
                           n_3967);
   clk_r_REG3708_S3 : DFFR_X1 port map( D => n3425, CK => CLK, RN => RST, Q => 
                           n3424, QN => n_3968);
   clk_r_REG5721_S2 : DFF_X1 port map( D => n1655, CK => CLK, Q => n3423, QN =>
                           n_3969);
   clk_r_REG5722_S3 : DFFR_X1 port map( D => n3423, CK => CLK, RN => RST, Q => 
                           n3422, QN => n_3970);
   clk_r_REG3760_S2 : DFF_X1 port map( D => n1653, CK => CLK, Q => n3421, QN =>
                           n_3971);
   clk_r_REG3761_S3 : DFFR_X1 port map( D => n3421, CK => CLK, RN => RST, Q => 
                           n3420, QN => n_3972);
   clk_r_REG5383_S2 : DFF_X1 port map( D => n1651, CK => CLK, Q => n3419, QN =>
                           n_3973);
   clk_r_REG5384_S3 : DFFR_X1 port map( D => n3419, CK => CLK, RN => RST, Q => 
                           n3418, QN => n_3974);
   clk_r_REG5447_S2 : DFF_X1 port map( D => n1649, CK => CLK, Q => n3417, QN =>
                           n_3975);
   clk_r_REG5448_S3 : DFFR_X1 port map( D => n3417, CK => CLK, RN => RST, Q => 
                           n3416, QN => n_3976);
   clk_r_REG5512_S2 : DFF_X1 port map( D => n1647, CK => CLK, Q => n3415, QN =>
                           n_3977);
   clk_r_REG5513_S3 : DFFR_X1 port map( D => n3415, CK => CLK, RN => RST, Q => 
                           n3414, QN => n_3978);
   clk_r_REG6002_S2 : DFF_X1 port map( D => n1645, CK => CLK, Q => n3413, QN =>
                           n_3979);
   clk_r_REG6003_S3 : DFFR_X1 port map( D => n3413, CK => CLK, RN => RST, Q => 
                           n3412, QN => n_3980);
   clk_r_REG6067_S2 : DFF_X1 port map( D => n1643, CK => CLK, Q => n3411, QN =>
                           n_3981);
   clk_r_REG6068_S3 : DFFR_X1 port map( D => n3411, CK => CLK, RN => RST, Q => 
                           n3410, QN => n_3982);
   clk_r_REG5130_S2 : DFF_X1 port map( D => n1641, CK => CLK, Q => n3409, QN =>
                           n_3983);
   clk_r_REG5131_S3 : DFFR_X1 port map( D => n3409, CK => CLK, RN => RST, Q => 
                           n3408, QN => n_3984);
   clk_r_REG3889_S2 : DFF_X1 port map( D => n1639, CK => CLK, Q => n3407, QN =>
                           n_3985);
   clk_r_REG3890_S3 : DFFR_X1 port map( D => n3407, CK => CLK, RN => RST, Q => 
                           n3406, QN => n_3986);
   clk_r_REG3960_S2 : DFF_X1 port map( D => n1637, CK => CLK, Q => n3405, QN =>
                           n_3987);
   clk_r_REG3961_S3 : DFFR_X1 port map( D => n3405, CK => CLK, RN => RST, Q => 
                           n3404, QN => n_3988);
   clk_r_REG5194_S2 : DFF_X1 port map( D => n1635, CK => CLK, Q => n3403, QN =>
                           n_3989);
   clk_r_REG5195_S3 : DFFR_X1 port map( D => n3403, CK => CLK, RN => RST, Q => 
                           n3402, QN => n_3990);
   clk_r_REG5065_S2 : DFF_X1 port map( D => n1633, CK => CLK, Q => n3401, QN =>
                           n_3991);
   clk_r_REG5066_S3 : DFFR_X1 port map( D => n3401, CK => CLK, RN => RST, Q => 
                           n3400, QN => n_3992);
   clk_r_REG5847_S2 : DFF_X1 port map( D => n1631, CK => CLK, Q => n3399, QN =>
                           n_3993);
   clk_r_REG5848_S3 : DFFR_X1 port map( D => n3399, CK => CLK, RN => RST, Q => 
                           n3398, QN => n_3994);
   clk_r_REG4093_S2 : DFF_X1 port map( D => n1629, CK => CLK, Q => n3397, QN =>
                           n_3995);
   clk_r_REG4094_S3 : DFFR_X1 port map( D => n3397, CK => CLK, RN => RST, Q => 
                           n3396, QN => n_3996);
   clk_r_REG6516_S2 : DFF_X1 port map( D => n1627, CK => CLK, Q => n3395, QN =>
                           n_3997);
   clk_r_REG6517_S3 : DFFR_X1 port map( D => n3395, CK => CLK, RN => RST, Q => 
                           n3394, QN => n_3998);
   clk_r_REG4149_S2 : DFF_X1 port map( D => n1625, CK => CLK, Q => n3393, QN =>
                           n_3999);
   clk_r_REG4150_S3 : DFFR_X1 port map( D => n3393, CK => CLK, RN => RST, Q => 
                           n3392, QN => n_4000);
   clk_r_REG6580_S2 : DFF_X1 port map( D => n1623, CK => CLK, Q => n3391, QN =>
                           n_4001);
   clk_r_REG6581_S3 : DFFR_X1 port map( D => n3391, CK => CLK, RN => RST, Q => 
                           n3390, QN => n_4002);
   clk_r_REG4706_S2 : DFF_X1 port map( D => n1621, CK => CLK, Q => n3389, QN =>
                           n_4003);
   clk_r_REG4707_S3 : DFFR_X1 port map( D => n3389, CK => CLK, RN => RST, Q => 
                           n3388, QN => n_4004);
   clk_r_REG4489_S2 : DFF_X1 port map( D => n1619, CK => CLK, Q => n3387, QN =>
                           n_4005);
   clk_r_REG4781_S2 : DFF_X1 port map( D => n1617, CK => CLK, Q => n3386, QN =>
                           n_4006);
   clk_r_REG4927_S2 : DFF_X1 port map( D => n1615, CK => CLK, Q => n3385, QN =>
                           n_4007);
   clk_r_REG5583_S2 : DFF_X1 port map( D => n1614, CK => CLK, Q => n3384, QN =>
                           n_4008);
   clk_r_REG6131_S2 : DFF_X1 port map( D => n1613, CK => CLK, Q => n3383, QN =>
                           n_4009);
   clk_r_REG3581_S2 : DFF_X1 port map( D => n1611, CK => CLK, Q => n3382, QN =>
                           n_4010);
   clk_r_REG3582_S3 : DFFR_X1 port map( D => n3382, CK => CLK, RN => RST, Q => 
                           n3381, QN => n_4011);
   clk_r_REG3583_S4 : DFFR_X1 port map( D => n3381, CK => CLK, RN => RST, Q => 
                           n3380, QN => n_4012);
   clk_r_REG3573_S2 : DFF_X1 port map( D => n1608, CK => CLK, Q => n3379, QN =>
                           n_4013);
   clk_r_REG3574_S3 : DFFR_X1 port map( D => n3379, CK => CLK, RN => RST, Q => 
                           n3378, QN => n_4014);
   clk_r_REG3575_S4 : DFFR_X1 port map( D => n3378, CK => CLK, RN => RST, Q => 
                           n3377, QN => n_4015);
   clk_r_REG3629_S2 : DFF_X1 port map( D => n1605, CK => CLK, Q => n3376, QN =>
                           n_4016);
   clk_r_REG3630_S3 : DFFR_X1 port map( D => n3376, CK => CLK, RN => RST, Q => 
                           n3375, QN => n_4017);
   clk_r_REG3631_S4 : DFFR_X1 port map( D => n3375, CK => CLK, RN => RST, Q => 
                           n3374, QN => n_4018);
   clk_r_REG3677_S2 : DFF_X1 port map( D => n1602, CK => CLK, Q => n3373, QN =>
                           n_4019);
   clk_r_REG3678_S3 : DFFR_X1 port map( D => n3373, CK => CLK, RN => RST, Q => 
                           n3372, QN => n_4020);
   clk_r_REG3679_S4 : DFFR_X1 port map( D => n3372, CK => CLK, RN => RST, Q => 
                           n3371, QN => n_4021);
   clk_r_REG3563_S2 : DFF_X1 port map( D => n1599, CK => CLK, Q => n3370, QN =>
                           n_4022);
   clk_r_REG3564_S3 : DFFR_X1 port map( D => n3370, CK => CLK, RN => RST, Q => 
                           n3369, QN => n_4023);
   clk_r_REG3565_S4 : DFFR_X1 port map( D => n3369, CK => CLK, RN => RST, Q => 
                           n3368, QN => n_4024);
   clk_r_REG3554_S2 : DFF_X1 port map( D => n1596, CK => CLK, Q => n3367, QN =>
                           n_4025);
   clk_r_REG3555_S3 : DFFR_X1 port map( D => n3367, CK => CLK, RN => RST, Q => 
                           n3366, QN => n_4026);
   clk_r_REG3556_S4 : DFFR_X1 port map( D => n3366, CK => CLK, RN => RST, Q => 
                           n3365, QN => n_4027);
   clk_r_REG3769_S2 : DFF_X1 port map( D => n1593, CK => CLK, Q => n3364, QN =>
                           n_4028);
   clk_r_REG3770_S3 : DFFR_X1 port map( D => n3364, CK => CLK, RN => RST, Q => 
                           n3363, QN => n_4029);
   clk_r_REG3771_S4 : DFFR_X1 port map( D => n3363, CK => CLK, RN => RST, Q => 
                           n3362, QN => n_4030);
   clk_r_REG3546_S2 : DFF_X1 port map( D => n1590, CK => CLK, Q => n3361, QN =>
                           n_4031);
   clk_r_REG3547_S3 : DFFR_X1 port map( D => n3361, CK => CLK, RN => RST, Q => 
                           n3360, QN => n_4032);
   clk_r_REG3548_S4 : DFFR_X1 port map( D => n3360, CK => CLK, RN => RST, Q => 
                           n3359, QN => n_4033);
   clk_r_REG3702_S2 : DFF_X1 port map( D => n1587, CK => CLK, Q => n3358, QN =>
                           n_4034);
   clk_r_REG3703_S3 : DFFR_X1 port map( D => n3358, CK => CLK, RN => RST, Q => 
                           n3357, QN => n_4035);
   clk_r_REG3704_S4 : DFFR_X1 port map( D => n3357, CK => CLK, RN => RST, Q => 
                           n3356, QN => n_4036);
   clk_r_REG3695_S2 : DFF_X1 port map( D => n1584, CK => CLK, Q => n3355, QN =>
                           n_4037);
   clk_r_REG3696_S3 : DFFR_X1 port map( D => n3355, CK => CLK, RN => RST, Q => 
                           n3354, QN => n_4038);
   clk_r_REG3697_S4 : DFFR_X1 port map( D => n3354, CK => CLK, RN => RST, Q => 
                           n3353, QN => n_4039);
   clk_r_REG3754_S2 : DFF_X1 port map( D => n1581, CK => CLK, Q => n3352, QN =>
                           n_4040);
   clk_r_REG3755_S3 : DFFR_X1 port map( D => n3352, CK => CLK, RN => RST, Q => 
                           n3351, QN => n_4041);
   clk_r_REG3756_S4 : DFFR_X1 port map( D => n3351, CK => CLK, RN => RST, Q => 
                           n3350, QN => n_4042);
   clk_r_REG3747_S2 : DFF_X1 port map( D => n1578, CK => CLK, Q => n3349, QN =>
                           n_4043);
   clk_r_REG3748_S3 : DFFR_X1 port map( D => n3349, CK => CLK, RN => RST, Q => 
                           n3348, QN => n_4044);
   clk_r_REG3749_S4 : DFFR_X1 port map( D => n3348, CK => CLK, RN => RST, Q => 
                           n3347, QN => n_4045);
   clk_r_REG3740_S2 : DFF_X1 port map( D => n1575, CK => CLK, Q => n3346, QN =>
                           n_4046);
   clk_r_REG3741_S3 : DFFR_X1 port map( D => n3346, CK => CLK, RN => RST, Q => 
                           n3345, QN => n_4047);
   clk_r_REG3742_S4 : DFFR_X1 port map( D => n3345, CK => CLK, RN => RST, Q => 
                           n3344, QN => n_4048);
   clk_r_REG3733_S2 : DFF_X1 port map( D => n1572, CK => CLK, Q => n3343, QN =>
                           n_4049);
   clk_r_REG3734_S3 : DFFR_X1 port map( D => n3343, CK => CLK, RN => RST, Q => 
                           n3342, QN => n_4050);
   clk_r_REG3735_S4 : DFFR_X1 port map( D => n3342, CK => CLK, RN => RST, Q => 
                           n3341, QN => n_4051);
   clk_r_REG3617_S2 : DFF_X1 port map( D => n1569, CK => CLK, Q => n3340, QN =>
                           n_4052);
   clk_r_REG3618_S3 : DFFR_X1 port map( D => n3340, CK => CLK, RN => RST, Q => 
                           n3339, QN => n_4053);
   clk_r_REG3619_S4 : DFFR_X1 port map( D => n3339, CK => CLK, RN => RST, Q => 
                           n3338, QN => n_4054);
   clk_r_REG3610_S2 : DFF_X1 port map( D => n1566, CK => CLK, Q => n3337, QN =>
                           n_4055);
   clk_r_REG3611_S3 : DFFR_X1 port map( D => n3337, CK => CLK, RN => RST, Q => 
                           n3336, QN => n_4056);
   clk_r_REG3612_S4 : DFFR_X1 port map( D => n3336, CK => CLK, RN => RST, Q => 
                           n3335, QN => n_4057);
   clk_r_REG3831_S2 : DFF_X1 port map( D => n1563, CK => CLK, Q => n3334, QN =>
                           n_4058);
   clk_r_REG3832_S3 : DFFR_X1 port map( D => n3334, CK => CLK, RN => RST, Q => 
                           n3333, QN => n_4059);
   clk_r_REG3833_S4 : DFFR_X1 port map( D => n3333, CK => CLK, RN => RST, Q => 
                           n3332, QN => n_4060);
   clk_r_REG3881_S2 : DFF_X1 port map( D => n1560, CK => CLK, Q => n3331, QN =>
                           n_4061);
   clk_r_REG3882_S3 : DFFR_X1 port map( D => n3331, CK => CLK, RN => RST, Q => 
                           n3330, QN => n_4062);
   clk_r_REG3883_S4 : DFFR_X1 port map( D => n3330, CK => CLK, RN => RST, Q => 
                           n3329, QN => n_4063);
   clk_r_REG3950_S2 : DFF_X1 port map( D => n1557, CK => CLK, Q => n3328, QN =>
                           n_4064);
   clk_r_REG3951_S3 : DFFR_X1 port map( D => n3328, CK => CLK, RN => RST, Q => 
                           n3327, QN => n_4065);
   clk_r_REG3952_S4 : DFFR_X1 port map( D => n3327, CK => CLK, RN => RST, Q => 
                           n3326, QN => n_4066);
   clk_r_REG3785_S2 : DFF_X1 port map( D => n1554, CK => CLK, Q => n3325, QN =>
                           n_4067);
   clk_r_REG3786_S3 : DFFR_X1 port map( D => n3325, CK => CLK, RN => RST, Q => 
                           n3324, QN => n_4068);
   clk_r_REG3787_S4 : DFFR_X1 port map( D => n3324, CK => CLK, RN => RST, Q => 
                           n3323, QN => n_4069);
   clk_r_REG3856_S2 : DFF_X1 port map( D => n1551, CK => CLK, Q => n3322, QN =>
                           n_4070);
   clk_r_REG3857_S3 : DFFR_X1 port map( D => n3322, CK => CLK, RN => RST, Q => 
                           n3321, QN => n_4071);
   clk_r_REG3858_S4 : DFFR_X1 port map( D => n3321, CK => CLK, RN => RST, Q => 
                           n3320, QN => n_4072);
   clk_r_REG3659_S2 : DFF_X1 port map( D => n1548, CK => CLK, Q => n3319, QN =>
                           n_4073);
   clk_r_REG3660_S3 : DFFR_X1 port map( D => n3319, CK => CLK, RN => RST, Q => 
                           n3318, QN => n_4074);
   clk_r_REG3661_S4 : DFFR_X1 port map( D => n3318, CK => CLK, RN => RST, Q => 
                           n3317, QN => n_4075);
   clk_r_REG4062_S2 : DFF_X1 port map( D => n1545, CK => CLK, Q => n3316, QN =>
                           n_4076);
   clk_r_REG4063_S3 : DFFR_X1 port map( D => n3316, CK => CLK, RN => RST, Q => 
                           n3315, QN => n_4077);
   clk_r_REG4064_S4 : DFFR_X1 port map( D => n3315, CK => CLK, RN => RST, Q => 
                           n3314, QN => n_4078);
   clk_r_REG3532_S2 : DFF_X1 port map( D => n1542, CK => CLK, Q => n3313, QN =>
                           n_4079);
   clk_r_REG3533_S3 : DFFR_X1 port map( D => n3313, CK => CLK, RN => RST, Q => 
                           n3312, QN => n_4080);
   clk_r_REG3534_S4 : DFFR_X1 port map( D => n3312, CK => CLK, RN => RST, Q => 
                           n3311, QN => n_4081);
   clk_r_REG4129_S2 : DFF_X1 port map( D => n1539, CK => CLK, Q => n3310, QN =>
                           n_4082);
   clk_r_REG4130_S3 : DFFR_X1 port map( D => n3310, CK => CLK, RN => RST, Q => 
                           n3309, QN => n_4083);
   clk_r_REG4131_S4 : DFFR_X1 port map( D => n3309, CK => CLK, RN => RST, Q => 
                           n3308, QN => n_4084);
   clk_r_REG3519_S2 : DFF_X1 port map( D => n1536, CK => CLK, Q => n3307, QN =>
                           n_4085);
   clk_r_REG3520_S3 : DFFR_X1 port map( D => n3307, CK => CLK, RN => RST, Q => 
                           n3306, QN => n_4086);
   clk_r_REG3521_S4 : DFFR_X1 port map( D => n3306, CK => CLK, RN => RST, Q => 
                           n3305, QN => n_4087);
   clk_r_REG3994_S2 : DFF_X1 port map( D => n1533, CK => CLK, Q => n3304, QN =>
                           n_4088);
   clk_r_REG3995_S3 : DFFR_X1 port map( D => n3304, CK => CLK, RN => RST, Q => 
                           n3303, QN => n_4089);
   clk_r_REG3996_S4 : DFFR_X1 port map( D => n3303, CK => CLK, RN => RST, Q => 
                           n3302, QN => n_4090);
   clk_r_REG4049_S2 : DFF_X1 port map( D => n1530, CK => CLK, Q => n3301, QN =>
                           n_4091);
   clk_r_REG4050_S3 : DFFR_X1 port map( D => n3301, CK => CLK, RN => RST, Q => 
                           n3300, QN => n_4092);
   clk_r_REG4051_S4 : DFFR_X1 port map( D => n3300, CK => CLK, RN => RST, Q => 
                           n3299, QN => n_4093);
   clk_r_REG3980_S2 : DFF_X1 port map( D => n1527, CK => CLK, Q => n3298, QN =>
                           n_4094);
   clk_r_REG3981_S3 : DFFR_X1 port map( D => n3298, CK => CLK, RN => RST, Q => 
                           n3297, QN => n_4095);
   clk_r_REG3982_S4 : DFFR_X1 port map( D => n3297, CK => CLK, RN => RST, Q => 
                           n3296, QN => n_4096);
   clk_r_REG3937_S2 : DFF_X1 port map( D => n1524, CK => CLK, Q => n3295, QN =>
                           n_4097);
   clk_r_REG3938_S3 : DFFR_X1 port map( D => n3295, CK => CLK, RN => RST, Q => 
                           n3294, QN => n_4098);
   clk_r_REG3939_S4 : DFFR_X1 port map( D => n3294, CK => CLK, RN => RST, Q => 
                           n3293, QN => n_4099);
   clk_r_REG3716_S2 : DFF_X1 port map( D => n1521, CK => CLK, Q => n3292, QN =>
                           n_4100);
   clk_r_REG3717_S3 : DFFR_X1 port map( D => n3292, CK => CLK, RN => RST, Q => 
                           n3291, QN => n_4101);
   clk_r_REG3718_S4 : DFFR_X1 port map( D => n3291, CK => CLK, RN => RST, Q => 
                           n3290, QN => n_4102);
   clk_r_REG3590_S2 : DFF_X1 port map( D => n1518, CK => CLK, Q => n3289, QN =>
                           n_4103);
   clk_r_REG3591_S3 : DFFR_X1 port map( D => n3289, CK => CLK, RN => RST, Q => 
                           n3288, QN => n_4104);
   clk_r_REG3592_S4 : DFFR_X1 port map( D => n3288, CK => CLK, RN => RST, Q => 
                           n3287, QN => n_4105);
   clk_r_REG6821_S8 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port, CK =>
                           CLK, RN => RST, Q => n3286, QN => n_4106);
   clk_r_REG6824_S8 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port, CK =>
                           CLK, RN => RST, Q => n3285, QN => n_4107);
   clk_r_REG6904_S3 : DFFR_X1 port map( D => n1513, CK => CLK, RN => RST, Q => 
                           n3284, QN => n4429);
   clk_r_REG6905_S5 : DFFR_X1 port map( D => n1512, CK => CLK, RN => RST, Q => 
                           n4417, QN => n3670);
   clk_r_REG6784_S3 : DFFS_X1 port map( D => n4039, CK => CLK, SN => RST, Q => 
                           n_4108, QN => n3282);
   clk_r_REG6906_S3 : DFFR_X1 port map( D => n1510, CK => CLK, RN => RST, Q => 
                           n3281, QN => n4418);
   clk_r_REG6823_S8 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port, CK =>
                           CLK, RN => RST, Q => n3280, QN => n_4109);
   clk_r_REG6646_S3 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port, CK =>
                           CLK, RN => RST, Q => n3279, QN => n_4110);
   clk_r_REG6658_S2 : DFFR_X1 port map( D => n3635, CK => CLK, RN => RST, Q => 
                           n4421, QN => n3277);
   clk_r_REG6710_S3 : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => CLK, 
                           RN => RST, Q => n3276, QN => n_4111);
   clk_r_REG6864_S6 : DFFR_X1 port map( D => n4055, CK => CLK, RN => RST, Q => 
                           n_4112, QN => n3275);
   clk_r_REG6863_S6 : DFFS_X1 port map( D => n474, CK => CLK, SN => RST, Q => 
                           n_4113, QN => n3639);
   clk_r_REG6857_S3 : DFFS_X1 port map( D => n4059, CK => CLK, SN => RST, Q => 
                           n_4114, QN => n3273);
   clk_r_REG6775_S3 : DFFR_X1 port map( D => cu_i_n135, CK => CLK, RN => RST, Q
                           => n3272, QN => n_4115);
   clk_r_REG6855_S6 : DFFR_X1 port map( D => n1500, CK => CLK, RN => RST, Q => 
                           n3271, QN => n_4116);
   clk_r_REG6859_S6 : DFFS_X1 port map( D => n2299, CK => CLK, SN => RST, Q => 
                           n_4117, QN => n3638);
   clk_r_REG6663_S3 : DFFR_X1 port map( D => n1498, CK => CLK, RN => RST, Q => 
                           n3269, QN => n_4118);
   clk_r_REG6785_S3 : DFFS_X1 port map( D => n4038, CK => CLK, SN => RST, Q => 
                           n_4119, QN => n3268);
   clk_r_REG6782_S1 : DFFS_X1 port map( D => n4048, CK => CLK, SN => RST, Q => 
                           n3643, QN => n_4120);
   clk_r_REG6715_S5 : DFFS_X1 port map( D => n3658, CK => CLK, SN => RST, Q => 
                           n_4121, QN => n3266);
   clk_r_REG4233_S5 : DFFR_X1 port map( D => n2359, CK => CLK, RN => RST, Q => 
                           n3265, QN => n_4122);
   clk_r_REG4238_S5 : DFFS_X1 port map( D => n2358, CK => CLK, SN => RST, Q => 
                           n3264, QN => n_4123);
   clk_r_REG4239_S5 : DFFR_X1 port map( D => n2363, CK => CLK, RN => RST, Q => 
                           n3263, QN => n_4124);
   clk_r_REG4571_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_5_port, CK => CLK, RN
                           => RST, Q => n3262, QN => n3674);
   clk_r_REG4568_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_4_port, CK => CLK, RN
                           => RST, Q => n3260, QN => n3644);
   clk_r_REG3646_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_6_port, CK => CLK, RN
                           => RST, Q => n3259, QN => n3675);
   clk_r_REG5927_S3 : DFFS_X1 port map( D => n1758, CK => CLK, SN => RST, Q => 
                           n3258, QN => n_4125);
   clk_r_REG3643_S3 : DFFS_X1 port map( D => n1505, CK => CLK, SN => RST, Q => 
                           n_4126, QN => n3654);
   clk_r_REG6644_S1 : DFFS_X1 port map( D => n477, CK => CLK, SN => RST, Q => 
                           n3253, QN => n_4127);
   clk_r_REG6908_S2 : DFFS_X1 port map( D => n2416, CK => CLK, SN => RST, Q => 
                           n3252, QN => n_4128);
   clk_r_REG4004_S8 : DFFS_X1 port map( D => n2483, CK => CLK, SN => RST, Q => 
                           n3251, QN => n_4129);
   clk_r_REG4006_S8 : DFFR_X1 port map( D => n2486, CK => CLK, RN => RST, Q => 
                           n3250, QN => n_4130);
   clk_r_REG4007_S8 : DFFS_X1 port map( D => n2485, CK => CLK, SN => RST, Q => 
                           n3249, QN => n_4131);
   clk_r_REG6826_S6 : DFFR_X1 port map( D => n1477, CK => CLK, RN => RST, Q => 
                           n3248, QN => n_4132);
   clk_r_REG6820_S6 : DFFS_X1 port map( D => n492, CK => CLK, SN => RST, Q => 
                           n3247, QN => n_4133);
   clk_r_REG6656_S1 : DFFR_X1 port map( D => n1475, CK => CLK, RN => RST, Q => 
                           n3246, QN => n4423);
   clk_r_REG6657_S2 : DFFR_X1 port map( D => n3246, CK => CLK, RN => RST, Q => 
                           n3245, QN => n_4134);
   clk_r_REG4852_S5 : DFFR_X1 port map( D => n1328, CK => CLK, RN => RST, Q => 
                           n3244, QN => n3673);
   clk_r_REG4618_S7 : DFFS_X1 port map( D => n1460, CK => CLK, SN => RST, Q => 
                           n3243, QN => n_4135);
   clk_r_REG3640_S2 : DFF_X1 port map( D => n2530, CK => CLK, Q => n3242, QN =>
                           n_4136);
   clk_r_REG6774_S3 : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK => CLK, 
                           RN => RST, Q => n3240, QN => n_4137);
   clk_r_REG6858_S6 : DFFS_X1 port map( D => n464, CK => CLK, SN => RST, Q => 
                           n3239, QN => n_4138);
   clk_r_REG6819_S6 : DFFR_X1 port map( D => n1394, CK => CLK, RN => RST, Q => 
                           n3238, QN => n_4139);
   clk_r_REG6825_S6 : DFFR_X1 port map( D => n1390, CK => CLK, RN => RST, Q => 
                           n3237, QN => n3664);
   clk_r_REG6827_S6 : DFFR_X1 port map( D => n1393, CK => CLK, RN => RST, Q => 
                           n3236, QN => n_4140);
   clk_r_REG6786_S3 : DFFS_X1 port map( D => n1458, CK => CLK, SN => RST, Q => 
                           n3235, QN => n_4141);
   clk_r_REG6877_S6 : DFFR_X1 port map( D => curr_instruction_to_cu_i_19_port, 
                           CK => CLK, RN => RST, Q => n3234, QN => n_4142);
   clk_r_REG6880_S6 : DFFR_X1 port map( D => n1404, CK => CLK, RN => RST, Q => 
                           n3233, QN => n_4143);
   clk_r_REG6881_S6 : DFFR_X1 port map( D => curr_instruction_to_cu_i_17_port, 
                           CK => CLK, RN => RST, Q => n3232, QN => n_4144);
   clk_r_REG6882_S6 : DFFR_X1 port map( D => n1402, CK => CLK, RN => RST, Q => 
                           n3231, QN => n_4145);
   clk_r_REG6883_S6 : DFFR_X1 port map( D => curr_instruction_to_cu_i_20_port, 
                           CK => CLK, RN => RST, Q => n3230, QN => n_4146);
   clk_r_REG6886_S6 : DFFR_X1 port map( D => curr_instruction_to_cu_i_16_port, 
                           CK => CLK, RN => RST, Q => n3228, QN => n_4147);
   clk_r_REG6828_S6 : DFFR_X1 port map( D => n1401, CK => CLK, RN => RST, Q => 
                           n3227, QN => n_4148);
   clk_r_REG6645_S1 : DFFS_X1 port map( D => n3629, CK => CLK, SN => RST, Q => 
                           IRAM_ENABLE, QN => n_4149);
   clk_r_REG4247_S12 : DFFS_X1 port map( D => n4110, CK => CLK, SN => RST, Q =>
                           n_4150, QN => n3225);
   clk_r_REG4009_S15 : DFFS_X1 port map( D => n4108, CK => CLK, SN => RST, Q =>
                           n_4151, QN => n3224);
   clk_r_REG4014_S5 : DFFS_X1 port map( D => n4101, CK => CLK, SN => RST, Q => 
                           n_4152, QN => n3223);
   clk_r_REG4020_S5 : DFFS_X1 port map( D => n4095, CK => CLK, SN => RST, Q => 
                           n_4153, QN => n3222);
   clk_r_REG4026_S12 : DFFS_X1 port map( D => n4094, CK => CLK, SN => RST, Q =>
                           n_4154, QN => n3221);
   clk_r_REG4032_S12 : DFFS_X1 port map( D => n4093, CK => CLK, SN => RST, Q =>
                           n_4155, QN => n3220);
   clk_r_REG4038_S6 : DFFS_X1 port map( D => n4092, CK => CLK, SN => RST, Q => 
                           n_4156, QN => n3219);
   clk_r_REG4582_S5 : DFFS_X1 port map( D => n4091, CK => CLK, SN => RST, Q => 
                           n_4157, QN => n3218);
   clk_r_REG4588_S12 : DFFS_X1 port map( D => n4090, CK => CLK, SN => RST, Q =>
                           n_4158, QN => n3217);
   clk_r_REG4594_S6 : DFFS_X1 port map( D => n4089, CK => CLK, SN => RST, Q => 
                           n_4159, QN => n3216);
   clk_r_REG4600_S12 : DFFS_X1 port map( D => n4088, CK => CLK, SN => RST, Q =>
                           n_4160, QN => n3215);
   clk_r_REG4616_S6 : DFFR_X1 port map( D => n1916, CK => CLK, RN => RST, Q => 
                           n3214, QN => n_4161);
   clk_r_REG4608_S6 : DFFS_X1 port map( D => n4087, CK => CLK, SN => RST, Q => 
                           n_4162, QN => n3213);
   clk_r_REG6778_S4 : DFFS_X1 port map( D => n4041, CK => CLK, SN => RST, Q => 
                           n_4163, QN => n3212);
   clk_r_REG6712_S4 : DFFR_X1 port map( D => n1425, CK => CLK, RN => RST, Q => 
                           n3211, QN => n_4164);
   clk_r_REG6709_S4 : DFFR_X1 port map( D => n1424, CK => CLK, RN => RST, Q => 
                           n3210, QN => n_4165);
   clk_r_REG6699_S4 : DFFR_X1 port map( D => n1423, CK => CLK, RN => RST, Q => 
                           n3209, QN => n_4166);
   clk_r_REG6664_S4 : DFFR_X1 port map( D => n1422, CK => CLK, RN => RST, Q => 
                           n3208, QN => n4424);
   clk_r_REG6829_S6 : DFFR_X1 port map( D => n1415, CK => CLK, RN => RST, Q => 
                           n3207, QN => n_4167);
   clk_r_REG6847_S6 : DFFR_X1 port map( D => n1414, CK => CLK, RN => RST, Q => 
                           n3206, QN => n_4168);
   clk_r_REG6887_S6 : DFFR_X1 port map( D => n1413, CK => CLK, RN => RST, Q => 
                           n3205, QN => n_4169);
   clk_r_REG6902_S6 : DFFR_X1 port map( D => n1412, CK => CLK, RN => RST, Q => 
                           n3204, QN => n_4170);
   clk_r_REG6903_S6 : DFFR_X1 port map( D => n1411, CK => CLK, RN => RST, Q => 
                           n3203, QN => n_4171);
   clk_r_REG6850_S6 : DFFR_X1 port map( D => n1400, CK => CLK, RN => RST, Q => 
                           n3202, QN => n_4172);
   clk_r_REG6851_S6 : DFFR_X1 port map( D => n1399, CK => CLK, RN => RST, Q => 
                           n3201, QN => n_4173);
   clk_r_REG6852_S6 : DFFR_X1 port map( D => n1398, CK => CLK, RN => RST, Q => 
                           n3200, QN => n_4174);
   clk_r_REG6853_S6 : DFFR_X1 port map( D => n1397, CK => CLK, RN => RST, Q => 
                           n3199, QN => n_4175);
   clk_r_REG6854_S6 : DFFR_X1 port map( D => n1396, CK => CLK, RN => RST, Q => 
                           n3198, QN => n_4176);
   clk_r_REG6739_S4 : DFFR_X1 port map( D => n1383, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3197, QN => n_4177);
   clk_r_REG6740_S4 : DFFR_X1 port map( D => n1382, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3196, QN => n_4178);
   clk_r_REG6741_S4 : DFFR_X1 port map( D => n1381, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3195, QN => n_4179);
   clk_r_REG6742_S4 : DFFR_X1 port map( D => n1380, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3194, QN => n_4180);
   clk_r_REG6743_S4 : DFFR_X1 port map( D => n1379, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3193, QN => n_4181);
   clk_r_REG6744_S4 : DFFR_X1 port map( D => n1378, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3192, QN => n_4182);
   clk_r_REG6745_S4 : DFFR_X1 port map( D => n1377, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3191, QN => n_4183);
   clk_r_REG6746_S4 : DFFR_X1 port map( D => n1376, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3190, QN => n_4184);
   clk_r_REG6747_S4 : DFFR_X1 port map( D => n1375, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3189, QN => n_4185);
   clk_r_REG6748_S4 : DFFR_X1 port map( D => n1374, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3188, QN => n_4186);
   clk_r_REG6749_S4 : DFFR_X1 port map( D => n1373, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3187, QN => n_4187);
   clk_r_REG6750_S4 : DFFR_X1 port map( D => n1372, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3186, QN => n_4188);
   clk_r_REG6751_S4 : DFFR_X1 port map( D => n1371, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3185, QN => n_4189);
   clk_r_REG6752_S4 : DFFR_X1 port map( D => n1370, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3184, QN => n_4190);
   clk_r_REG6753_S4 : DFFR_X1 port map( D => n1369, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3183, QN => n_4191);
   clk_r_REG6754_S4 : DFFR_X1 port map( D => n1368, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3182, QN => n_4192);
   clk_r_REG6755_S4 : DFFR_X1 port map( D => n1367, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3181, QN => n_4193);
   clk_r_REG6756_S4 : DFFR_X1 port map( D => n1366, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3180, QN => n_4194);
   clk_r_REG6757_S4 : DFFR_X1 port map( D => n1365, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3179, QN => n_4195);
   clk_r_REG6758_S4 : DFFR_X1 port map( D => n1364, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3178, QN => n_4196);
   clk_r_REG6759_S4 : DFFR_X1 port map( D => n1363, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3177, QN => n_4197);
   clk_r_REG6760_S4 : DFFR_X1 port map( D => n1362, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3176, QN => n_4198);
   clk_r_REG6761_S4 : DFFR_X1 port map( D => n1361, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3175, QN => n_4199);
   clk_r_REG6762_S4 : DFFR_X1 port map( D => n1360, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3174, QN => n_4200);
   clk_r_REG6763_S4 : DFFR_X1 port map( D => n1359, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3173, QN => n_4201);
   clk_r_REG6764_S4 : DFFR_X1 port map( D => n1358, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3172, QN => n_4202);
   clk_r_REG6765_S4 : DFFR_X1 port map( D => n1357, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3171, QN => n_4203);
   clk_r_REG6766_S4 : DFFR_X1 port map( D => n1356, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3170, QN => n_4204);
   clk_r_REG6767_S4 : DFFR_X1 port map( D => n1355, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3169, QN => n_4205);
   clk_r_REG6768_S4 : DFFR_X1 port map( D => n1354, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3168, QN => n_4206);
   clk_r_REG6769_S4 : DFFR_X1 port map( D => n1353, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3167, QN => n_4207);
   clk_r_REG6770_S4 : DFFR_X1 port map( D => n1352, CK => 
                           datapath_i_decode_stage_dp_clk_immediate, RN => RST,
                           Q => n3166, QN => n_4208);
   clk_r_REG5918_S5 : DFFR_X1 port map( D => n3628, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_0_port, QN => n_4209);
   clk_r_REG5919_S5 : DFFR_X1 port map( D => n1388, CK => CLK, RN => RST, Q => 
                           n3164, QN => n3676);
   clk_r_REG5654_S5 : DFFR_X1 port map( D => n3627, CK => CLK, RN => RST, Q => 
                           IRAM_ADDRESS_1_port, QN => n_4210);
   clk_r_REG5655_S5 : DFFR_X1 port map( D => n1385, CK => CLK, RN => RST, Q => 
                           n3162, QN => n3671);
   clk_r_REG5001_S5 : DFFR_X1 port map( D => n2547, CK => CLK, RN => RST, Q => 
                           n3161, QN => n_4211);
   clk_r_REG6700_S5 : DFFR_X1 port map( D => n1779, CK => CLK, RN => RST, Q => 
                           n3160, QN => n_4212);
   clk_r_REG6861_S6 : DFFR_X1 port map( D => n4064, CK => CLK, RN => RST, Q => 
                           n_4213, QN => n3159);
   clk_r_REG6867_S6 : DFFR_X1 port map( D => n4061, CK => CLK, RN => RST, Q => 
                           n4427, QN => n3158);
   clk_r_REG6704_S3 : DFFR_X1 port map( D => n4044, CK => CLK, RN => RST, Q => 
                           n_4214, QN => n4426);
   clk_r_REG6862_S1 : DFFR_X1 port map( D => n1350, CK => CLK, RN => RST, Q => 
                           n3155, QN => n_4215);
   clk_r_REG6856_S6 : DFFR_X1 port map( D => n4060, CK => CLK, RN => RST, Q => 
                           n_4216, QN => n3154);
   clk_r_REG6870_S6 : DFFR_X1 port map( D => n4051, CK => CLK, RN => RST, Q => 
                           n_4217, QN => n3153);
   clk_r_REG6872_S6 : DFFR_X1 port map( D => n4050, CK => CLK, RN => RST, Q => 
                           n_4218, QN => n3152);
   clk_r_REG6874_S6 : DFFR_X1 port map( D => n4049, CK => CLK, RN => RST, Q => 
                           n_4219, QN => n3151);
   clk_r_REG4234_S5 : DFFR_X1 port map( D => n2350, CK => CLK, RN => RST, Q => 
                           n3150, QN => n_4220);
   clk_r_REG4490_S3 : DFFS_X1 port map( D => n2398, CK => CLK, SN => RST, Q => 
                           n3149, QN => n_4221);
   clk_r_REG4256_S6 : DFFR_X1 port map( D => n1346, CK => CLK, RN => RST, Q => 
                           n3148, QN => n_4222);
   clk_r_REG4579_S5 : DFFR_X1 port map( D => n1345, CK => CLK, RN => RST, Q => 
                           n3147, QN => n_4223);
   clk_r_REG4243_S9 : DFFR_X1 port map( D => n1344, CK => CLK, RN => RST, Q => 
                           n3146, QN => n_4224);
   clk_r_REG4692_S6 : DFFR_X1 port map( D => n1343, CK => CLK, RN => RST, Q => 
                           n3145, QN => n_4225);
   clk_r_REG4683_S6 : DFFR_X1 port map( D => n1342, CK => CLK, RN => RST, Q => 
                           n3144, QN => n_4226);
   clk_r_REG4674_S6 : DFFR_X1 port map( D => n1341, CK => CLK, RN => RST, Q => 
                           n3143, QN => n_4227);
   clk_r_REG4665_S7 : DFFR_X1 port map( D => n1340, CK => CLK, RN => RST, Q => 
                           n3142, QN => n_4228);
   clk_r_REG4657_S6 : DFFR_X1 port map( D => n1339, CK => CLK, RN => RST, Q => 
                           n3141, QN => n_4229);
   clk_r_REG4650_S6 : DFFR_X1 port map( D => n1338, CK => CLK, RN => RST, Q => 
                           n3140, QN => n_4230);
   clk_r_REG4644_S6 : DFFR_X1 port map( D => n1337, CK => CLK, RN => RST, Q => 
                           n3139, QN => n_4231);
   clk_r_REG4638_S6 : DFFR_X1 port map( D => n1336, CK => CLK, RN => RST, Q => 
                           n3138, QN => n_4232);
   clk_r_REG4629_S7 : DFFR_X1 port map( D => n1335, CK => CLK, RN => RST, Q => 
                           n3137, QN => n_4233);
   clk_r_REG4623_S7 : DFFR_X1 port map( D => n1334, CK => CLK, RN => RST, Q => 
                           n3136, QN => n_4234);
   clk_r_REG6780_S1 : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK => CLK, 
                           RN => RST, Q => n3134, QN => n_4235);
   clk_r_REG4855_S5 : DFFS_X1 port map( D => n2478, CK => CLK, SN => RST, Q => 
                           n3133, QN => n_4236);
   clk_r_REG4578_S5 : DFFS_X1 port map( D => n1325, CK => CLK, SN => RST, Q => 
                           n3132, QN => n_4237);
   clk_r_REG4005_S8 : DFFS_X1 port map( D => n1324, CK => CLK, SN => RST, Q => 
                           n3131, QN => n_4238);
   clk_r_REG4249_S9 : DFFS_X1 port map( D => n1323, CK => CLK, SN => RST, Q => 
                           n3130, QN => n_4239);
   clk_r_REG4008_S9 : DFFS_X1 port map( D => n1322, CK => CLK, SN => RST, Q => 
                           n3129, QN => n_4240);
   clk_r_REG4016_S6 : DFFS_X1 port map( D => n1321, CK => CLK, SN => RST, Q => 
                           n3128, QN => n_4241);
   clk_r_REG4022_S6 : DFFS_X1 port map( D => n1320, CK => CLK, SN => RST, Q => 
                           n3127, QN => n_4242);
   clk_r_REG4028_S13 : DFFS_X1 port map( D => n1319, CK => CLK, SN => RST, Q =>
                           n3126, QN => n_4243);
   clk_r_REG4034_S13 : DFFS_X1 port map( D => n1318, CK => CLK, SN => RST, Q =>
                           n3125, QN => n_4244);
   clk_r_REG4040_S7 : DFFS_X1 port map( D => n1317, CK => CLK, SN => RST, Q => 
                           n3124, QN => n_4245);
   clk_r_REG4584_S6 : DFFS_X1 port map( D => n1316, CK => CLK, SN => RST, Q => 
                           n3123, QN => n_4246);
   clk_r_REG4590_S13 : DFFS_X1 port map( D => n1315, CK => CLK, SN => RST, Q =>
                           n3122, QN => n_4247);
   clk_r_REG4596_S7 : DFFS_X1 port map( D => n1314, CK => CLK, SN => RST, Q => 
                           n3121, QN => n_4248);
   clk_r_REG4602_S13 : DFFS_X1 port map( D => n1313, CK => CLK, SN => RST, Q =>
                           n3120, QN => n_4249);
   clk_r_REG4610_S7 : DFFS_X1 port map( D => n1312, CK => CLK, SN => RST, Q => 
                           n3119, QN => n_4250);
   clk_r_REG3641_S3 : DFFS_X1 port map( D => n4040, CK => CLK, SN => RST, Q => 
                           n_4251, QN => n3118);
   clk_r_REG5929_S4 : DFFR_X1 port map( D => n3118, CK => CLK, RN => RST, Q => 
                           n3117, QN => n4420);
   clk_r_REG4998_S5 : DFFR_X1 port map( D => n1330, CK => CLK, RN => RST, Q => 
                           n3116, QN => n3672);
   clk_r_REG5933_S5 : DFFS_X1 port map( D => n3115, CK => CLK, SN => RST, Q => 
                           n3114, QN => n_4252);
   clk_r_REG6713_S3 : DFFR_X1 port map( D => n1302, CK => CLK, RN => RST, Q => 
                           n3113, QN => n_4253);
   clk_r_REG6714_S4 : DFFR_X1 port map( D => n3113, CK => CLK, RN => RST, Q => 
                           n3112, QN => n_4254);
   clk_r_REG6662_S3 : DFFR_X1 port map( D => n302, CK => CLK, RN => RST, Q => 
                           n3111, QN => n_4255);
   clk_r_REG4042_S5 : DFFR_X1 port map( D => n4086, CK => CLK, RN => RST, Q => 
                           n_4256, QN => n3110);
   clk_r_REG4041_S5 : DFFS_X1 port map( D => n4086, CK => CLK, SN => RST, Q => 
                           n_4257, QN => n3109);
   clk_r_REG4036_S5 : DFFR_X1 port map( D => n4085, CK => CLK, RN => RST, Q => 
                           n_4258, QN => n3108);
   clk_r_REG4035_S5 : DFFS_X1 port map( D => n4085, CK => CLK, SN => RST, Q => 
                           n_4259, QN => n3107);
   clk_r_REG4030_S6 : DFFR_X1 port map( D => n4084, CK => CLK, RN => RST, Q => 
                           n_4260, QN => n3106);
   clk_r_REG4029_S6 : DFFS_X1 port map( D => n4084, CK => CLK, SN => RST, Q => 
                           n_4261, QN => n3105);
   clk_r_REG4018_S5 : DFFR_X1 port map( D => n4083, CK => CLK, RN => RST, Q => 
                           n_4262, QN => n3104);
   clk_r_REG4017_S5 : DFFS_X1 port map( D => n4083, CK => CLK, SN => RST, Q => 
                           n_4263, QN => n3103);
   clk_r_REG4024_S5 : DFFR_X1 port map( D => n4082, CK => CLK, RN => RST, Q => 
                           n_4264, QN => n3102);
   clk_r_REG4023_S5 : DFFS_X1 port map( D => n4082, CK => CLK, SN => RST, Q => 
                           n_4265, QN => n3101);
   clk_r_REG4586_S5 : DFFR_X1 port map( D => n4081, CK => CLK, RN => RST, Q => 
                           n_4266, QN => n3100);
   clk_r_REG4585_S5 : DFFS_X1 port map( D => n4081, CK => CLK, SN => RST, Q => 
                           n_4267, QN => n3099);
   clk_r_REG4592_S5 : DFFR_X1 port map( D => n4080, CK => CLK, RN => RST, Q => 
                           n_4268, QN => n3098);
   clk_r_REG4591_S5 : DFFS_X1 port map( D => n4080, CK => CLK, SN => RST, Q => 
                           n_4269, QN => n3097);
   clk_r_REG4231_S5 : DFFR_X1 port map( D => n4116, CK => CLK, RN => RST, Q => 
                           n_4270, QN => n3096);
   clk_r_REG4241_S5 : DFFR_X1 port map( D => n4115, CK => CLK, RN => RST, Q => 
                           n_4271, QN => n3095);
   clk_r_REG4240_S5 : DFFS_X1 port map( D => n4115, CK => CLK, SN => RST, Q => 
                           n_4272, QN => n3094);
   clk_r_REG4012_S5 : DFFR_X1 port map( D => n4114, CK => CLK, RN => RST, Q => 
                           n_4273, QN => n3093);
   clk_r_REG4011_S5 : DFFS_X1 port map( D => n4114, CK => CLK, SN => RST, Q => 
                           n_4274, QN => n3092);
   clk_r_REG4598_S6 : DFFR_X1 port map( D => n4079, CK => CLK, RN => RST, Q => 
                           n_4275, QN => n3091);
   clk_r_REG4597_S6 : DFFS_X1 port map( D => n4079, CK => CLK, SN => RST, Q => 
                           n_4276, QN => n3090);
   clk_r_REG4604_S6 : DFFR_X1 port map( D => n4078, CK => CLK, RN => RST, Q => 
                           n_4277, QN => n3089);
   clk_r_REG4603_S6 : DFFS_X1 port map( D => n4078, CK => CLK, SN => RST, Q => 
                           n_4278, QN => n3088);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => n3580, ADD_WR(3) => n3584, ADD_WR(2) =>
                           n3112, ADD_WR(1) => n3582, ADD_WR(0) => n3578, 
                           ADD_RD1(4) => n1415, ADD_RD1(3) => n1414, ADD_RD1(2)
                           => n1413, ADD_RD1(1) => n1412, ADD_RD1(0) => n1411, 
                           ADD_RD2(4) => curr_instruction_to_cu_i_20_port, 
                           ADD_RD2(3) => curr_instruction_to_cu_i_19_port, 
                           ADD_RD2(2) => n4113, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n43, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n44, OUT1(31) => n1673, 
                           OUT1(30) => n1671, OUT1(29) => n1669, OUT1(28) => 
                           n1667, OUT1(27) => n1665, OUT1(26) => n1663, 
                           OUT1(25) => n1661, OUT1(24) => n1659, OUT1(23) => 
                           n1657, OUT1(22) => n1655, OUT1(21) => n1653, 
                           OUT1(20) => n1651, OUT1(19) => n1649, OUT1(18) => 
                           n1647, OUT1(17) => n1645, OUT1(16) => n1643, 
                           OUT1(15) => n1641, OUT1(14) => n1639, OUT1(13) => 
                           n1637, OUT1(12) => n1635, OUT1(11) => n1633, 
                           OUT1(10) => n1631, OUT1(9) => n1629, OUT1(8) => 
                           n1627, OUT1(7) => n1625, OUT1(6) => n1623, OUT1(5) 
                           => n1621, OUT1(4) => n1619, OUT1(3) => n1617, 
                           OUT1(2) => n1615, OUT1(1) => n1614, OUT1(0) => n1613
                           , OUT2(31) => n1611, OUT2(30) => n1608, OUT2(29) => 
                           n1605, OUT2(28) => n1602, OUT2(27) => n1599, 
                           OUT2(26) => n1596, OUT2(25) => n1593, OUT2(24) => 
                           n1590, OUT2(23) => n1587, OUT2(22) => n1584, 
                           OUT2(21) => n1581, OUT2(20) => n1578, OUT2(19) => 
                           n1575, OUT2(18) => n1572, OUT2(17) => n1569, 
                           OUT2(16) => n1566, OUT2(15) => n1563, OUT2(14) => 
                           n1560, OUT2(13) => n1557, OUT2(12) => n1554, 
                           OUT2(11) => n1551, OUT2(10) => n1548, OUT2(9) => 
                           n1545, OUT2(8) => n1542, OUT2(7) => n1539, OUT2(6) 
                           => n1536, OUT2(5) => n1533, OUT2(4) => n1530, 
                           OUT2(3) => n1527, OUT2(2) => n1524, OUT2(1) => n1521
                           , OUT2(0) => n1518, RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_4279, mul_exeception => 
                           n_4280, FUNC(0) => n4033, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_4281, 
                           OUTALU(31) => datapath_i_alu_output_val_i_31_port, 
                           OUTALU(30) => datapath_i_alu_output_val_i_30_port, 
                           OUTALU(29) => datapath_i_alu_output_val_i_29_port, 
                           OUTALU(28) => datapath_i_alu_output_val_i_28_port, 
                           OUTALU(27) => datapath_i_alu_output_val_i_27_port, 
                           OUTALU(26) => datapath_i_alu_output_val_i_26_port, 
                           OUTALU(25) => datapath_i_alu_output_val_i_25_port, 
                           OUTALU(24) => datapath_i_alu_output_val_i_24_port, 
                           OUTALU(23) => datapath_i_alu_output_val_i_23_port, 
                           OUTALU(22) => datapath_i_alu_output_val_i_22_port, 
                           OUTALU(21) => datapath_i_alu_output_val_i_21_port, 
                           OUTALU(20) => datapath_i_alu_output_val_i_20_port, 
                           OUTALU(19) => datapath_i_alu_output_val_i_19_port, 
                           OUTALU(18) => datapath_i_alu_output_val_i_18_port, 
                           OUTALU(17) => datapath_i_alu_output_val_i_17_port, 
                           OUTALU(16) => datapath_i_alu_output_val_i_16_port, 
                           OUTALU(15) => datapath_i_alu_output_val_i_15_port, 
                           OUTALU(14) => datapath_i_alu_output_val_i_14_port, 
                           OUTALU(13) => datapath_i_alu_output_val_i_13_port, 
                           OUTALU(12) => datapath_i_alu_output_val_i_12_port, 
                           OUTALU(11) => datapath_i_alu_output_val_i_11_port, 
                           OUTALU(10) => datapath_i_alu_output_val_i_10_port, 
                           OUTALU(9) => datapath_i_alu_output_val_i_9_port, 
                           OUTALU(8) => datapath_i_alu_output_val_i_8_port, 
                           OUTALU(7) => datapath_i_alu_output_val_i_7_port, 
                           OUTALU(6) => datapath_i_alu_output_val_i_6_port, 
                           OUTALU(5) => datapath_i_alu_output_val_i_5_port, 
                           OUTALU(4) => datapath_i_alu_output_val_i_4_port, 
                           OUTALU(3) => datapath_i_alu_output_val_i_3_port, 
                           OUTALU(2) => datapath_i_alu_output_val_i_2_port, 
                           OUTALU(1) => datapath_i_alu_output_val_i_1_port, 
                           OUTALU(0) => datapath_i_alu_output_val_i_0_port, 
                           rst_BAR => RST);
   U1672 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_31_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(31), ZN => n3857
                           );
   U1674 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_30_port, A2 => 
                           n4433, B1 => n4434, B2 => DRAM_DATA(30), ZN => n3858
                           );
   U1676 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_29_port, A2 => 
                           n3889, B1 => n4434, B2 => DRAM_DATA(29), ZN => n3859
                           );
   U1678 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_28_port, A2 => 
                           n3889, B1 => n4434, B2 => DRAM_DATA(28), ZN => n3860
                           );
   U1680 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_27_port, A2 => 
                           n4433, B1 => n4434, B2 => DRAM_DATA(27), ZN => n3861
                           );
   U1682 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_26_port, A2 => 
                           n3889, B1 => n4434, B2 => DRAM_DATA(26), ZN => n3862
                           );
   U1684 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_25_port, A2 => 
                           n4433, B1 => n4434, B2 => DRAM_DATA(25), ZN => n3863
                           );
   U1686 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_24_port, A2 => 
                           n4433, B1 => n4434, B2 => DRAM_DATA(24), ZN => n3864
                           );
   U1688 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_23_port, A2 => 
                           n4433, B1 => n4434, B2 => DRAM_DATA(23), ZN => n3865
                           );
   U1690 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_22_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(22), ZN => n3866
                           );
   U1692 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_21_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(21), ZN => n3867
                           );
   U1694 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_20_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(20), ZN => n3868
                           );
   U1696 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_19_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(19), ZN => n3869
                           );
   U1698 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_18_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(18), ZN => n3870
                           );
   U1700 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_17_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(17), ZN => n3871
                           );
   U1702 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(16), B1 => n4433, B2
                           => datapath_i_alu_output_val_i_16_port, ZN => n3872)
                           ;
   U1704 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(15), B1 => n4433, B2
                           => datapath_i_alu_output_val_i_15_port, ZN => n3873)
                           ;
   U1706 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(14), B1 => n4433, B2
                           => datapath_i_alu_output_val_i_14_port, ZN => n3874)
                           ;
   U1708 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(13), B1 => n4433, B2
                           => datapath_i_alu_output_val_i_13_port, ZN => n3875)
                           ;
   U1710 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(12), B1 => n4433, B2
                           => datapath_i_alu_output_val_i_12_port, ZN => n3876)
                           ;
   U1712 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(11), B1 => n4433, B2
                           => datapath_i_alu_output_val_i_11_port, ZN => n3877)
                           ;
   U1714 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(10), B1 => n4433, B2
                           => datapath_i_alu_output_val_i_10_port, ZN => n3878)
                           ;
   U1716 : AOI22_X1 port map( A1 => n3888, A2 => DRAM_DATA(9), B1 => n4433, B2 
                           => datapath_i_alu_output_val_i_9_port, ZN => n3879);
   U1718 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_8_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(8), ZN => n3880)
                           ;
   U1720 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_7_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(7), ZN => n3881)
                           ;
   U1722 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_6_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(6), ZN => n3882)
                           ;
   U1724 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_5_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(5), ZN => n3883)
                           ;
   U1726 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_4_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(4), ZN => n3884)
                           ;
   U1728 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_3_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(3), ZN => n3885)
                           ;
   U1730 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_2_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(2), ZN => n3886)
                           ;
   U1732 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_1_port, A2 => 
                           n3889, B1 => n3888, B2 => DRAM_DATA(1), ZN => n3887)
                           ;
   U1734 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_0_port, A2 => 
                           n4433, B1 => n3888, B2 => DRAM_DATA(0), ZN => n3890)
                           ;
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   clk_r_REG4617_S6 : DFFR_X1 port map( D => n1916, CK => CLK, RN => RST, Q => 
                           n3692, QN => n_4282);
   clk_r_REG6706_S3 : DFFS_X1 port map( D => n1497, CK => CLK, SN => RST, Q => 
                           n3576, QN => n_4283);
   clk_r_REG6194_S2 : DFF_X1 port map( D => n1673, CK => CLK, Q => n3441, QN =>
                           n_4284);
   clk_r_REG5928_S4 : DFFS_X1 port map( D => n3258, CK => CLK, SN => RST, Q => 
                           n3257, QN => n4425);
   clk_r_REG6705_S3 : DFFS_X1 port map( D => n1497, CK => CLK, SN => RST, Q => 
                           n3254, QN => n4422);
   clk_r_REG6773_S5 : DFFR_X1 port map( D => n1727, CK => CLK, RN => RST, Q => 
                           n3241, QN => n_4285);
   clk_r_REG6661_S3 : DFFS_X1 port map( D => n1728, CK => CLK, SN => RST, Q => 
                           n3135, QN => n_4286);
   clk_r_REG6725_S3 : DFFR_X1 port map( D => n4432, CK => CLK, RN => RST, Q => 
                           n3587, QN => n_4287);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => n3235, Q => 
                           n1801);
   clk_r_REG6885_S6 : DFFR_X1 port map( D => n1405, CK => CLK, RN => RST, Q => 
                           n3229, QN => n_4288);
   clk_r_REG5931_S4 : DFFR_X1 port map( D => n4042, CK => CLK, RN => RST, Q => 
                           n3554, QN => n_4289);
   clk_r_REG5930_S4 : DFFR_X1 port map( D => n4042, CK => CLK, RN => RST, Q => 
                           n_4290, QN => n3115);
   clk_r_REG3644_S4 : DFFR_X1 port map( D => n3654, CK => CLK, RN => RST, Q => 
                           n_4291, QN => n3255);
   clk_r_REG6771_S5 : DFFS_X1 port map( D => n1507, CK => CLK, SN => RST, Q => 
                           n3261, QN => n_4292);
   clk_r_REG6776_S3 : DFFR_X1 port map( D => n4043, CK => CLK, RN => RST, Q => 
                           n_4293, QN => n3156);
   clk_r_REG6787_S5 : DFFS_X1 port map( D => n4047, CK => CLK, SN => RST, Q => 
                           n_4294, QN => n3278);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X2 port map( A => 
                           n3335, EN => n3254, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X2 port map( A => 
                           n3326, EN => n3576, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X2 port map( A => 
                           n3329, EN => n4431, Z => DRAM_DATA(14));
   clk_r_REG6716_S5 : DFFS_X2 port map( D => n3658, CK => CLK, SN => RST, Q => 
                           n3596, QN => n_4295);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X2 port map( A => 
                           n3332, EN => n3576, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X2 port map( A => 
                           n3320, EN => n3576, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X2 port map( A => 
                           n3314, EN => n3576, Z => DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X2 port map( A => 
                           n3323, EN => n4431, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X2 port map( A => 
                           n3317, EN => n4431, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X2 port map( A => 
                           n3377, EN => n3576, Z => DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X2 port map( A => 
                           n3371, EN => n3576, Z => DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X2 port map( A => 
                           n3365, EN => n3576, Z => DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X2 port map( A => 
                           n3359, EN => n3576, Z => DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X2 port map( A => 
                           n3353, EN => n3576, Z => DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X2 port map( A => 
                           n3311, EN => n3576, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X2 port map( A => 
                           n3287, EN => n3576, Z => DRAM_DATA(0));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X2 port map( A => 
                           n3380, EN => n3254, Z => DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X2 port map( A => 
                           n3374, EN => n3254, Z => DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X2 port map( A => 
                           n3368, EN => n3254, Z => DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X2 port map( A => 
                           n3356, EN => n3254, Z => DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X2 port map( A => 
                           n3350, EN => n3254, Z => DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X2 port map( A => 
                           n3347, EN => n3254, Z => DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X2 port map( A => 
                           n3344, EN => n3254, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X2 port map( A => 
                           n3341, EN => n3254, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X2 port map( A => 
                           n3308, EN => n3254, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X2 port map( A => 
                           n3302, EN => n3254, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X2 port map( A => 
                           n3299, EN => n3254, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X2 port map( A => 
                           n3362, EN => n4431, Z => DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X2 port map( A => 
                           n3338, EN => n4431, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X2 port map( A => 
                           n3305, EN => n4431, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X2 port map( A => 
                           n3296, EN => n4431, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X2 port map( A => 
                           n3293, EN => n4431, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X2 port map( A => 
                           n3290, EN => n4431, Z => DRAM_DATA(1));
   U1952 : OAI21_X2 port map( B1 => n3261, B2 => n3496, A => n4274, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U1953 : OAI21_X2 port map( B1 => n3559, B2 => n3492, A => n4280, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U1954 : OAI21_X2 port map( B1 => n3559, B2 => n3469, A => n4270, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U1955 : OAI21_X2 port map( B1 => n3261, B2 => n3465, A => n4278, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U1956 : OAI21_X2 port map( B1 => n3559, B2 => n3474, A => n4261, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U1957 : CLKBUF_X1 port map( A => n3692, Z => n4132);
   U1958 : AOI22_X1 port map( A1 => n3278, A2 => cu_i_cmd_alu_op_type_3_port, 
                           B1 => n3456, B2 => n3285, ZN => n4203);
   U1959 : AOI22_X1 port map( A1 => n3278, A2 => cu_i_cmd_alu_op_type_2_port, 
                           B1 => n3456, B2 => n3286, ZN => n4204);
   U1960 : AOI22_X1 port map( A1 => n3278, A2 => cu_i_cmd_alu_op_type_0_port, 
                           B1 => n3456, B2 => n3280, ZN => n4207);
   U1961 : CLKBUF_X1 port map( A => n3135, Z => n4379);
   U1962 : CLKBUF_X1 port map( A => n3587, Z => n4378);
   U1963 : NOR2_X1 port map( A1 => n4204, A2 => n4205, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U1964 : MUX2_X1 port map( A => n3168, B => n3300, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U1965 : MUX2_X1 port map( A => IRAM_DATA(23), B => n3205, S => n3278, Z => 
                           n1413);
   U1966 : INV_X1 port map( A => n1801, ZN => n4047);
   U1967 : NOR2_X1 port map( A1 => n1801, A2 => n3272, ZN => n4188);
   U1968 : AOI21_X1 port map( B1 => n1801, B2 => n3527, A => n4188, ZN => n4133
                           );
   U1969 : INV_X1 port map( A => n4133, ZN => n4041);
   U1970 : AOI22_X1 port map( A1 => n3278, A2 => n3535, B1 => n3552, B2 => 
                           IRAM_DATA(13), ZN => n4364);
   U1971 : INV_X1 port map( A => n4364, ZN => n4112);
   U1972 : AOI22_X1 port map( A1 => n3555, A2 => n3538, B1 => n3593, B2 => 
                           IRAM_DATA(1), ZN => n4326);
   U1973 : INV_X1 port map( A => n4326, ZN => n4050);
   U1974 : AOI22_X1 port map( A1 => n3555, A2 => n3537, B1 => n3593, B2 => 
                           IRAM_DATA(2), ZN => n4328);
   U1975 : INV_X1 port map( A => n4328, ZN => n4051);
   U1976 : AOI22_X1 port map( A1 => n3555, A2 => n3530, B1 => n3593, B2 => 
                           IRAM_DATA(29), ZN => n4362);
   U1977 : INV_X1 port map( A => n4362, ZN => n4065);
   U1978 : AOI22_X1 port map( A1 => n3555, A2 => n3529, B1 => n3593, B2 => 
                           IRAM_DATA(30), ZN => n4144);
   U1979 : INV_X1 port map( A => n4144, ZN => n4062);
   U1980 : AOI22_X1 port map( A1 => n3555, A2 => n3528, B1 => n3593, B2 => 
                           IRAM_DATA(31), ZN => n4162);
   U1981 : NAND3_X1 port map( A1 => n4065, A2 => n4062, A3 => n4162, ZN => 
                           n4136);
   U1982 : INV_X1 port map( A => n4136, ZN => n1500);
   U1983 : AOI22_X1 port map( A1 => n3278, A2 => n3534, B1 => n3552, B2 => 
                           IRAM_DATA(18), ZN => n4366);
   U1984 : INV_X1 port map( A => n4366, ZN => n4113);
   U1985 : AOI22_X1 port map( A1 => n3555, A2 => n3531, B1 => n3593, B2 => 
                           IRAM_DATA(28), ZN => n4327);
   U1986 : INV_X1 port map( A => n4327, ZN => n4061);
   U1987 : AOI22_X1 port map( A1 => n3555, A2 => n3533, B1 => n3593, B2 => 
                           IRAM_DATA(26), ZN => n4414);
   U1988 : INV_X1 port map( A => n4414, ZN => n4064);
   U1989 : INV_X1 port map( A => n4162, ZN => n4063);
   U1990 : AOI22_X1 port map( A1 => n3555, A2 => n3532, B1 => n3593, B2 => 
                           IRAM_DATA(27), ZN => n4332);
   U1991 : NOR3_X1 port map( A1 => n4332, A2 => n4062, A3 => n4061, ZN => n4138
                           );
   U1992 : NAND3_X1 port map( A1 => n4138, A2 => n4064, A3 => n4063, ZN => 
                           n4164);
   U1993 : NOR2_X1 port map( A1 => n4421, A2 => n4164, ZN => n4056);
   U1994 : INV_X1 port map( A => n4056, ZN => n4361);
   U1995 : NOR2_X1 port map( A1 => n4065, A2 => n4361, ZN => 
                           cu_i_cmd_word_3_port);
   U1996 : NAND2_X1 port map( A1 => n4332, A2 => n4414, ZN => n4055);
   U1997 : INV_X1 port map( A => n4055, ZN => n4161);
   U1998 : NOR2_X1 port map( A1 => n4065, A2 => n4063, ZN => n4143);
   U1999 : NAND4_X1 port map( A1 => n4161, A2 => n4143, A3 => n4144, A4 => 
                           n4327, ZN => n4053);
   U2000 : NOR2_X1 port map( A1 => n4053, A2 => n4421, ZN => n4054);
   U2001 : NOR2_X1 port map( A1 => n3555, A2 => IRAM_DATA(0), ZN => n4134);
   U2002 : AOI21_X1 port map( B1 => n3664, B2 => n3555, A => n4134, ZN => n1390
                           );
   U2003 : MUX2_X1 port map( A => IRAM_DATA(3), B => n3236, S => n3555, Z => 
                           n1393);
   U2004 : MUX2_X1 port map( A => IRAM_DATA(4), B => n3238, S => n3555, Z => 
                           n1394);
   U2005 : AOI22_X1 port map( A1 => n3555, A2 => n3536, B1 => n3593, B2 => 
                           IRAM_DATA(5), ZN => n4135);
   U2006 : INV_X1 port map( A => n4135, ZN => n4049);
   U2007 : INV_X1 port map( A => n4332, ZN => n4058);
   U2008 : AOI211_X1 port map( C1 => n4327, C2 => n4414, A => n4058, B => n4136
                           , ZN => n4060);
   U2009 : NAND2_X1 port map( A1 => n4143, A2 => n4061, ZN => n4137);
   U2010 : NOR3_X1 port map( A1 => n4144, A2 => n4064, A3 => n4137, ZN => n1350
                           );
   U2011 : AND2_X1 port map( A1 => n4143, A2 => n4138, ZN => n4165);
   U2012 : NAND2_X1 port map( A1 => n3277, A2 => n4165, ZN => n4363);
   U2013 : INV_X1 port map( A => n4054, ZN => n4329);
   U2014 : NAND4_X1 port map( A1 => n1390, A2 => n1393, A3 => n1394, A4 => 
                           n4049, ZN => n4139);
   U2015 : NOR3_X1 port map( A1 => n4326, A2 => n4328, A3 => n4139, ZN => n4190
                           );
   U2016 : NOR3_X1 port map( A1 => n4362, A2 => n4063, A3 => n4062, ZN => n4415
                           );
   U2017 : OAI21_X1 port map( B1 => n4327, B2 => n4058, A => n4064, ZN => n4140
                           );
   U2018 : AOI211_X1 port map( C1 => n4415, C2 => n4140, A => n4060, B => n1350
                           , ZN => n4240);
   U2019 : OAI222_X1 port map( A1 => n4363, A2 => n4414, B1 => n4329, B2 => 
                           n4190, C1 => n4240, C2 => n3589, ZN => n302);
   U2020 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n302, ZN => n1498
                           );
   U2021 : OAI22_X1 port map( A1 => n4047, A2 => cu_i_cmd_word_3_port, B1 => 
                           n3211, B2 => n1801, ZN => n4301);
   U2022 : INV_X1 port map( A => n4301, ZN => n4045);
   U2023 : OAI22_X1 port map( A1 => n4047, A2 => n4056, B1 => n3210, B2 => 
                           n1801, ZN => n1760);
   U2024 : INV_X1 port map( A => n1760, ZN => n4044);
   U2025 : NAND2_X1 port map( A1 => n3224, A2 => n3263, ZN => n4234);
   U2026 : NOR2_X1 port map( A1 => n3093, A2 => n4234, ZN => n4233);
   U2027 : NAND2_X1 port map( A1 => n4233, A2 => n3223, ZN => n4231);
   U2028 : NOR2_X1 port map( A1 => n3104, A2 => n4231, ZN => n4230);
   U2029 : NAND2_X1 port map( A1 => n4230, A2 => n3222, ZN => n4228);
   U2030 : NOR2_X1 port map( A1 => n3102, A2 => n4228, ZN => n4227);
   U2031 : NAND2_X1 port map( A1 => n4227, A2 => n3221, ZN => n4225);
   U2032 : OAI211_X1 port map( C1 => n4227, C2 => n3221, A => n3553, B => n4225
                           , ZN => n4141);
   U2033 : NAND2_X1 port map( A1 => n3126, A2 => n4141, ZN => n4271);
   U2034 : INV_X1 port map( A => n4271, ZN => n4102);
   U2035 : INV_X1 port map( A => datapath_i_alu_output_val_i_16_port, ZN => 
                           n4142);
   U2036 : OAI222_X1 port map( A1 => n4142, A2 => n4419, B1 => n3255, B2 => 
                           n3498, C1 => n4425, C2 => n4102, ZN => n1441);
   U2037 : INV_X1 port map( A => n1441, ZN => n4094);
   U2038 : NAND4_X1 port map( A1 => n4144, A2 => n4143, A3 => n3277, A4 => 
                           n4061, ZN => n4145);
   U2039 : OAI21_X1 port map( B1 => n4055, B2 => n4145, A => n4363, ZN => 
                           cu_i_cmd_word_6_port);
   U2040 : NAND2_X1 port map( A1 => n4332, A2 => n4064, ZN => n474);
   U2041 : OAI221_X1 port map( B1 => n1801, B2 => n3240, C1 => n4047, C2 => 
                           cu_i_cmd_word_6_port, A => n3242, ZN => n4147);
   U2042 : NOR2_X1 port map( A1 => n4145, A2 => n474, ZN => n4187);
   U2043 : AOI22_X1 port map( A1 => n1801, A2 => n4187, B1 => n3273, B2 => 
                           n4047, ZN => n4146);
   U2044 : MUX2_X1 port map( A => n3242, B => n4147, S => n4146, Z => n4040);
   U2045 : NOR2_X1 port map( A1 => n3106, A2 => n4225, ZN => n4224);
   U2046 : NAND2_X1 port map( A1 => n4224, A2 => n3220, ZN => n4222);
   U2047 : OAI211_X1 port map( C1 => n4224, C2 => n3220, A => n3553, B => n4222
                           , ZN => n4148);
   U2048 : NAND2_X1 port map( A1 => n3125, A2 => n4148, ZN => n4262);
   U2049 : INV_X1 port map( A => n4262, ZN => n4099);
   U2050 : INV_X1 port map( A => datapath_i_alu_output_val_i_18_port, ZN => 
                           n4149);
   U2051 : OAI222_X1 port map( A1 => n4149, A2 => n4419, B1 => n3255, B2 => 
                           n3500, C1 => n4425, C2 => n4099, ZN => n1439);
   U2052 : INV_X1 port map( A => n1439, ZN => n4093);
   U2053 : NOR2_X1 port map( A1 => n1512, A2 => n1513, ZN => n4150);
   U2054 : NAND3_X1 port map( A1 => n1510, A2 => n4150, A3 => cu_i_n151, ZN => 
                           n1458);
   U2055 : INV_X1 port map( A => cu_i_n151, ZN => n4039);
   U2056 : OR2_X1 port map( A1 => n4150, A2 => n4039, ZN => n4038);
   U2057 : MUX2_X1 port map( A => IRAM_DATA(16), B => n3228, S => n3278, Z => 
                           curr_instruction_to_cu_i_16_port);
   U2058 : MUX2_X1 port map( A => IRAM_DATA(11), B => n3227, S => n3555, Z => 
                           n1401);
   U2059 : INV_X1 port map( A => n4363, ZN => n4057);
   U2060 : CLKBUF_X1 port map( A => n4057, Z => n4432);
   U2061 : NAND2_X1 port map( A1 => n1458, A2 => n4038, ZN => n4191);
   U2062 : AOI21_X1 port map( B1 => n4191, B2 => n4190, A => n4329, ZN => n4367
                           );
   U2063 : INV_X1 port map( A => n4367, ZN => n4365);
   U2064 : AOI221_X1 port map( B1 => n4365, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n4367, C2 =>
                           n1401, A => n4432, ZN => n4151);
   U2065 : INV_X1 port map( A => n4151, ZN => n4034);
   U2066 : MUX2_X1 port map( A => IRAM_DATA(20), B => n3230, S => n3278, Z => 
                           curr_instruction_to_cu_i_20_port);
   U2067 : MUX2_X1 port map( A => IRAM_DATA(15), B => n3229, S => n3278, Z => 
                           n1405);
   U2068 : AOI221_X1 port map( B1 => n4365, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n4367, C2 =>
                           n1405, A => n4432, ZN => n4152);
   U2069 : INV_X1 port map( A => n4152, ZN => n4035);
   U2070 : MUX2_X1 port map( A => IRAM_DATA(19), B => n3234, S => n3278, Z => 
                           curr_instruction_to_cu_i_19_port);
   U2071 : MUX2_X1 port map( A => IRAM_DATA(14), B => n3233, S => n3278, Z => 
                           n1404);
   U2072 : AOI221_X1 port map( B1 => n4365, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n4367, C2 =>
                           n1404, A => n4432, ZN => n4153);
   U2073 : INV_X1 port map( A => n4153, ZN => n4037);
   U2074 : MUX2_X1 port map( A => IRAM_DATA(17), B => n3232, S => n3278, Z => 
                           curr_instruction_to_cu_i_17_port);
   U2075 : MUX2_X1 port map( A => IRAM_DATA(12), B => n3231, S => n3278, Z => 
                           n1402);
   U2076 : AOI221_X1 port map( B1 => n4365, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n4367, C2 =>
                           n1402, A => n4432, ZN => n4154);
   U2077 : INV_X1 port map( A => n4154, ZN => n4036);
   U2078 : OAI211_X1 port map( C1 => n4233, C2 => n3223, A => n3553, B => n4231
                           , ZN => n4155);
   U2079 : NAND2_X1 port map( A1 => n3128, A2 => n4155, ZN => n4275);
   U2080 : INV_X1 port map( A => n4275, ZN => n4100);
   U2081 : INV_X1 port map( A => datapath_i_alu_output_val_i_12_port, ZN => 
                           n4156);
   U2082 : OAI222_X1 port map( A1 => n4156, A2 => n4420, B1 => n3255, B2 => 
                           n3494, C1 => n4425, C2 => n4100, ZN => n1445);
   U2083 : INV_X1 port map( A => n1445, ZN => n4101);
   U2084 : OAI211_X1 port map( C1 => n4230, C2 => n3222, A => n3553, B => n4228
                           , ZN => n4157);
   U2085 : NAND2_X1 port map( A1 => n3127, A2 => n4157, ZN => n4273);
   U2086 : INV_X1 port map( A => n4273, ZN => n4106);
   U2087 : INV_X1 port map( A => datapath_i_alu_output_val_i_14_port, ZN => 
                           n4158);
   U2088 : OAI222_X1 port map( A1 => n4158, A2 => n4419, B1 => n3255, B2 => 
                           n3496, C1 => n4425, C2 => n4106, ZN => n1443);
   U2089 : INV_X1 port map( A => n1443, ZN => n4095);
   U2090 : NOR2_X1 port map( A1 => n3108, A2 => n4222, ZN => n4221);
   U2091 : NAND2_X1 port map( A1 => n4221, A2 => n3219, ZN => n4219);
   U2092 : OAI211_X1 port map( C1 => n4221, C2 => n3219, A => n3553, B => n4219
                           , ZN => n4159);
   U2093 : NAND2_X1 port map( A1 => n3124, A2 => n4159, ZN => n4292);
   U2094 : INV_X1 port map( A => n4292, ZN => n4105);
   U2095 : INV_X1 port map( A => datapath_i_alu_output_val_i_20_port, ZN => 
                           n4160);
   U2096 : OAI222_X1 port map( A1 => n4160, A2 => n4419, B1 => n3255, B2 => 
                           n3502, C1 => n4425, C2 => n4105, ZN => n1437);
   U2097 : INV_X1 port map( A => n1437, ZN => n4092);
   U2098 : INV_X1 port map( A => n4187, ZN => n4059);
   U2099 : NAND3_X1 port map( A1 => n4162, A2 => n4161, A3 => n4061, ZN => 
                           n4163);
   U2100 : NAND3_X1 port map( A1 => n4240, A2 => n4164, A3 => n4163, ZN => 
                           n4169);
   U2101 : NOR2_X1 port map( A1 => n4165, A2 => n4169, ZN => n4245);
   U2102 : OAI21_X1 port map( B1 => n3589, B2 => n4245, A => n4059, ZN => n301)
                           ;
   U2103 : CLKBUF_X1 port map( A => n301, Z => n4435);
   U2104 : NAND2_X1 port map( A1 => n4054, A2 => n4190, ZN => n4048);
   U2105 : NOR2_X1 port map( A1 => n4038, A2 => n4048, ZN => n4166);
   U2106 : NOR2_X1 port map( A1 => n4166, A2 => n3160, ZN => n4175);
   U2107 : AND3_X1 port map( A1 => n4175, A2 => n3596, A3 => DRAM_READY, ZN => 
                           n3888);
   U2108 : CLKBUF_X1 port map( A => n3888, Z => n4434);
   U2109 : NOR2_X1 port map( A1 => n3110, A2 => n4219, ZN => n4218);
   U2110 : NAND2_X1 port map( A1 => n4218, A2 => n3218, ZN => n4216);
   U2111 : OAI211_X1 port map( C1 => n4218, C2 => n3218, A => n3553, B => n4216
                           , ZN => n4167);
   U2112 : NAND2_X1 port map( A1 => n3123, A2 => n4167, ZN => n4386);
   U2113 : INV_X1 port map( A => n4386, ZN => n4098);
   U2114 : INV_X1 port map( A => datapath_i_alu_output_val_i_22_port, ZN => 
                           n4168);
   U2115 : OAI222_X1 port map( A1 => n4168, A2 => n4419, B1 => n3255, B2 => 
                           n3504, C1 => n4425, C2 => n4098, ZN => n1435);
   U2116 : INV_X1 port map( A => n1435, ZN => n4091);
   U2117 : INV_X1 port map( A => n4169, ZN => n4170);
   U2118 : OAI211_X1 port map( C1 => n4170, C2 => n4421, A => n4059, B => n4365
                           , ZN => enable_rf_i);
   U2119 : OAI21_X1 port map( B1 => n4038, B2 => n4048, A => n4416, ZN => 
                           write_rf_i);
   U2120 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U2121 : OAI211_X1 port map( C1 => n3265, C2 => n3225, A => n3553, B => n3264
                           , ZN => n4171);
   U2122 : NAND2_X1 port map( A1 => n3130, A2 => n4171, ZN => n4287);
   U2123 : INV_X1 port map( A => n4287, ZN => n4109);
   U2124 : INV_X1 port map( A => datapath_i_alu_output_val_i_8_port, ZN => 
                           n4172);
   U2125 : OAI222_X1 port map( A1 => n4172, A2 => n4420, B1 => n3255, B2 => 
                           n3490, C1 => n4425, C2 => n4109, ZN => n1449);
   U2126 : INV_X1 port map( A => n1449, ZN => n4110);
   U2127 : OAI211_X1 port map( C1 => n3224, C2 => n3263, A => n3553, B => n4234
                           , ZN => n4173);
   U2128 : NAND2_X1 port map( A1 => n3129, A2 => n4173, ZN => n4279);
   U2129 : INV_X1 port map( A => n4279, ZN => n4107);
   U2130 : INV_X1 port map( A => datapath_i_alu_output_val_i_10_port, ZN => 
                           n4174);
   U2131 : OAI222_X1 port map( A1 => n4174, A2 => n4420, B1 => n3255, B2 => 
                           n3492, C1 => n4425, C2 => n4107, ZN => n1447);
   U2132 : INV_X1 port map( A => n1447, ZN => n4108);
   U2133 : NOR2_X1 port map( A1 => n4175, A2 => n3266, ZN => n3889);
   U2134 : CLKBUF_X1 port map( A => n3889, Z => n4433);
   U2135 : NOR2_X1 port map( A1 => n3100, A2 => n4216, ZN => n4215);
   U2136 : NAND2_X1 port map( A1 => n4215, A2 => n3217, ZN => n4213);
   U2137 : OAI211_X1 port map( C1 => n4215, C2 => n3217, A => n3553, B => n4213
                           , ZN => n4176);
   U2138 : NAND2_X1 port map( A1 => n3122, A2 => n4176, ZN => n4258);
   U2139 : INV_X1 port map( A => n4258, ZN => n4103);
   U2140 : INV_X1 port map( A => datapath_i_alu_output_val_i_24_port, ZN => 
                           n4177);
   U2141 : OAI222_X1 port map( A1 => n4177, A2 => n4419, B1 => n3255, B2 => 
                           n3506, C1 => n4425, C2 => n4103, ZN => n1433);
   U2142 : INV_X1 port map( A => n1433, ZN => n4090);
   U2143 : NOR2_X1 port map( A1 => n3098, A2 => n4213, ZN => n4212);
   U2144 : NAND2_X1 port map( A1 => n4212, A2 => n3216, ZN => n4210);
   U2145 : OAI211_X1 port map( C1 => n4212, C2 => n3216, A => n3553, B => n4210
                           , ZN => n4178);
   U2146 : NAND2_X1 port map( A1 => n3121, A2 => n4178, ZN => n4254);
   U2147 : INV_X1 port map( A => n4254, ZN => n4104);
   U2148 : INV_X1 port map( A => datapath_i_alu_output_val_i_26_port, ZN => 
                           n4179);
   U2149 : OAI222_X1 port map( A1 => n4179, A2 => n4419, B1 => n3255, B2 => 
                           n3508, C1 => n4425, C2 => n4104, ZN => n1431);
   U2150 : INV_X1 port map( A => n1431, ZN => n4089);
   U2151 : NOR2_X1 port map( A1 => n3091, A2 => n4210, ZN => n4209);
   U2152 : NAND2_X1 port map( A1 => n4209, A2 => n3215, ZN => n4199);
   U2153 : OAI211_X1 port map( C1 => n4209, C2 => n3215, A => n3553, B => n4199
                           , ZN => n4180);
   U2154 : NAND2_X1 port map( A1 => n3120, A2 => n4180, ZN => n4252);
   U2155 : INV_X1 port map( A => n4252, ZN => n4111);
   U2156 : INV_X1 port map( A => datapath_i_alu_output_val_i_28_port, ZN => 
                           n4181);
   U2157 : OAI222_X1 port map( A1 => n4181, A2 => n4419, B1 => n3255, B2 => 
                           n3510, C1 => n4425, C2 => n4111, ZN => n1429);
   U2158 : INV_X1 port map( A => n1429, ZN => n4088);
   U2159 : NOR2_X1 port map( A1 => n3089, A2 => n4199, ZN => n4198);
   U2160 : NAND2_X1 port map( A1 => n4198, A2 => n3213, ZN => n4184);
   U2161 : OAI211_X1 port map( C1 => n4198, C2 => n3213, A => n3553, B => n4184
                           , ZN => n4182);
   U2162 : NAND2_X1 port map( A1 => n3119, A2 => n4182, ZN => n4250);
   U2163 : INV_X1 port map( A => n4250, ZN => n4096);
   U2164 : INV_X1 port map( A => datapath_i_alu_output_val_i_30_port, ZN => 
                           n4183);
   U2165 : OAI222_X1 port map( A1 => n4183, A2 => n4419, B1 => n3255, B2 => 
                           n3512, C1 => n4425, C2 => n4096, ZN => n1427);
   U2166 : INV_X1 port map( A => n1427, ZN => n4087);
   U2167 : XOR2_X1 port map( A => n3214, B => n4184, Z => n4185);
   U2168 : AOI22_X1 port map( A1 => n3553, A2 => n4185, B1 => n3114, B2 => 
                           n3243, ZN => n4395);
   U2169 : INV_X1 port map( A => n4395, ZN => n4097);
   U2170 : AOI22_X1 port map( A1 => n3257, A2 => n3116, B1 => n3557, B2 => 
                           datapath_i_alu_output_val_i_2_port, ZN => n4186);
   U2171 : OAI21_X1 port map( B1 => n3255, B2 => n3545, A => n4186, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U2172 : OR2_X1 port map( A1 => cu_i_cmd_word_6_port, A2 => n4187, ZN => 
                           cu_i_n135);
   U2173 : NOR2_X1 port map( A1 => n4047, A2 => cu_i_n135, ZN => n4189);
   U2174 : NOR2_X1 port map( A1 => n4189, A2 => n4188, ZN => n4043);
   U2175 : INV_X1 port map( A => n4043, ZN => n1802);
   U2176 : AOI221_X1 port map( B1 => n3212, B2 => n4047, C1 => cu_i_n135, C2 =>
                           n1801, A => n3118, ZN => n4337);
   U2177 : INV_X1 port map( A => n4337, ZN => n4042);
   U2178 : INV_X1 port map( A => n4053, ZN => n4243);
   U2179 : NAND2_X1 port map( A1 => n4243, A2 => n4190, ZN => n477);
   U2180 : AOI22_X1 port map( A1 => n3277, A2 => n477, B1 => n4054, B2 => n4191
                           , ZN => n4192);
   U2181 : AOI21_X1 port map( B1 => n3252, B2 => n4192, A => n1801, ZN => n3629
                           );
   U2182 : INV_X1 port map( A => datapath_i_alu_output_val_i_5_port, ZN => 
                           n4194);
   U2183 : AOI22_X1 port map( A1 => n3257, A2 => n3262, B1 => n3457, B2 => 
                           n3455, ZN => n4193);
   U2184 : OAI21_X1 port map( B1 => n4420, B2 => n4194, A => n4193, ZN => n4117
                           );
   U2185 : AOI211_X1 port map( C1 => n3264, C2 => n3094, A => n3263, B => n3114
                           , ZN => n4195);
   U2186 : NOR2_X1 port map( A1 => n3146, A2 => n4195, ZN => n4118);
   U2187 : AOI22_X1 port map( A1 => n3117, A2 => 
                           datapath_i_alu_output_val_i_9_port, B1 => n3457, B2 
                           => n3453, ZN => n4196);
   U2188 : OAI21_X1 port map( B1 => n4118, B2 => n4425, A => n4196, ZN => n4115
                           );
   U2189 : NOR2_X1 port map( A1 => n3148, A2 => n3150, ZN => n4130);
   U2190 : AOI22_X1 port map( A1 => n3117, A2 => 
                           datapath_i_alu_output_val_i_7_port, B1 => n3457, B2 
                           => n3454, ZN => n4197);
   U2191 : OAI21_X1 port map( B1 => n4130, B2 => n4425, A => n4197, ZN => n4116
                           );
   U2192 : AOI211_X1 port map( C1 => n3088, C2 => n4199, A => n3114, B => n4198
                           , ZN => n4200);
   U2193 : NOR2_X1 port map( A1 => n3136, A2 => n4200, ZN => n4119);
   U2194 : AOI22_X1 port map( A1 => n3278, A2 => cu_i_cmd_alu_op_type_1_port, 
                           B1 => n3456, B2 => n3279, ZN => n4206);
   U2195 : AOI21_X1 port map( B1 => n4204, B2 => n4206, A => n4203, ZN => n4201
                           );
   U2196 : NOR2_X1 port map( A1 => n4207, A2 => n4201, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U2197 : AOI21_X1 port map( B1 => n4204, B2 => n4207, A => n4203, ZN => n4202
                           );
   U2198 : NOR2_X1 port map( A1 => n4206, A2 => n4202, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U2199 : INV_X1 port map( A => n4203, ZN => n4205);
   U2200 : OAI211_X1 port map( C1 => n4207, C2 => n4206, A => n4205, B => n4204
                           , ZN => n4208);
   U2201 : INV_X1 port map( A => n4208, ZN => n4033);
   U2202 : AOI211_X1 port map( C1 => n3090, C2 => n4210, A => n3114, B => n4209
                           , ZN => n4211);
   U2203 : NOR2_X1 port map( A1 => n3137, A2 => n4211, ZN => n4120);
   U2204 : AOI211_X1 port map( C1 => n3097, C2 => n4213, A => n3114, B => n4212
                           , ZN => n4214);
   U2205 : NOR2_X1 port map( A1 => n3138, A2 => n4214, ZN => n4121);
   U2206 : AOI211_X1 port map( C1 => n3099, C2 => n4216, A => n3114, B => n4215
                           , ZN => n4217);
   U2207 : NOR2_X1 port map( A1 => n3139, A2 => n4217, ZN => n4122);
   U2208 : AOI211_X1 port map( C1 => n3109, C2 => n4219, A => n3114, B => n4218
                           , ZN => n4220);
   U2209 : NOR2_X1 port map( A1 => n3140, A2 => n4220, ZN => n4123);
   U2210 : AOI211_X1 port map( C1 => n3107, C2 => n4222, A => n3114, B => n4221
                           , ZN => n4223);
   U2211 : NOR2_X1 port map( A1 => n3141, A2 => n4223, ZN => n4124);
   U2212 : AOI211_X1 port map( C1 => n3105, C2 => n4225, A => n3114, B => n4224
                           , ZN => n4226);
   U2213 : NOR2_X1 port map( A1 => n3142, A2 => n4226, ZN => n4125);
   U2214 : AOI211_X1 port map( C1 => n3101, C2 => n4228, A => n3114, B => n4227
                           , ZN => n4229);
   U2215 : NOR2_X1 port map( A1 => n3143, A2 => n4229, ZN => n4126);
   U2216 : AOI211_X1 port map( C1 => n3103, C2 => n4231, A => n3114, B => n4230
                           , ZN => n4232);
   U2217 : NOR2_X1 port map( A1 => n3144, A2 => n4232, ZN => n4127);
   U2218 : AOI211_X1 port map( C1 => n3092, C2 => n4234, A => n3114, B => n4233
                           , ZN => n4235);
   U2219 : NOR2_X1 port map( A1 => n3145, A2 => n4235, ZN => n4128);
   U2220 : MUX2_X1 port map( A => n3167, B => n3303, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U2221 : CLKBUF_X1 port map( A => n4426, Z => n4430);
   U2222 : AOI22_X1 port map( A1 => n3257, A2 => n3260, B1 => n3117, B2 => 
                           datapath_i_alu_output_val_i_4_port, ZN => n4236);
   U2223 : OAI21_X1 port map( B1 => n3255, B2 => n3486, A => n4236, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U2224 : AOI22_X1 port map( A1 => n3257, A2 => n3244, B1 => n3557, B2 => 
                           datapath_i_alu_output_val_i_3_port, ZN => n4237);
   U2225 : OAI21_X1 port map( B1 => n3255, B2 => n3547, A => n4237, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U2226 : INV_X1 port map( A => n4117, ZN => n4302);
   U2227 : NAND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_2_port,
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, ZN
                           => n4400);
   U2228 : INV_X1 port map( A => n4400, ZN => n4294);
   U2229 : NAND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port,
                           A2 => n4294, ZN => n4285);
   U2230 : NOR2_X1 port map( A1 => n4302, A2 => n4285, ZN => n4298);
   U2231 : AOI211_X1 port map( C1 => n4302, C2 => n4285, A => n3115, B => n4298
                           , ZN => n4238);
   U2232 : OR2_X1 port map( A1 => n3147, A2 => n4238, ZN => 
                           datapath_i_new_pc_value_decode_5_port);
   U2233 : NOR4_X1 port map( A1 => n1402, A2 => n1404, A3 => n1401, A4 => n1405
                           , ZN => n4239);
   U2234 : NAND2_X1 port map( A1 => n4364, A2 => n4239, ZN => n4244);
   U2235 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_17_port, A2 => 
                           curr_instruction_to_cu_i_19_port, A3 => 
                           curr_instruction_to_cu_i_16_port, A4 => 
                           curr_instruction_to_cu_i_20_port, ZN => n4241);
   U2236 : AOI21_X1 port map( B1 => n4366, B2 => n4241, A => n4240, ZN => n4242
                           );
   U2237 : AOI221_X1 port map( B1 => n4245, B2 => n4053, C1 => n4244, C2 => 
                           n4243, A => n4242, ZN => n4246);
   U2238 : OAI21_X1 port map( B1 => n3589, B2 => n4246, A => n4361, ZN => n4247
                           );
   U2239 : AOI211_X1 port map( C1 => n3544, C2 => n3245, A => cu_i_n135, B => 
                           n4247, ZN => n4052);
   U2240 : OR2_X1 port map( A1 => n3246, A2 => n4052, ZN => n3635);
   U2241 : INV_X1 port map( A => n4422, ZN => n4431);
   U2242 : OR2_X1 port map( A1 => n3577, A2 => n3458, ZN => cu_i_N278);
   U2243 : INV_X1 port map( A => n3655, ZN => IRAM_ADDRESS_8_port);
   U2244 : INV_X1 port map( A => n3667, ZN => IRAM_ADDRESS_10_port);
   U2245 : INV_X1 port map( A => n3666, ZN => IRAM_ADDRESS_12_port);
   U2246 : INV_X1 port map( A => n3668, ZN => IRAM_ADDRESS_14_port);
   U2247 : INV_X1 port map( A => n3665, ZN => IRAM_ADDRESS_16_port);
   U2248 : INV_X1 port map( A => n3661, ZN => IRAM_ADDRESS_18_port);
   U2249 : INV_X1 port map( A => n3656, ZN => IRAM_ADDRESS_20_port);
   U2250 : INV_X1 port map( A => n3657, ZN => IRAM_ADDRESS_22_port);
   U2251 : INV_X1 port map( A => n3660, ZN => IRAM_ADDRESS_24_port);
   U2252 : INV_X1 port map( A => n3663, ZN => IRAM_ADDRESS_26_port);
   U2253 : INV_X1 port map( A => n3662, ZN => IRAM_ADDRESS_28_port);
   U2254 : INV_X1 port map( A => n3659, ZN => IRAM_ADDRESS_30_port);
   U2255 : CLKBUF_X1 port map( A => n3241, Z => n4389);
   U2256 : INV_X1 port map( A => n4119, ZN => n4248);
   U2257 : AOI22_X1 port map( A1 => n4389, A2 => n4248, B1 => n3558, B2 => 
                           n3436, ZN => n4249);
   U2258 : OAI21_X1 port map( B1 => n3559, B2 => n3484, A => n4249, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U2259 : AOI22_X1 port map( A1 => n3241, A2 => n4250, B1 => n3156, B2 => 
                           n3438, ZN => n4251);
   U2260 : OAI21_X1 port map( B1 => n3512, B2 => n3559, A => n4251, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U2261 : AOI22_X1 port map( A1 => n4389, A2 => n4252, B1 => n3156, B2 => 
                           n3434, ZN => n4253);
   U2262 : OAI21_X1 port map( B1 => n3559, B2 => n3510, A => n4253, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U2263 : AOI22_X1 port map( A1 => n3241, A2 => n4254, B1 => n3156, B2 => 
                           n3430, ZN => n4255);
   U2264 : OAI21_X1 port map( B1 => n3559, B2 => n3508, A => n4255, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U2265 : INV_X1 port map( A => n4121, ZN => n4256);
   U2266 : AOI22_X1 port map( A1 => n3241, A2 => n4256, B1 => n3558, B2 => 
                           n3428, ZN => n4257);
   U2267 : OAI21_X1 port map( B1 => n3559, B2 => n3480, A => n4257, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U2268 : AOI22_X1 port map( A1 => n3241, A2 => n4258, B1 => n3558, B2 => 
                           n3426, ZN => n4259);
   U2269 : OAI21_X1 port map( B1 => n3261, B2 => n3506, A => n4259, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U2270 : INV_X1 port map( A => n4124, ZN => n4260);
   U2271 : AOI22_X1 port map( A1 => n3241, A2 => n4260, B1 => n3558, B2 => 
                           n3416, ZN => n4261);
   U2272 : AOI22_X1 port map( A1 => n3241, A2 => n4262, B1 => n3156, B2 => 
                           n3414, ZN => n4263);
   U2273 : OAI21_X1 port map( B1 => n3261, B2 => n3500, A => n4263, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U2274 : AOI22_X1 port map( A1 => n3241, A2 => n3259, B1 => n3558, B2 => 
                           n3390, ZN => n4264);
   U2275 : OAI21_X1 port map( B1 => n3261, B2 => n3488, A => n4264, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);
   U2276 : INV_X1 port map( A => n4130, ZN => n4265);
   U2277 : AOI22_X1 port map( A1 => n3241, A2 => n4265, B1 => n3156, B2 => 
                           n3392, ZN => n4266);
   U2278 : OAI21_X1 port map( B1 => n3559, B2 => n3459, A => n4266, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U2279 : INV_X1 port map( A => n4118, ZN => n4267);
   U2280 : AOI22_X1 port map( A1 => n4389, A2 => n4267, B1 => n3156, B2 => 
                           n3396, ZN => n4268);
   U2281 : OAI21_X1 port map( B1 => n3261, B2 => n3463, A => n4268, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U2282 : INV_X1 port map( A => n4126, ZN => n4269);
   U2283 : AOI22_X1 port map( A1 => n3241, A2 => n4269, B1 => n3156, B2 => 
                           n3408, ZN => n4270);
   U2284 : AOI22_X1 port map( A1 => n3241, A2 => n4271, B1 => n3558, B2 => 
                           n3410, ZN => n4272);
   U2285 : OAI21_X1 port map( B1 => n3261, B2 => n3498, A => n4272, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U2286 : AOI22_X1 port map( A1 => n3241, A2 => n4273, B1 => n3558, B2 => 
                           n3406, ZN => n4274);
   U2287 : AOI22_X1 port map( A1 => n4389, A2 => n4275, B1 => n3558, B2 => 
                           n3402, ZN => n4276);
   U2288 : OAI21_X1 port map( B1 => n3261, B2 => n3494, A => n4276, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U2289 : INV_X1 port map( A => n4128, ZN => n4277);
   U2290 : AOI22_X1 port map( A1 => n3241, A2 => n4277, B1 => n3156, B2 => 
                           n3400, ZN => n4278);
   U2291 : AOI22_X1 port map( A1 => n3241, A2 => n4279, B1 => n3558, B2 => 
                           n3398, ZN => n4280);
   U2292 : MUX2_X1 port map( A => n3170, B => n3294, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U2293 : MUX2_X1 port map( A => n3169, B => n3297, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U2294 : NAND2_X1 port map( A1 => n3281, A2 => n3284, ZN => n4324);
   U2295 : INV_X1 port map( A => n4324, ZN => n4325);
   U2296 : NAND2_X1 port map( A1 => n4325, A2 => n4417, ZN => n4281);
   U2297 : NOR2_X1 port map( A1 => n3643, A2 => n4281, ZN => n4283);
   U2298 : OAI22_X1 port map( A1 => n4417, A2 => n3473, B1 => n4325, B2 => 
                           n3643, ZN => n4282);
   U2299 : MUX2_X1 port map( A => n4283, B => n4282, S => n3282, Z => cu_i_N277
                           );
   datapath_i_execute_stage_dp_n9 <= '0';
   U2301 : MUX2_X1 port map( A => n3177, B => n3288, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U2302 : AOI22_X1 port map( A1 => n3257, A2 => n3259, B1 => n3117, B2 => 
                           datapath_i_alu_output_val_i_6_port, ZN => n4284);
   U2303 : OAI21_X1 port map( B1 => n3255, B2 => n3488, A => n4284, ZN => n1453
                           );
   U2304 : INV_X1 port map( A => n4116, ZN => n4303);
   U2305 : INV_X1 port map( A => n4285, ZN => n4296);
   U2306 : NAND3_X1 port map( A1 => n4296, A2 => n1453, A3 => n4117, ZN => 
                           n4297);
   U2307 : NOR2_X1 port map( A1 => n4303, A2 => n4297, ZN => n2359);
   U2308 : NAND2_X1 port map( A1 => n2359, A2 => n1449, ZN => n2358);
   U2309 : INV_X1 port map( A => n4115, ZN => n4286);
   U2310 : NOR2_X1 port map( A1 => n4286, A2 => n2358, ZN => n2363);
   U2311 : AOI211_X1 port map( C1 => n4303, C2 => n4297, A => n3115, B => n2359
                           , ZN => n2350);
   U2312 : AOI22_X1 port map( A1 => n3241, A2 => n4287, B1 => n3156, B2 => 
                           n3394, ZN => n4288);
   U2313 : OAI21_X1 port map( B1 => n3261, B2 => n3490, A => n4288, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U2314 : NAND2_X1 port map( A1 => n4043, A2 => n3586, ZN => n1507);
   U2315 : AOI22_X1 port map( A1 => n3257, A2 => n3162, B1 => n3557, B2 => 
                           datapath_i_alu_output_val_i_1_port, ZN => n4289);
   U2316 : OAI21_X1 port map( B1 => n3255, B2 => n3541, A => n4289, ZN => n3627
                           );
   U2317 : MUX2_X1 port map( A => n3627, B => IRAM_ADDRESS_1_port, S => n3115, 
                           Z => n1385);
   U2318 : NOR2_X1 port map( A1 => n3586, A2 => n1802, ZN => n1727);
   U2319 : AOI22_X1 port map( A1 => n1385, A2 => n1727, B1 => n3384, B2 => 
                           n1802, ZN => n4290);
   U2320 : OAI21_X1 port map( B1 => n3542, B2 => n1507, A => n4290, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U2321 : AOI22_X1 port map( A1 => n3241, A2 => n3262, B1 => n3156, B2 => 
                           n3388, ZN => n4291);
   U2322 : OAI21_X1 port map( B1 => n3559, B2 => n3461, A => n4291, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U2323 : AOI22_X1 port map( A1 => n4389, A2 => n4292, B1 => n3156, B2 => 
                           n3418, ZN => n4293);
   U2324 : OAI21_X1 port map( B1 => n3559, B2 => n3502, A => n4293, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U2325 : MUX2_X1 port map( A => n3171, B => n3291, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U2326 : OAI21_X1 port map( B1 => n4294, B2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n3554, ZN => n4295);
   U2327 : OAI21_X1 port map( B1 => n4296, B2 => n4295, A => n3132, ZN => 
                           datapath_i_new_pc_value_decode_4_port);
   U2328 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_4_port, B1 => n3387, 
                           B2 => n1802, ZN => n2398);
   U2329 : OAI21_X1 port map( B1 => n3261, B2 => n3486, A => n3149, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U2330 : OAI211_X1 port map( C1 => n4298, C2 => n1453, A => n3554, B => n4297
                           , ZN => n4299);
   U2331 : NAND2_X1 port map( A1 => n3131, A2 => n4299, ZN => 
                           datapath_i_new_pc_value_decode_6_port);
   U2332 : INV_X1 port map( A => n4040, ZN => n4300);
   U2333 : NOR2_X1 port map( A1 => n4378, A2 => n4300, ZN => n1758);
   U2334 : NAND2_X1 port map( A1 => n3587, A2 => n4040, ZN => n1505);
   U2335 : NAND2_X1 port map( A1 => n4044, A2 => n4301, ZN => n1497);
   U2336 : NAND2_X1 port map( A1 => n3246, A2 => n4052, ZN => n2416);
   U2337 : AOI211_X1 port map( C1 => n3251, C2 => n3096, A => n3554, B => n3250
                           , ZN => n1346);
   U2338 : INV_X1 port map( A => n3629, ZN => n4397);
   U2339 : NOR2_X1 port map( A1 => n4400, A2 => n4397, ZN => n4336);
   U2340 : NAND2_X1 port map( A1 => n4336, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n4335);
   U2341 : NOR2_X1 port map( A1 => n4302, A2 => n4335, ZN => n4338);
   U2342 : AOI211_X1 port map( C1 => n4302, C2 => n4335, A => n4338, B => n4042
                           , ZN => n1345);
   U2343 : NAND2_X1 port map( A1 => n4338, A2 => n1453, ZN => n2483);
   U2344 : NOR2_X1 port map( A1 => n4303, A2 => n2483, ZN => n2486);
   U2345 : NAND2_X1 port map( A1 => n2486, A2 => n1449, ZN => n2485);
   U2346 : NOR2_X1 port map( A1 => n3249, A2 => n3095, ZN => n4340);
   U2347 : AOI211_X1 port map( C1 => n3095, C2 => n3249, A => n4340, B => n3554
                           , ZN => n1344);
   U2348 : NAND2_X1 port map( A1 => n3224, A2 => n4340, ZN => n4339);
   U2349 : NOR2_X1 port map( A1 => n3093, A2 => n4339, ZN => n4342);
   U2350 : AOI211_X1 port map( C1 => n3093, C2 => n4339, A => n4342, B => n3554
                           , ZN => n1343);
   U2351 : NAND2_X1 port map( A1 => n3223, A2 => n4342, ZN => n4341);
   U2352 : NOR2_X1 port map( A1 => n3104, A2 => n4341, ZN => n4344);
   U2353 : AOI211_X1 port map( C1 => n3104, C2 => n4341, A => n4344, B => n3554
                           , ZN => n1342);
   U2354 : NAND2_X1 port map( A1 => n3222, A2 => n4344, ZN => n4343);
   U2355 : NOR2_X1 port map( A1 => n3102, A2 => n4343, ZN => n4346);
   U2356 : AOI211_X1 port map( C1 => n3102, C2 => n4343, A => n4346, B => n3554
                           , ZN => n1341);
   U2357 : NAND2_X1 port map( A1 => n3221, A2 => n4346, ZN => n4345);
   U2358 : NOR2_X1 port map( A1 => n3106, A2 => n4345, ZN => n4348);
   U2359 : AOI211_X1 port map( C1 => n3106, C2 => n4345, A => n4348, B => n3554
                           , ZN => n1340);
   U2360 : NAND2_X1 port map( A1 => n3220, A2 => n4348, ZN => n4347);
   U2361 : NOR2_X1 port map( A1 => n3108, A2 => n4347, ZN => n4350);
   U2362 : AOI211_X1 port map( C1 => n3108, C2 => n4347, A => n4350, B => n3554
                           , ZN => n1339);
   U2363 : NAND2_X1 port map( A1 => n3219, A2 => n4350, ZN => n4349);
   U2364 : NOR2_X1 port map( A1 => n3110, A2 => n4349, ZN => n4352);
   U2365 : AOI211_X1 port map( C1 => n3110, C2 => n4349, A => n4352, B => n3554
                           , ZN => n1338);
   U2366 : NAND2_X1 port map( A1 => n3218, A2 => n4352, ZN => n4351);
   U2367 : NOR2_X1 port map( A1 => n3100, A2 => n4351, ZN => n4354);
   U2368 : AOI211_X1 port map( C1 => n3100, C2 => n4351, A => n4354, B => n3554
                           , ZN => n1337);
   U2369 : NAND2_X1 port map( A1 => n3217, A2 => n4354, ZN => n4353);
   U2370 : NOR2_X1 port map( A1 => n3098, A2 => n4353, ZN => n4356);
   U2371 : AOI211_X1 port map( C1 => n3098, C2 => n4353, A => n4356, B => n3554
                           , ZN => n1336);
   U2372 : NAND2_X1 port map( A1 => n3216, A2 => n4356, ZN => n4355);
   U2373 : NOR2_X1 port map( A1 => n3091, A2 => n4355, ZN => n4358);
   U2374 : AOI211_X1 port map( C1 => n3091, C2 => n4355, A => n4358, B => n3554
                           , ZN => n1335);
   U2375 : NAND2_X1 port map( A1 => n3215, A2 => n4358, ZN => n4357);
   U2376 : NOR2_X1 port map( A1 => n3089, A2 => n4357, ZN => n4359);
   U2377 : AOI211_X1 port map( C1 => n3089, C2 => n4357, A => n4359, B => n3554
                           , ZN => n1334);
   U2378 : AOI22_X1 port map( A1 => n1801, A2 => n4435, B1 => n3577, B2 => 
                           n4047, ZN => n1728);
   U2379 : INV_X1 port map( A => datapath_i_alu_output_val_i_31_port, ZN => 
                           n4304);
   U2380 : OAI222_X1 port map( A1 => n4304, A2 => n4420, B1 => n3255, B2 => 
                           n3549, C1 => n4425, C2 => n4097, ZN => n1916);
   U2381 : NOR4_X1 port map( A1 => n3236, A2 => n3238, A3 => n3588, A4 => n3151
                           , ZN => n4319);
   U2382 : NOR2_X1 port map( A1 => n3153, A2 => n3237, ZN => n4316);
   U2383 : NAND2_X1 port map( A1 => n3247, A2 => n4428, ZN => n4311);
   U2384 : INV_X1 port map( A => n4319, ZN => n4306);
   U2385 : NOR3_X1 port map( A1 => n3238, A2 => n3588, A3 => n3151, ZN => n4305
                           );
   U2386 : NAND3_X1 port map( A1 => n3236, A2 => n4305, A3 => n3152, ZN => 
                           n4323);
   U2387 : OAI211_X1 port map( C1 => n3152, C2 => n4311, A => n4306, B => n4323
                           , ZN => n4307);
   U2388 : AOI22_X1 port map( A1 => n4319, A2 => n3248, B1 => n4316, B2 => 
                           n4307, ZN => n4310);
   U2389 : NAND3_X1 port map( A1 => n3271, A2 => n3275, A3 => n4427, ZN => 
                           n4309);
   U2390 : NAND2_X1 port map( A1 => n3532, A2 => n3155, ZN => n4308);
   U2391 : NAND4_X1 port map( A1 => n3239, A2 => n4310, A3 => n4309, A4 => 
                           n4308, ZN => cu_i_N264);
   U2392 : NOR2_X1 port map( A1 => n4311, A2 => n3536, ZN => n4312);
   U2393 : AOI21_X1 port map( B1 => n4312, B2 => n4316, A => n3155, ZN => n4321
                           );
   U2394 : NOR3_X1 port map( A1 => n3537, A2 => n3664, A3 => n4323, ZN => n4315
                           );
   U2395 : NAND3_X1 port map( A1 => n3158, A2 => n3639, A3 => n3271, ZN => 
                           n4313);
   U2396 : NAND2_X1 port map( A1 => n4313, A2 => n3253, ZN => n4314);
   U2397 : AOI211_X1 port map( C1 => n3275, C2 => n3638, A => n4315, B => n4314
                           , ZN => n4318);
   U2398 : NAND3_X1 port map( A1 => n4319, A2 => n4316, A3 => n3152, ZN => 
                           n4317);
   U2399 : NAND3_X1 port map( A1 => n4321, A2 => n4318, A3 => n4317, ZN => 
                           cu_i_N265);
   U2400 : OAI221_X1 port map( B1 => n3248, B2 => n3152, C1 => n3248, C2 => 
                           n3237, A => n4319, ZN => n4322);
   U2401 : OAI221_X1 port map( B1 => n3639, B2 => n3532, C1 => n3639, C2 => 
                           n3159, A => n3638, ZN => n4320);
   U2402 : OAI211_X1 port map( C1 => n3153, C2 => n4322, A => n4321, B => n4320
                           , ZN => cu_i_N266);
   U2403 : OAI221_X1 port map( B1 => n4323, B2 => n3153, C1 => n4323, C2 => 
                           n3664, A => n3154, ZN => cu_i_N267);
   U2404 : NAND2_X1 port map( A1 => n3278, A2 => n3473, ZN => cu_i_N274);
   U2405 : AOI211_X1 port map( C1 => n4418, C2 => n4429, A => n3473, B => n4325
                           , ZN => cu_i_N275);
   U2406 : NOR2_X1 port map( A1 => n3281, A2 => n3473, ZN => cu_i_N273);
   U2407 : AOI221_X1 port map( B1 => n4325, B2 => n4417, C1 => n4324, C2 => 
                           n3670, A => n3643, ZN => cu_i_N276);
   U2408 : AOI211_X1 port map( C1 => n3278, C2 => n3235, A => n3473, B => n3268
                           , ZN => cu_i_N279);
   U2409 : NOR2_X1 port map( A1 => n4326, A2 => n1390, ZN => n1477);
   U2410 : NOR2_X1 port map( A1 => n1393, A2 => n1394, ZN => n492);
   U2411 : NAND4_X1 port map( A1 => n4414, A2 => n4327, A3 => n3277, A4 => 
                           n4415, ZN => n4331);
   U2412 : NAND4_X1 port map( A1 => n4328, A2 => n1477, A3 => n492, A4 => n4049
                           , ZN => n4330);
   U2413 : OAI22_X1 port map( A1 => n4332, A2 => n4331, B1 => n4330, B2 => 
                           n4329, ZN => cu_i_cmd_word_8_port);
   U2414 : MUX2_X1 port map( A => n3134, B => cu_i_cmd_word_8_port, S => n1801,
                           Z => alu_cin_i);
   U2415 : MUX2_X1 port map( A => n3276, B => n3211, S => n1801, Z => n1425);
   U2416 : MUX2_X1 port map( A => n3590, B => n3210, S => n1801, Z => n1424);
   U2417 : NOR2_X1 port map( A1 => n4052, A2 => n4423, ZN => n1475);
   U2418 : MUX2_X1 port map( A => n3111, B => n3209, S => n1801, Z => n1423);
   U2419 : MUX2_X1 port map( A => n3269, B => n3208, S => n1801, Z => n1422);
   U2420 : MUX2_X1 port map( A => IRAM_DATA(25), B => n3207, S => n3555, Z => 
                           n1415);
   U2421 : MUX2_X1 port map( A => IRAM_DATA(24), B => n3206, S => n3555, Z => 
                           n1414);
   U2422 : MUX2_X1 port map( A => IRAM_DATA(22), B => n3204, S => n3278, Z => 
                           n1412);
   U2423 : MUX2_X1 port map( A => IRAM_DATA(21), B => n3203, S => n3278, Z => 
                           n1411);
   U2424 : MUX2_X1 port map( A => IRAM_DATA(10), B => n3202, S => n3555, Z => 
                           n1400);
   U2425 : MUX2_X1 port map( A => IRAM_DATA(9), B => n3201, S => n3555, Z => 
                           n1399);
   U2426 : MUX2_X1 port map( A => IRAM_DATA(8), B => n3200, S => n3555, Z => 
                           n1398);
   U2427 : MUX2_X1 port map( A => IRAM_DATA(7), B => n3199, S => n3555, Z => 
                           n1397);
   U2428 : MUX2_X1 port map( A => IRAM_DATA(6), B => n3198, S => n3555, Z => 
                           n1396);
   U2429 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_2_port, ZN
                           => n4398);
   U2430 : NOR2_X1 port map( A1 => n4398, A2 => n4397, ZN => n4334);
   U2431 : INV_X1 port map( A => n4336, ZN => n4333);
   U2432 : OAI211_X1 port map( C1 => n4334, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, A => 
                           n4337, B => n4333, ZN => n2478);
   U2433 : OAI211_X1 port map( C1 => n4336, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n4337, B => n4335, ZN => n1325);
   U2434 : OAI211_X1 port map( C1 => n4338, C2 => n1453, A => n4337, B => n2483
                           , ZN => n1324);
   U2435 : OAI211_X1 port map( C1 => n3250, C2 => IRAM_ADDRESS_8_port, A => 
                           n3249, B => n3115, ZN => n1323);
   U2436 : OAI211_X1 port map( C1 => n4340, C2 => IRAM_ADDRESS_10_port, A => 
                           n3115, B => n4339, ZN => n1322);
   U2437 : OAI211_X1 port map( C1 => n4342, C2 => IRAM_ADDRESS_12_port, A => 
                           n3115, B => n4341, ZN => n1321);
   U2438 : OAI211_X1 port map( C1 => n4344, C2 => IRAM_ADDRESS_14_port, A => 
                           n3115, B => n4343, ZN => n1320);
   U2439 : OAI211_X1 port map( C1 => n4346, C2 => IRAM_ADDRESS_16_port, A => 
                           n3115, B => n4345, ZN => n1319);
   U2440 : OAI211_X1 port map( C1 => n4348, C2 => IRAM_ADDRESS_18_port, A => 
                           n3115, B => n4347, ZN => n1318);
   U2441 : OAI211_X1 port map( C1 => n4350, C2 => IRAM_ADDRESS_20_port, A => 
                           n3115, B => n4349, ZN => n1317);
   U2442 : OAI211_X1 port map( C1 => n4352, C2 => IRAM_ADDRESS_22_port, A => 
                           n3115, B => n4351, ZN => n1316);
   U2443 : OAI211_X1 port map( C1 => n4354, C2 => IRAM_ADDRESS_24_port, A => 
                           n3115, B => n4353, ZN => n1315);
   U2444 : OAI211_X1 port map( C1 => n4356, C2 => IRAM_ADDRESS_26_port, A => 
                           n3115, B => n4355, ZN => n1314);
   U2445 : OAI211_X1 port map( C1 => n4358, C2 => IRAM_ADDRESS_28_port, A => 
                           n3115, B => n4357, ZN => n1313);
   U2446 : NAND2_X1 port map( A1 => n3213, A2 => n4359, ZN => n4360);
   U2447 : OAI211_X1 port map( C1 => n4359, C2 => IRAM_ADDRESS_30_port, A => 
                           n3115, B => n4360, ZN => n1312);
   U2448 : XOR2_X1 port map( A => n4132, B => n4360, Z => n1460);
   U2449 : AND2_X1 port map( A1 => n3577, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U2450 : OAI21_X1 port map( B1 => n4362, B2 => n4361, A => n4365, ZN => 
                           read_rf_p2_i);
   U2451 : OAI221_X1 port map( B1 => n4367, B2 => n4366, C1 => n4365, C2 => 
                           n4364, A => n4363, ZN => n1302);
   U2452 : OAI21_X1 port map( B1 => n3540, B2 => n3596, A => n3890, ZN => 
                           datapath_i_decode_stage_dp_n44);
   U2453 : OAI21_X1 port map( B1 => n3542, B2 => n3596, A => n3887, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U2454 : OAI21_X1 port map( B1 => n3546, B2 => n3596, A => n3886, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U2455 : OAI21_X1 port map( B1 => n3548, B2 => n3596, A => n3885, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U2456 : OAI21_X1 port map( B1 => n3596, B2 => n3487, A => n3884, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U2457 : OAI21_X1 port map( B1 => n3596, B2 => n3462, A => n3883, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U2458 : OAI21_X1 port map( B1 => n3596, B2 => n3489, A => n3882, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U2459 : OAI21_X1 port map( B1 => n3596, B2 => n3460, A => n3881, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U2460 : OAI21_X1 port map( B1 => n3596, B2 => n3491, A => n3880, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U2461 : OAI21_X1 port map( B1 => n3596, B2 => n3464, A => n3879, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U2462 : OAI21_X1 port map( B1 => n3596, B2 => n3493, A => n3878, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U2463 : OAI21_X1 port map( B1 => n3596, B2 => n3466, A => n3877, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U2464 : OAI21_X1 port map( B1 => n3596, B2 => n3495, A => n3876, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U2465 : OAI21_X1 port map( B1 => n3596, B2 => n3468, A => n3875, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U2466 : OAI21_X1 port map( B1 => n3596, B2 => n3497, A => n3874, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U2467 : OAI21_X1 port map( B1 => n3596, B2 => n3470, A => n3873, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U2468 : OAI21_X1 port map( B1 => n3596, B2 => n3499, A => n3872, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U2469 : OAI21_X1 port map( B1 => n3596, B2 => n3472, A => n3871, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U2470 : OAI21_X1 port map( B1 => n3596, B2 => n3501, A => n3870, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U2471 : OAI21_X1 port map( B1 => n3596, B2 => n3475, A => n3869, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U2472 : OAI21_X1 port map( B1 => n3596, B2 => n3503, A => n3868, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U2473 : OAI21_X1 port map( B1 => n3596, B2 => n3477, A => n3867, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U2474 : OAI21_X1 port map( B1 => n3596, B2 => n3505, A => n3866, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U2475 : OAI21_X1 port map( B1 => n3596, B2 => n3479, A => n3865, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U2476 : OAI21_X1 port map( B1 => n3596, B2 => n3507, A => n3864, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U2477 : OAI21_X1 port map( B1 => n3596, B2 => n3481, A => n3863, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U2478 : OAI21_X1 port map( B1 => n3596, B2 => n3509, A => n3862, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U2479 : OAI21_X1 port map( B1 => n3596, B2 => n3483, A => n3861, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U2480 : OAI21_X1 port map( B1 => n3596, B2 => n3511, A => n3860, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U2481 : OAI21_X1 port map( B1 => n3596, B2 => n3485, A => n3859, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U2482 : OAI21_X1 port map( B1 => n3596, B2 => n3513, A => n3858, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U2483 : OAI21_X1 port map( B1 => n3596, B2 => n3550, A => n3857, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U2484 : NOR4_X1 port map( A1 => n1641, A2 => n1643, A3 => n1645, A4 => n1647
                           , ZN => n4371);
   U2485 : NOR4_X1 port map( A1 => n1649, A2 => n1651, A3 => n1653, A4 => n1655
                           , ZN => n4370);
   U2486 : NOR4_X1 port map( A1 => n1625, A2 => n1627, A3 => n1629, A4 => n1631
                           , ZN => n4369);
   U2487 : NOR4_X1 port map( A1 => n1633, A2 => n1635, A3 => n1637, A4 => n1639
                           , ZN => n4368);
   U2488 : NAND4_X1 port map( A1 => n4371, A2 => n4370, A3 => n4369, A4 => 
                           n4368, ZN => n4377);
   U2489 : NOR4_X1 port map( A1 => n1663, A2 => n1617, A3 => n1619, A4 => n1621
                           , ZN => n4375);
   U2490 : NOR4_X1 port map( A1 => n1613, A2 => n1614, A3 => n1615, A4 => n1661
                           , ZN => n4374);
   U2491 : NOR4_X1 port map( A1 => n1667, A2 => n1669, A3 => n1657, A4 => n1659
                           , ZN => n4373);
   U2492 : NOR4_X1 port map( A1 => n1623, A2 => n1671, A3 => n1673, A4 => n1665
                           , ZN => n4372);
   U2493 : NAND4_X1 port map( A1 => n4375, A2 => n4374, A3 => n4373, A4 => 
                           n4372, ZN => n4376);
   U2494 : NOR2_X1 port map( A1 => n4377, A2 => n4376, ZN => n2530);
   U2495 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, S 
                           => n4378, Z => n1383);
   U2496 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, S 
                           => n4378, Z => n1382);
   U2497 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, S 
                           => n4378, Z => n1381);
   U2498 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, S 
                           => n4378, Z => n1380);
   U2499 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, S 
                           => n3587, Z => n1379);
   U2500 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, S 
                           => n3587, Z => n1378);
   U2501 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, S 
                           => n3587, Z => n1377);
   U2502 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, S 
                           => n3587, Z => n1376);
   U2503 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, S 
                           => n3587, Z => n1375);
   U2504 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, S 
                           => n3587, Z => n1374);
   U2505 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, S 
                           => n3587, Z => n1373);
   U2506 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, S 
                           => n3587, Z => n1372);
   U2507 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, S 
                           => n3587, Z => n1371);
   U2508 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, S 
                           => n3587, Z => n1370);
   U2509 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, S 
                           => n4378, Z => n1369);
   U2510 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, S 
                           => n4378, Z => n1368);
   U2511 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, S 
                           => n4378, Z => n1367);
   U2512 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, S 
                           => n4378, Z => n1366);
   U2513 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, S 
                           => n4378, Z => n1365);
   U2514 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, S 
                           => n4378, Z => n1364);
   U2515 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, S 
                           => n3587, Z => n1363);
   U2516 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, S 
                           => n3587, Z => n1362);
   U2517 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, S 
                           => n3587, Z => n1361);
   U2518 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, S 
                           => n3587, Z => n1360);
   U2519 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, S 
                           => n3587, Z => n1359);
   U2520 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, S 
                           => n3587, Z => n1358);
   U2521 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, S 
                           => n3587, Z => n1357);
   U2522 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, S 
                           => n3587, Z => n1356);
   U2523 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, S 
                           => n3587, Z => n1355);
   U2524 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, S 
                           => n3587, Z => n1354);
   U2525 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, S 
                           => n3587, Z => n1353);
   U2526 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, S 
                           => n4378, Z => n1352);
   U2527 : MUX2_X1 port map( A => n3197, B => n3309, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U2528 : MUX2_X1 port map( A => n3196, B => n3312, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U2529 : MUX2_X1 port map( A => n3195, B => n3315, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U2530 : MUX2_X1 port map( A => n3194, B => n3318, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_10_port);
   U2531 : MUX2_X1 port map( A => n3193, B => n3321, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_11_port);
   U2532 : MUX2_X1 port map( A => n3192, B => n3324, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_12_port);
   U2533 : MUX2_X1 port map( A => n3191, B => n3327, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_13_port);
   U2534 : MUX2_X1 port map( A => n3190, B => n3330, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_14_port);
   U2535 : MUX2_X1 port map( A => n3189, B => n3333, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_15_port);
   U2536 : MUX2_X1 port map( A => n3188, B => n3336, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_16_port);
   U2537 : MUX2_X1 port map( A => n3187, B => n3339, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_17_port);
   U2538 : MUX2_X1 port map( A => n3186, B => n3342, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_18_port);
   U2539 : MUX2_X1 port map( A => n3185, B => n3345, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_19_port);
   U2540 : MUX2_X1 port map( A => n3184, B => n3348, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_20_port);
   U2541 : MUX2_X1 port map( A => n3183, B => n3351, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_21_port);
   U2542 : MUX2_X1 port map( A => n3182, B => n3354, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_22_port);
   U2543 : MUX2_X1 port map( A => n3181, B => n3357, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_23_port);
   U2544 : MUX2_X1 port map( A => n3180, B => n3360, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_24_port);
   U2545 : MUX2_X1 port map( A => n3179, B => n3363, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U2546 : MUX2_X1 port map( A => n3178, B => n3366, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U2547 : MUX2_X1 port map( A => n3176, B => n3369, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U2548 : MUX2_X1 port map( A => n3175, B => n3372, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U2549 : MUX2_X1 port map( A => n3174, B => n3375, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U2550 : MUX2_X1 port map( A => n3173, B => n3378, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U2551 : MUX2_X1 port map( A => n3172, B => n3381, S => n4379, Z => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U2552 : MUX2_X1 port map( A => n3166, B => n3306, S => n3135, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U2553 : INV_X1 port map( A => n4127, ZN => n4380);
   U2554 : AOI22_X1 port map( A1 => n3241, A2 => n4380, B1 => n3156, B2 => 
                           n3404, ZN => n4381);
   U2555 : OAI21_X1 port map( B1 => n3261, B2 => n3467, A => n4381, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U2556 : INV_X1 port map( A => n4125, ZN => n4382);
   U2557 : AOI22_X1 port map( A1 => n4389, A2 => n4382, B1 => n3558, B2 => 
                           n3412, ZN => n4383);
   U2558 : OAI21_X1 port map( B1 => n3261, B2 => n3471, A => n4383, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U2559 : INV_X1 port map( A => n4123, ZN => n4384);
   U2560 : AOI22_X1 port map( A1 => n3241, A2 => n4384, B1 => n3156, B2 => 
                           n3420, ZN => n4385);
   U2561 : OAI21_X1 port map( B1 => n3559, B2 => n3476, A => n4385, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U2562 : AOI22_X1 port map( A1 => n3241, A2 => n4386, B1 => n3156, B2 => 
                           n3422, ZN => n4387);
   U2563 : OAI21_X1 port map( B1 => n3261, B2 => n3504, A => n4387, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U2564 : INV_X1 port map( A => n4122, ZN => n4388);
   U2565 : AOI22_X1 port map( A1 => n4389, A2 => n4388, B1 => n3558, B2 => 
                           n3424, ZN => n4390);
   U2566 : OAI21_X1 port map( B1 => n3261, B2 => n3478, A => n4390, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U2567 : AOI22_X1 port map( A1 => n3257, A2 => n3164, B1 => n3117, B2 => 
                           datapath_i_alu_output_val_i_0_port, ZN => n4391);
   U2568 : OAI21_X1 port map( B1 => n3255, B2 => n3539, A => n4391, ZN => n3628
                           );
   U2569 : MUX2_X1 port map( A => n3628, B => IRAM_ADDRESS_0_port, S => n3115, 
                           Z => n1388);
   U2570 : AOI22_X1 port map( A1 => n1388, A2 => n1727, B1 => n3383, B2 => 
                           n1802, ZN => n4392);
   U2571 : OAI21_X1 port map( B1 => n3540, B2 => n1507, A => n4392, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U2572 : INV_X1 port map( A => n4120, ZN => n4393);
   U2573 : AOI22_X1 port map( A1 => n3241, A2 => n4393, B1 => n3156, B2 => 
                           n3432, ZN => n4394);
   U2574 : OAI21_X1 port map( B1 => n3261, B2 => n3482, A => n4394, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U2575 : AOI22_X1 port map( A1 => n4395, A2 => n3241, B1 => n3156, B2 => 
                           n3440, ZN => n4396);
   U2576 : OAI21_X1 port map( B1 => n3549, B2 => n3261, A => n4396, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U2577 : AOI22_X1 port map( A1 => n4398, A2 => n3629, B1 => n4397, B2 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, ZN => 
                           n2547);
   U2578 : AOI22_X1 port map( A1 => n3115, A2 => n3161, B1 => n3554, B2 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, ZN => 
                           n1330);
   U2579 : AOI22_X1 port map( A1 => n1330, A2 => n1727, B1 => n3385, B2 => 
                           n1802, ZN => n4399);
   U2580 : OAI21_X1 port map( B1 => n3546, B2 => n1507, A => n4399, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U2581 : OAI211_X1 port map( C1 => datapath_i_new_pc_value_mem_stage_i_2_port
                           , C2 => datapath_i_new_pc_value_mem_stage_i_3_port, 
                           A => n3554, B => n4400, ZN => n4401);
   U2582 : NAND2_X1 port map( A1 => n3133, A2 => n4401, ZN => n1328);
   U2583 : AOI22_X1 port map( A1 => n1727, A2 => n1328, B1 => n3386, B2 => 
                           n1802, ZN => n4402);
   U2584 : OAI21_X1 port map( B1 => n3548, B2 => n1507, A => n4402, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U2585 : MUX2_X1 port map( A => n3209, B => n3160, S => n1801, Z => n1779);
   U2586 : AND4_X1 port map( A1 => n3584, A2 => n3582, A3 => n3578, A4 => n3112
                           , ZN => n4403);
   U2587 : NAND2_X1 port map( A1 => n3580, A2 => n4403, ZN => n3658);
   U2588 : AOI22_X1 port map( A1 => n3117, A2 => 
                           datapath_i_alu_output_val_i_11_port, B1 => n3457, B2
                           => n3452, ZN => n4404);
   U2589 : OAI21_X1 port map( B1 => n4128, B2 => n4425, A => n4404, ZN => n4114
                           );
   U2590 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_21_port, B1 => n3457, B2
                           => n3448, ZN => n4405);
   U2591 : OAI21_X1 port map( B1 => n4123, B2 => n4425, A => n4405, ZN => n4086
                           );
   U2592 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_19_port, B1 => n3457, B2
                           => n3556, ZN => n4406);
   U2593 : OAI21_X1 port map( B1 => n4124, B2 => n4425, A => n4406, ZN => n4085
                           );
   U2594 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_17_port, B1 => n3457, B2
                           => n3449, ZN => n4407);
   U2595 : OAI21_X1 port map( B1 => n4125, B2 => n4425, A => n4407, ZN => n4084
                           );
   U2596 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_13_port, B1 => n3457, B2
                           => n3451, ZN => n4408);
   U2597 : OAI21_X1 port map( B1 => n4127, B2 => n4425, A => n4408, ZN => n4083
                           );
   U2598 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_15_port, B1 => n3457, B2
                           => n3450, ZN => n4409);
   U2599 : OAI21_X1 port map( B1 => n4126, B2 => n4425, A => n4409, ZN => n4082
                           );
   U2600 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_23_port, B1 => n3457, B2
                           => n3447, ZN => n4410);
   U2601 : OAI21_X1 port map( B1 => n4122, B2 => n4425, A => n4410, ZN => n4081
                           );
   U2602 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_25_port, B1 => n3457, B2
                           => n3446, ZN => n4411);
   U2603 : OAI21_X1 port map( B1 => n4121, B2 => n4425, A => n4411, ZN => n4080
                           );
   U2604 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_27_port, B1 => n3443, B2
                           => n3445, ZN => n4412);
   U2605 : OAI21_X1 port map( B1 => n4120, B2 => n4425, A => n4412, ZN => n4079
                           );
   U2606 : AOI22_X1 port map( A1 => n3557, A2 => 
                           datapath_i_alu_output_val_i_29_port, B1 => n3443, B2
                           => n3444, ZN => n4413);
   U2607 : OAI21_X1 port map( B1 => n4119, B2 => n4425, A => n4413, ZN => n4078
                           );
   U2608 : OAI211_X1 port map( C1 => n4058, C2 => n4061, A => n4414, B => n4415
                           , ZN => n464);
   U2609 : NAND2_X1 port map( A1 => n4415, A2 => n4061, ZN => n2299);
   U2610 : AOI22_X1 port map( A1 => n1801, A2 => n4416, B1 => n4424, B2 => 
                           n4047, ZN => n4046);

end SYN_dlx_rtl;
