
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, dataout_mul_31_port, dataout_mul_30_port, 
      dataout_mul_29_port, dataout_mul_28_port, dataout_mul_27_port, 
      dataout_mul_26_port, dataout_mul_25_port, dataout_mul_24_port, 
      dataout_mul_23_port, dataout_mul_22_port, dataout_mul_21_port, 
      dataout_mul_20_port, dataout_mul_19_port, dataout_mul_18_port, 
      dataout_mul_17_port, dataout_mul_16_port, dataout_mul_15_port, 
      dataout_mul_13_port, dataout_mul_12_port, dataout_mul_11_port, 
      dataout_mul_10_port, dataout_mul_9_port, dataout_mul_8_port, 
      dataout_mul_7_port, dataout_mul_6_port, dataout_mul_5_port, 
      dataout_mul_4_port, dataout_mul_3_port, dataout_mul_2_port, 
      dataout_mul_1_port, dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521
      , N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n553, 
      boothmul_pipelined_i_muxes_in_7_232_port, 
      boothmul_pipelined_i_muxes_in_7_231_port, 
      boothmul_pipelined_i_muxes_in_7_230_port, 
      boothmul_pipelined_i_muxes_in_7_229_port, 
      boothmul_pipelined_i_muxes_in_7_228_port, 
      boothmul_pipelined_i_muxes_in_7_227_port, 
      boothmul_pipelined_i_muxes_in_7_226_port, 
      boothmul_pipelined_i_muxes_in_7_225_port, 
      boothmul_pipelined_i_muxes_in_7_224_port, 
      boothmul_pipelined_i_muxes_in_7_223_port, 
      boothmul_pipelined_i_muxes_in_7_222_port, 
      boothmul_pipelined_i_muxes_in_7_221_port, 
      boothmul_pipelined_i_muxes_in_7_220_port, 
      boothmul_pipelined_i_muxes_in_7_219_port, 
      boothmul_pipelined_i_muxes_in_7_218_port, 
      boothmul_pipelined_i_muxes_in_7_217_port, 
      boothmul_pipelined_i_muxes_in_7_76_port, 
      boothmul_pipelined_i_muxes_in_7_75_port, 
      boothmul_pipelined_i_muxes_in_7_74_port, 
      boothmul_pipelined_i_muxes_in_7_73_port, 
      boothmul_pipelined_i_muxes_in_7_72_port, 
      boothmul_pipelined_i_muxes_in_7_71_port, 
      boothmul_pipelined_i_muxes_in_7_70_port, 
      boothmul_pipelined_i_muxes_in_7_69_port, 
      boothmul_pipelined_i_muxes_in_7_68_port, 
      boothmul_pipelined_i_muxes_in_7_67_port, 
      boothmul_pipelined_i_muxes_in_7_66_port, 
      boothmul_pipelined_i_muxes_in_7_65_port, 
      boothmul_pipelined_i_muxes_in_7_64_port, 
      boothmul_pipelined_i_muxes_in_7_63_port, 
      boothmul_pipelined_i_muxes_in_7_62_port, 
      boothmul_pipelined_i_muxes_in_6_218_port, 
      boothmul_pipelined_i_muxes_in_6_217_port, 
      boothmul_pipelined_i_muxes_in_6_216_port, 
      boothmul_pipelined_i_muxes_in_6_215_port, 
      boothmul_pipelined_i_muxes_in_6_214_port, 
      boothmul_pipelined_i_muxes_in_6_213_port, 
      boothmul_pipelined_i_muxes_in_6_212_port, 
      boothmul_pipelined_i_muxes_in_6_211_port, 
      boothmul_pipelined_i_muxes_in_6_210_port, 
      boothmul_pipelined_i_muxes_in_6_209_port, 
      boothmul_pipelined_i_muxes_in_6_208_port, 
      boothmul_pipelined_i_muxes_in_6_207_port, 
      boothmul_pipelined_i_muxes_in_6_206_port, 
      boothmul_pipelined_i_muxes_in_6_205_port, 
      boothmul_pipelined_i_muxes_in_6_204_port, 
      boothmul_pipelined_i_muxes_in_6_203_port, 
      boothmul_pipelined_i_muxes_in_6_73_port, 
      boothmul_pipelined_i_muxes_in_6_72_port, 
      boothmul_pipelined_i_muxes_in_6_71_port, 
      boothmul_pipelined_i_muxes_in_6_70_port, 
      boothmul_pipelined_i_muxes_in_6_69_port, 
      boothmul_pipelined_i_muxes_in_6_68_port, 
      boothmul_pipelined_i_muxes_in_6_67_port, 
      boothmul_pipelined_i_muxes_in_6_66_port, 
      boothmul_pipelined_i_muxes_in_6_65_port, 
      boothmul_pipelined_i_muxes_in_6_64_port, 
      boothmul_pipelined_i_muxes_in_6_63_port, 
      boothmul_pipelined_i_muxes_in_6_62_port, 
      boothmul_pipelined_i_muxes_in_6_61_port, 
      boothmul_pipelined_i_muxes_in_6_60_port, 
      boothmul_pipelined_i_muxes_in_6_59_port, 
      boothmul_pipelined_i_muxes_in_6_58_port, 
      boothmul_pipelined_i_muxes_in_5_205_port, 
      boothmul_pipelined_i_muxes_in_5_204_port, 
      boothmul_pipelined_i_muxes_in_5_203_port, 
      boothmul_pipelined_i_muxes_in_5_202_port, 
      boothmul_pipelined_i_muxes_in_5_201_port, 
      boothmul_pipelined_i_muxes_in_5_200_port, 
      boothmul_pipelined_i_muxes_in_5_199_port, 
      boothmul_pipelined_i_muxes_in_5_198_port, 
      boothmul_pipelined_i_muxes_in_5_197_port, 
      boothmul_pipelined_i_muxes_in_5_196_port, 
      boothmul_pipelined_i_muxes_in_5_195_port, 
      boothmul_pipelined_i_muxes_in_5_194_port, 
      boothmul_pipelined_i_muxes_in_5_193_port, 
      boothmul_pipelined_i_muxes_in_5_192_port, 
      boothmul_pipelined_i_muxes_in_5_191_port, 
      boothmul_pipelined_i_muxes_in_5_190_port, 
      boothmul_pipelined_i_muxes_in_5_189_port, 
      boothmul_pipelined_i_muxes_in_5_68_port, 
      boothmul_pipelined_i_muxes_in_5_67_port, 
      boothmul_pipelined_i_muxes_in_5_66_port, 
      boothmul_pipelined_i_muxes_in_5_65_port, 
      boothmul_pipelined_i_muxes_in_5_64_port, 
      boothmul_pipelined_i_muxes_in_5_63_port, 
      boothmul_pipelined_i_muxes_in_5_62_port, 
      boothmul_pipelined_i_muxes_in_5_61_port, 
      boothmul_pipelined_i_muxes_in_5_60_port, 
      boothmul_pipelined_i_muxes_in_5_59_port, 
      boothmul_pipelined_i_muxes_in_5_58_port, 
      boothmul_pipelined_i_muxes_in_5_57_port, 
      boothmul_pipelined_i_muxes_in_5_56_port, 
      boothmul_pipelined_i_muxes_in_5_55_port, 
      boothmul_pipelined_i_muxes_in_5_54_port, 
      boothmul_pipelined_i_muxes_in_4_190_port, 
      boothmul_pipelined_i_muxes_in_4_189_port, 
      boothmul_pipelined_i_muxes_in_4_188_port, 
      boothmul_pipelined_i_muxes_in_4_187_port, 
      boothmul_pipelined_i_muxes_in_4_186_port, 
      boothmul_pipelined_i_muxes_in_4_185_port, 
      boothmul_pipelined_i_muxes_in_4_184_port, 
      boothmul_pipelined_i_muxes_in_4_183_port, 
      boothmul_pipelined_i_muxes_in_4_182_port, 
      boothmul_pipelined_i_muxes_in_4_181_port, 
      boothmul_pipelined_i_muxes_in_4_180_port, 
      boothmul_pipelined_i_muxes_in_4_179_port, 
      boothmul_pipelined_i_muxes_in_4_178_port, 
      boothmul_pipelined_i_muxes_in_4_177_port, 
      boothmul_pipelined_i_muxes_in_4_176_port, 
      boothmul_pipelined_i_muxes_in_4_175_port, 
      boothmul_pipelined_i_muxes_in_4_65_port, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_58_port, 
      boothmul_pipelined_i_muxes_in_4_57_port, 
      boothmul_pipelined_i_muxes_in_4_56_port, 
      boothmul_pipelined_i_muxes_in_4_55_port, 
      boothmul_pipelined_i_muxes_in_4_54_port, 
      boothmul_pipelined_i_muxes_in_4_53_port, 
      boothmul_pipelined_i_muxes_in_4_52_port, 
      boothmul_pipelined_i_muxes_in_4_51_port, 
      boothmul_pipelined_i_muxes_in_4_50_port, 
      boothmul_pipelined_i_muxes_in_3_177_port, 
      boothmul_pipelined_i_muxes_in_3_176_port, 
      boothmul_pipelined_i_muxes_in_3_175_port, 
      boothmul_pipelined_i_muxes_in_3_174_port, 
      boothmul_pipelined_i_muxes_in_3_173_port, 
      boothmul_pipelined_i_muxes_in_3_172_port, 
      boothmul_pipelined_i_muxes_in_3_171_port, 
      boothmul_pipelined_i_muxes_in_3_170_port, 
      boothmul_pipelined_i_muxes_in_3_169_port, 
      boothmul_pipelined_i_muxes_in_3_168_port, 
      boothmul_pipelined_i_muxes_in_3_167_port, 
      boothmul_pipelined_i_muxes_in_3_166_port, 
      boothmul_pipelined_i_muxes_in_3_165_port, 
      boothmul_pipelined_i_muxes_in_3_164_port, 
      boothmul_pipelined_i_muxes_in_3_163_port, 
      boothmul_pipelined_i_muxes_in_3_162_port, 
      boothmul_pipelined_i_muxes_in_3_161_port, 
      boothmul_pipelined_i_muxes_in_3_60_port, 
      boothmul_pipelined_i_muxes_in_3_59_port, 
      boothmul_pipelined_i_muxes_in_3_58_port, 
      boothmul_pipelined_i_muxes_in_3_57_port, 
      boothmul_pipelined_i_muxes_in_3_56_port, 
      boothmul_pipelined_i_muxes_in_3_55_port, 
      boothmul_pipelined_i_muxes_in_3_54_port, 
      boothmul_pipelined_i_muxes_in_3_53_port, 
      boothmul_pipelined_i_muxes_in_3_52_port, 
      boothmul_pipelined_i_muxes_in_3_51_port, 
      boothmul_pipelined_i_muxes_in_3_50_port, 
      boothmul_pipelined_i_muxes_in_3_49_port, 
      boothmul_pipelined_i_muxes_in_3_48_port, 
      boothmul_pipelined_i_muxes_in_3_47_port, 
      boothmul_pipelined_i_muxes_in_3_46_port, 
      boothmul_pipelined_i_sum_out_6_0_port, 
      boothmul_pipelined_i_sum_out_6_1_port, 
      boothmul_pipelined_i_sum_out_6_2_port, 
      boothmul_pipelined_i_sum_out_6_3_port, 
      boothmul_pipelined_i_sum_out_6_4_port, 
      boothmul_pipelined_i_sum_out_6_5_port, 
      boothmul_pipelined_i_sum_out_6_6_port, 
      boothmul_pipelined_i_sum_out_6_7_port, 
      boothmul_pipelined_i_sum_out_6_8_port, 
      boothmul_pipelined_i_sum_out_6_9_port, 
      boothmul_pipelined_i_sum_out_6_10_port, 
      boothmul_pipelined_i_sum_out_6_11_port, 
      boothmul_pipelined_i_sum_out_6_13_port, 
      boothmul_pipelined_i_sum_out_6_14_port, 
      boothmul_pipelined_i_sum_out_6_15_port, 
      boothmul_pipelined_i_sum_out_6_16_port, 
      boothmul_pipelined_i_sum_out_6_17_port, 
      boothmul_pipelined_i_sum_out_6_18_port, 
      boothmul_pipelined_i_sum_out_6_19_port, 
      boothmul_pipelined_i_sum_out_6_20_port, 
      boothmul_pipelined_i_sum_out_6_21_port, 
      boothmul_pipelined_i_sum_out_6_22_port, 
      boothmul_pipelined_i_sum_out_6_23_port, 
      boothmul_pipelined_i_sum_out_6_24_port, 
      boothmul_pipelined_i_sum_out_6_25_port, 
      boothmul_pipelined_i_sum_out_6_26_port, 
      boothmul_pipelined_i_sum_out_6_27_port, 
      boothmul_pipelined_i_sum_out_6_28_port, 
      boothmul_pipelined_i_sum_out_5_0_port, 
      boothmul_pipelined_i_sum_out_5_1_port, 
      boothmul_pipelined_i_sum_out_5_2_port, 
      boothmul_pipelined_i_sum_out_5_3_port, 
      boothmul_pipelined_i_sum_out_5_4_port, 
      boothmul_pipelined_i_sum_out_5_5_port, 
      boothmul_pipelined_i_sum_out_5_6_port, 
      boothmul_pipelined_i_sum_out_5_7_port, 
      boothmul_pipelined_i_sum_out_5_8_port, 
      boothmul_pipelined_i_sum_out_5_9_port, 
      boothmul_pipelined_i_sum_out_5_11_port, 
      boothmul_pipelined_i_sum_out_5_12_port, 
      boothmul_pipelined_i_sum_out_5_13_port, 
      boothmul_pipelined_i_sum_out_5_14_port, 
      boothmul_pipelined_i_sum_out_5_15_port, 
      boothmul_pipelined_i_sum_out_5_16_port, 
      boothmul_pipelined_i_sum_out_5_17_port, 
      boothmul_pipelined_i_sum_out_5_18_port, 
      boothmul_pipelined_i_sum_out_5_19_port, 
      boothmul_pipelined_i_sum_out_5_20_port, 
      boothmul_pipelined_i_sum_out_5_21_port, 
      boothmul_pipelined_i_sum_out_5_22_port, 
      boothmul_pipelined_i_sum_out_5_23_port, 
      boothmul_pipelined_i_sum_out_5_24_port, 
      boothmul_pipelined_i_sum_out_5_25_port, 
      boothmul_pipelined_i_sum_out_5_26_port, 
      boothmul_pipelined_i_sum_out_4_0_port, 
      boothmul_pipelined_i_sum_out_4_1_port, 
      boothmul_pipelined_i_sum_out_4_2_port, 
      boothmul_pipelined_i_sum_out_4_3_port, 
      boothmul_pipelined_i_sum_out_4_4_port, 
      boothmul_pipelined_i_sum_out_4_5_port, 
      boothmul_pipelined_i_sum_out_4_6_port, 
      boothmul_pipelined_i_sum_out_4_7_port, 
      boothmul_pipelined_i_sum_out_4_9_port, 
      boothmul_pipelined_i_sum_out_4_10_port, 
      boothmul_pipelined_i_sum_out_4_11_port, 
      boothmul_pipelined_i_sum_out_4_12_port, 
      boothmul_pipelined_i_sum_out_4_13_port, 
      boothmul_pipelined_i_sum_out_4_14_port, 
      boothmul_pipelined_i_sum_out_4_15_port, 
      boothmul_pipelined_i_sum_out_4_16_port, 
      boothmul_pipelined_i_sum_out_4_17_port, 
      boothmul_pipelined_i_sum_out_4_18_port, 
      boothmul_pipelined_i_sum_out_4_19_port, 
      boothmul_pipelined_i_sum_out_4_20_port, 
      boothmul_pipelined_i_sum_out_4_21_port, 
      boothmul_pipelined_i_sum_out_4_22_port, 
      boothmul_pipelined_i_sum_out_4_23_port, 
      boothmul_pipelined_i_sum_out_4_24_port, 
      boothmul_pipelined_i_sum_out_3_0_port, 
      boothmul_pipelined_i_sum_out_3_1_port, 
      boothmul_pipelined_i_sum_out_3_2_port, 
      boothmul_pipelined_i_sum_out_3_3_port, 
      boothmul_pipelined_i_sum_out_3_4_port, 
      boothmul_pipelined_i_sum_out_3_5_port, 
      boothmul_pipelined_i_sum_out_3_7_port, 
      boothmul_pipelined_i_sum_out_3_8_port, 
      boothmul_pipelined_i_sum_out_3_9_port, 
      boothmul_pipelined_i_sum_out_3_10_port, 
      boothmul_pipelined_i_sum_out_3_11_port, 
      boothmul_pipelined_i_sum_out_3_12_port, 
      boothmul_pipelined_i_sum_out_3_13_port, 
      boothmul_pipelined_i_sum_out_3_14_port, 
      boothmul_pipelined_i_sum_out_3_15_port, 
      boothmul_pipelined_i_sum_out_3_16_port, 
      boothmul_pipelined_i_sum_out_3_17_port, 
      boothmul_pipelined_i_sum_out_3_18_port, 
      boothmul_pipelined_i_sum_out_3_19_port, 
      boothmul_pipelined_i_sum_out_3_20_port, 
      boothmul_pipelined_i_sum_out_3_21_port, 
      boothmul_pipelined_i_sum_out_3_22_port, 
      boothmul_pipelined_i_sum_out_2_0_port, 
      boothmul_pipelined_i_sum_out_2_1_port, 
      boothmul_pipelined_i_sum_out_2_2_port, 
      boothmul_pipelined_i_sum_out_2_3_port, 
      boothmul_pipelined_i_sum_out_2_5_port, 
      boothmul_pipelined_i_sum_out_2_6_port, 
      boothmul_pipelined_i_sum_out_2_7_port, 
      boothmul_pipelined_i_sum_out_2_8_port, 
      boothmul_pipelined_i_sum_out_2_9_port, 
      boothmul_pipelined_i_sum_out_2_10_port, 
      boothmul_pipelined_i_sum_out_2_11_port, 
      boothmul_pipelined_i_sum_out_2_12_port, 
      boothmul_pipelined_i_sum_out_2_13_port, 
      boothmul_pipelined_i_sum_out_2_14_port, 
      boothmul_pipelined_i_sum_out_2_15_port, 
      boothmul_pipelined_i_sum_out_2_16_port, 
      boothmul_pipelined_i_sum_out_2_17_port, 
      boothmul_pipelined_i_sum_out_2_18_port, 
      boothmul_pipelined_i_sum_out_2_19_port, 
      boothmul_pipelined_i_sum_out_2_20_port, 
      boothmul_pipelined_i_sum_out_1_0_port, 
      boothmul_pipelined_i_sum_out_1_3_port, 
      boothmul_pipelined_i_sum_out_1_4_port, 
      boothmul_pipelined_i_sum_out_1_5_port, 
      boothmul_pipelined_i_sum_out_1_6_port, 
      boothmul_pipelined_i_sum_out_1_7_port, 
      boothmul_pipelined_i_sum_out_1_8_port, 
      boothmul_pipelined_i_sum_out_1_9_port, 
      boothmul_pipelined_i_sum_out_1_10_port, 
      boothmul_pipelined_i_sum_out_1_11_port, 
      boothmul_pipelined_i_sum_out_1_12_port, 
      boothmul_pipelined_i_sum_out_1_13_port, 
      boothmul_pipelined_i_sum_out_1_14_port, 
      boothmul_pipelined_i_sum_out_1_15_port, 
      boothmul_pipelined_i_sum_out_1_16_port, 
      boothmul_pipelined_i_sum_out_1_17_port, 
      boothmul_pipelined_i_sum_out_1_18_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_13_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_11_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_6_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_15_port, 
      boothmul_pipelined_i_multiplicand_pip_5_9_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_5_12_port, 
      boothmul_pipelined_i_multiplicand_pip_5_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_14_port, 
      boothmul_pipelined_i_multiplicand_pip_5_15_port, 
      boothmul_pipelined_i_multiplicand_pip_4_7_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_4_10_port, 
      boothmul_pipelined_i_multiplicand_pip_4_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_12_port, 
      boothmul_pipelined_i_multiplicand_pip_4_13_port, 
      boothmul_pipelined_i_multiplicand_pip_4_14_port, 
      boothmul_pipelined_i_multiplicand_pip_4_15_port, 
      boothmul_pipelined_i_multiplicand_pip_3_5_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_3_8_port, 
      boothmul_pipelined_i_multiplicand_pip_3_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_10_port, 
      boothmul_pipelined_i_multiplicand_pip_3_11_port, 
      boothmul_pipelined_i_multiplicand_pip_3_12_port, 
      boothmul_pipelined_i_multiplicand_pip_3_13_port, 
      boothmul_pipelined_i_multiplicand_pip_3_14_port, 
      boothmul_pipelined_i_multiplicand_pip_3_15_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_multiplicand_pip_2_6_port, 
      boothmul_pipelined_i_multiplicand_pip_2_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_8_port, 
      boothmul_pipelined_i_multiplicand_pip_2_9_port, 
      boothmul_pipelined_i_multiplicand_pip_2_10_port, 
      boothmul_pipelined_i_multiplicand_pip_2_11_port, 
      boothmul_pipelined_i_multiplicand_pip_2_12_port, 
      boothmul_pipelined_i_multiplicand_pip_2_13_port, 
      boothmul_pipelined_i_multiplicand_pip_2_14_port, 
      boothmul_pipelined_i_multiplicand_pip_2_15_port, 
      boothmul_pipelined_i_muxes_in_0_119_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n3076, 
      n3077, n3078, n3079, n3080, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n1995, n1996, 
      n1997, n5121, n5122, n5123, n5124, n5126, n5127, n5128, n5129, n5130, 
      n5131, n5132, n5133, n5134, n1991, n7164, n7165, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1992, n1993, n1994, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n11231, n11232, n11233, 
      n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, 
      n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, 
      n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, 
      n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, 
      n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, 
      n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, 
      n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, 
      n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, 
      n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, 
      n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, 
      n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, 
      n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, 
      n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, 
      n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, 
      n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, 
      n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, 
      n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, 
      n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, 
      n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, 
      n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, 
      n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, 
      n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, 
      n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, 
      n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, 
      n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, 
      n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, 
      n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, 
      n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, 
      n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, 
      n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, 
      n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, 
      n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, 
      n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, 
      n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, 
      n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, 
      n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, 
      n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, 
      n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, 
      n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, 
      n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, 
      n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, 
      n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, 
      n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, 
      n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, 
      n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, 
      n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, 
      n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, 
      n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, 
      n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, 
      n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, 
      n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, 
      n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, 
      n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, 
      n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, 
      n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, 
      n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, 
      n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, 
      n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, 
      n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, 
      n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, 
      n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, 
      n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, 
      n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, 
      n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, 
      n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, 
      n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, 
      n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, 
      n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, 
      n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, 
      n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, 
      n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, 
      n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, 
      n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, 
      n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, 
      n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, 
      n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, 
      n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, 
      n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, 
      n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, 
      n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, 
      n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, 
      n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, 
      n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, 
      n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, 
      n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, 
      n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, 
      n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, 
      n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, 
      n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, 
      n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, 
      n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, 
      n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, 
      n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, 
      n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, 
      n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, 
      n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, 
      n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, 
      n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, 
      n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, 
      n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, 
      n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, 
      n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, 
      n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, 
      n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, 
      n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, 
      n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, 
      n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, 
      n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, 
      n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, 
      n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, 
      n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, 
      n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, 
      n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, 
      n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, 
      n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, 
      n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, 
      n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, 
      n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, 
      n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, 
      n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, 
      n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, 
      n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, 
      n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, 
      n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, 
      n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, 
      n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, 
      n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, 
      n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, 
      n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, 
      n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, 
      n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, 
      n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, 
      n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, 
      n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, 
      n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, 
      n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, 
      n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, 
      n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, 
      n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, 
      n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, 
      n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, 
      n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, 
      n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, 
      n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, 
      n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, 
      n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, 
      n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, 
      n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, 
      n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, 
      n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, 
      n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, 
      n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, 
      n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, 
      n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, 
      n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, 
      n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, 
      n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, 
      n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, 
      n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, 
      n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, 
      n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, 
      n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, 
      n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, 
      n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, 
      n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, 
      n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, 
      n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, 
      n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, 
      n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, 
      n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, 
      n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, 
      n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, 
      n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, 
      n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, 
      n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, 
      n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, 
      n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, 
      n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, 
      n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, 
      n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, 
      n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, 
      n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, 
      n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, 
      n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, 
      n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, 
      n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, 
      n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, 
      n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, 
      n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, 
      n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, 
      n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, 
      n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, 
      n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, 
      n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, 
      n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, 
      n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, 
      n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, 
      n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, 
      n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, 
      n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, 
      n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, 
      n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, 
      n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, 
      n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, 
      n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, 
      n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, 
      n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, 
      n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, 
      n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, 
      n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, 
      n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, 
      n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, 
      n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, 
      n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, 
      n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, 
      n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, 
      n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, 
      n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, 
      n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, 
      n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, 
      n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, 
      n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, 
      n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, 
      n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, 
      n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, 
      n13259, n13260, n13261, n13262, n13263, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, 
      n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, 
      n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, 
      n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348 : 
      std_logic;

begin
   
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n2009, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n13259, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n2009, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n2009, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n13259, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n2009, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n13259, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n2009, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n2009, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n2009, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n2009, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n2009, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n13259, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n2009, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n13259, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n2009, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n13259, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n2009, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n2009, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n2009, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n13259, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n2009, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n13259, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n13259, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n13259, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n2009, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => n13263, GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => n13262, GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => n13261, GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => DATA1(3), GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => n13260, GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, CK 
                           => clk, RN => n11241, Q => n13258, QN => n7165);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, CK 
                           => clk, RN => n11241, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, QN 
                           => n_1004);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => n11245, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, QN 
                           => n_1005);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, CK 
                           => clk, RN => n11238, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, QN 
                           => n_1006);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, CK 
                           => clk, RN => n11241, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, QN 
                           => n_1007);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, CK 
                           => clk, RN => n11240, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, QN 
                           => n3080);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, CK 
                           => clk, RN => n11239, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, QN 
                           => n_1008);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => n11242, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, QN 
                           => n_1009);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, CK 
                           => clk, RN => n11238, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, QN 
                           => n_1010);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, CK 
                           => clk, RN => n11244, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, QN 
                           => n_1011);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, CK 
                           => clk, RN => n11231, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, QN 
                           => n_1012);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, QN 
                           => n_1013);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, CK 
                           => clk, RN => n11240, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, QN 
                           => n3079);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, CK 
                           => clk, RN => n11233, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, QN 
                           => n_1014);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => n11240, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, QN 
                           => n_1015);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, CK 
                           => clk, RN => n11231, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, QN 
                           => n_1016);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, CK 
                           => clk, RN => n11238, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, QN 
                           => n_1017);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, CK 
                           => clk, RN => n11245, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, QN 
                           => n_1018);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, CK 
                           => clk, RN => n11244, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, QN 
                           => n_1019);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, CK 
                           => clk, RN => n11238, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, QN 
                           => n_1020);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, CK 
                           => clk, RN => n11232, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, QN 
                           => n_1021);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, CK 
                           => clk, RN => n11243, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, QN 
                           => n3078);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, CK 
                           => clk, RN => n11239, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, QN 
                           => n_1022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => n11242, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, QN 
                           => n_1023);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, CK 
                           => clk, RN => n11239, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, QN 
                           => n_1024);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, CK 
                           => clk, RN => n11231, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, QN 
                           => n_1025);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, CK 
                           => clk, RN => n11235, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, QN 
                           => n_1026);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, CK 
                           => clk, RN => n11240, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, QN 
                           => n_1027);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, CK 
                           => clk, RN => n11234, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, QN 
                           => n_1028);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, CK 
                           => clk, RN => n11239, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, QN 
                           => n_1029);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, CK 
                           => clk, RN => n11241, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, QN 
                           => n_1030);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, CK 
                           => clk, RN => n11244, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, QN 
                           => n_1031);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, CK 
                           => clk, RN => n11243, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, QN 
                           => n3082);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, CK 
                           => clk, RN => n11231, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, QN 
                           => n_1032);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, CK 
                           => clk, RN => n11240, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, QN 
                           => n_1033);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_15_port, CK => clk, RN => n11239, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, QN 
                           => n_1034);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_14_port, CK => clk, RN => n11240, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, QN 
                           => n_1035);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_13_port, CK => clk, RN => n11233, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, QN 
                           => n_1036);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_12_port, CK => clk, RN => n11231, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, QN 
                           => n_1037);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_11_port, CK => clk, RN => n11233, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, QN 
                           => n_1038);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_10_port, CK => clk, RN => n11242, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, QN 
                           => n_1039);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_9_port, CK => clk, RN => n11243, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, QN 
                           => n_1040);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_8_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, QN 
                           => n_1041);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_7_port, CK => clk, RN => n11245, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, QN 
                           => n_1042);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_6_port, CK => clk, RN => n11236, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, QN 
                           => n_1043);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_5_port, CK => clk, RN => n11243, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, QN 
                           => n3076);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_4_port, CK => clk, RN => n11244, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, QN 
                           => n_1044);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_3_port, CK => clk, RN => n11233, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, QN 
                           => n_1045);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_28_port, CK => clk
                           , RN => n11232, Q => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, QN => 
                           n_1046);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_27_port, CK => clk
                           , RN => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, QN => 
                           n_1047);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_26_port, CK => clk
                           , RN => n11235, Q => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, QN => 
                           n_1048);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_25_port, CK => clk
                           , RN => n11237, Q => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, QN => 
                           n_1049);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_24_port, CK => clk
                           , RN => n11242, Q => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, QN => 
                           n_1050);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_23_port, CK => clk
                           , RN => n11236, Q => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, QN => 
                           n_1051);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_22_port, CK => clk
                           , RN => n11238, Q => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, QN => 
                           n_1052);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_21_port, CK => clk
                           , RN => n11240, Q => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, QN => 
                           n_1053);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_20_port, CK => clk
                           , RN => n11244, Q => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, QN => 
                           n_1054);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_19_port, CK => clk
                           , RN => n11243, Q => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, QN => 
                           n_1055);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_18_port, CK => clk
                           , RN => n11232, Q => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, QN => 
                           n_1056);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_17_port, CK => clk
                           , RN => n11240, Q => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, QN => 
                           n_1057);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_16_port, CK => clk
                           , RN => n11231, Q => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, QN => 
                           n_1058);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_15_port, CK => clk
                           , RN => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, QN => 
                           n_1059);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_14_port, CK => clk
                           , RN => n11243, Q => n_1060, QN => n5126);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_13_port, CK => clk
                           , RN => n11236, Q => dataout_mul_13_port, QN => 
                           n_1061);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => n3095, CK => clk, RN => n11240, Q => 
                           dataout_mul_12_port, QN => n_1062);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_11_port, CK => clk
                           , RN => n11236, Q => dataout_mul_11_port, QN => 
                           n_1063);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_10_port, CK => clk
                           , RN => n11241, Q => dataout_mul_10_port, QN => 
                           n_1064);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_9_port, CK => clk, RN
                           => n11240, Q => dataout_mul_9_port, QN => n_1065);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_8_port, CK => clk, RN
                           => n11237, Q => dataout_mul_8_port, QN => n_1066);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_7_port, CK => clk, RN
                           => n11232, Q => dataout_mul_7_port, QN => n_1067);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_6_port, CK => clk, RN
                           => n11236, Q => dataout_mul_6_port, QN => n_1068);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_5_port, CK => clk, RN
                           => n11241, Q => dataout_mul_5_port, QN => n_1069);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_4_port, CK => clk, RN
                           => n11238, Q => dataout_mul_4_port, QN => n_1070);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_3_port, CK => clk, RN
                           => n11244, Q => dataout_mul_3_port, QN => n_1071);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_2_port, CK => clk, RN
                           => n11233, Q => dataout_mul_2_port, QN => n_1072);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_1_port, CK => clk, RN
                           => n11241, Q => dataout_mul_1_port, QN => n_1073);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_0_port, CK => clk, RN
                           => n11242, Q => dataout_mul_0_port, QN => n_1074);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_58_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_7_62_port, QN => 
                           n_1075);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_59_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_63_port, QN => 
                           n_1076);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_60_port, CK => 
                           clk, RN => n11240, Q => 
                           boothmul_pipelined_i_muxes_in_7_64_port, QN => 
                           n_1077);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_61_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_7_65_port, QN => 
                           n_1078);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_62_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_7_66_port, QN => 
                           n_1079);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_63_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_7_67_port, QN => 
                           n_1080);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_64_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_7_68_port, QN => 
                           n_1081);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_65_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_7_69_port, QN => 
                           n_1082);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_66_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_7_70_port, QN => 
                           n_1083);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_67_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_7_71_port, QN => 
                           n_1084);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_68_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_7_72_port, QN => 
                           n_1085);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_69_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_7_73_port, QN => 
                           n_1086);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_178_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_70_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_7_74_port, QN => 
                           n_1087);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_177_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_71_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_7_75_port, QN => 
                           n_1088);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_176_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_72_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_7_76_port, QN => 
                           n_1089);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_203_port, CK => 
                           clk, RN => n11233, Q => 
                           boothmul_pipelined_i_muxes_in_7_217_port, QN => 
                           n_1090);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_204_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_7_218_port, QN => 
                           n_1091);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_205_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_7_219_port, QN => 
                           n_1092);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_42_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_206_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_7_220_port, QN => 
                           n_1093);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_41_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_207_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_7_221_port, QN => 
                           n_1094);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_40_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_208_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_7_222_port, QN => 
                           n_1095);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_39_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_209_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_7_223_port, QN => 
                           n_1096);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_38_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_210_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_224_port, QN => 
                           n_1097);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_37_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_211_port, CK => 
                           clk, RN => n11240, Q => 
                           boothmul_pipelined_i_muxes_in_7_225_port, QN => 
                           n_1098);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_36_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_212_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_7_226_port, QN => 
                           n_1099);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_35_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_213_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_7_227_port, QN => 
                           n_1100);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_34_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_214_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_7_228_port, QN => 
                           n_1101);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_33_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_215_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_7_229_port, QN => 
                           n_1102);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_216_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_7_230_port, QN => 
                           n_1103);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_217_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_7_231_port, QN => 
                           n_1104);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_218_port, CK => 
                           clk, RN => n11233, Q => 
                           boothmul_pipelined_i_muxes_in_7_232_port, QN => 
                           n_1105);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => n11243, Q => n_1106, QN => n5134);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_26_port, CK => clk
                           , RN => n11233, Q => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, QN => 
                           n_1107);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_25_port, CK => clk
                           , RN => n11234, Q => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, QN => 
                           n_1108);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_24_port, CK => clk
                           , RN => n11233, Q => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, QN => 
                           n_1109);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_23_port, CK => clk
                           , RN => n11233, Q => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, QN => 
                           n_1110);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_22_port, CK => clk
                           , RN => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, QN => 
                           n_1111);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_21_port, CK => clk
                           , RN => n11239, Q => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, QN => 
                           n_1112);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, QN => 
                           n_1113);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_19_port, CK => clk
                           , RN => n11238, Q => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, QN => 
                           n_1114);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_18_port, CK => clk
                           , RN => n11238, Q => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, QN => 
                           n_1115);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_17_port, CK => clk
                           , RN => n11239, Q => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, QN => 
                           n_1116);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_16_port, CK => clk
                           , RN => n11236, Q => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, QN => 
                           n_1117);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_15_port, CK => clk
                           , RN => n11237, Q => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, QN => 
                           n_1118);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_14_port, CK => clk
                           , RN => n11241, Q => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, QN => 
                           n_1119);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_13_port, CK => clk
                           , RN => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, QN => 
                           n_1120);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_12_port, CK => clk
                           , RN => n11244, Q => n_1121, QN => n5133);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_11_port, CK => clk
                           , RN => n11236, Q => 
                           boothmul_pipelined_i_sum_out_6_11_port, QN => n_1122
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => n3094, CK => clk, RN => n11239, Q => 
                           boothmul_pipelined_i_sum_out_6_10_port, QN => n_1123
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_9_port, CK => clk, RN
                           => n11235, Q => 
                           boothmul_pipelined_i_sum_out_6_9_port, QN => n_1124)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_8_port, CK => clk, RN
                           => n11236, Q => 
                           boothmul_pipelined_i_sum_out_6_8_port, QN => n_1125)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_7_port, CK => clk, RN
                           => n11233, Q => 
                           boothmul_pipelined_i_sum_out_6_7_port, QN => n_1126)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_6_6_port, QN => n_1127)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_5_port, CK => clk, RN
                           => n11241, Q => 
                           boothmul_pipelined_i_sum_out_6_5_port, QN => n_1128)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_4_port, CK => clk, RN
                           => n11239, Q => 
                           boothmul_pipelined_i_sum_out_6_4_port, QN => n_1129)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_3_port, CK => clk, RN
                           => n11241, Q => 
                           boothmul_pipelined_i_sum_out_6_3_port, QN => n_1130)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_2_port, CK => clk, RN
                           => n11234, Q => 
                           boothmul_pipelined_i_sum_out_6_2_port, QN => n_1131)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_1_port, CK => clk, RN
                           => n11238, Q => 
                           boothmul_pipelined_i_sum_out_6_1_port, QN => n_1132)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_0_port, CK => clk, RN
                           => n11236, Q => 
                           boothmul_pipelined_i_sum_out_6_0_port, QN => n_1133)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_54_port, CK => 
                           clk, RN => n11240, Q => 
                           boothmul_pipelined_i_muxes_in_6_58_port, QN => n5129
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_55_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_6_59_port, QN => 
                           n_1134);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_56_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_6_60_port, QN => 
                           n_1135);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_57_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_6_61_port, QN => 
                           n_1136);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_58_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_6_62_port, QN => 
                           n_1137);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_59_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_6_63_port, QN => 
                           n_1138);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_60_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_64_port, QN => 
                           n_1139);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_61_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_6_65_port, QN => 
                           n_1140);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_62_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_6_66_port, QN => 
                           n_1141);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_63_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_6_67_port, QN => 
                           n_1142);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_64_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_6_68_port, QN => 
                           n_1143);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_65_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_6_69_port, QN => 
                           n_1144);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_66_port, CK => 
                           clk, RN => n11241, Q => 
                           boothmul_pipelined_i_muxes_in_6_70_port, QN => 
                           n_1145);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_67_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_6_71_port, QN => 
                           n_1146);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_68_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_6_72_port, QN => 
                           n_1147);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_205_port, CK => 
                           clk, RN => n11240, Q => 
                           boothmul_pipelined_i_muxes_in_6_73_port, QN => n5123
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_189_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_6_203_port, QN => 
                           n_1148);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_190_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_6_204_port, QN => 
                           n_1149);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_191_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_6_205_port, QN => 
                           n_1150);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_56_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_192_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_6_206_port, QN => 
                           n_1151);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_55_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_193_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_6_207_port, QN => 
                           n_1152);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_54_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_194_port, CK => 
                           clk, RN => n11240, Q => 
                           boothmul_pipelined_i_muxes_in_6_208_port, QN => 
                           n_1153);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_53_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_195_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_6_209_port, QN => 
                           n_1154);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_52_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_196_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_6_210_port, QN => 
                           n_1155);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_51_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_197_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_6_211_port, QN => 
                           n_1156);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_50_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_198_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_6_212_port, QN => 
                           n_1157);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_49_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_199_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_6_213_port, QN => 
                           n_1158);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_48_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_200_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_6_214_port, QN => 
                           n_1159);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_47_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_201_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_6_215_port, QN => 
                           n_1160);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_46_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_202_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_6_216_port, QN => 
                           n_1161);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_203_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_6_217_port, QN => 
                           n_1162);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_204_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_6_218_port, QN => 
                           n_1163);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_24_port, CK => clk
                           , RN => n11236, Q => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, QN => 
                           n_1164);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_23_port, CK => clk
                           , RN => n11237, Q => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, QN => 
                           n_1165);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_22_port, CK => clk
                           , RN => n11239, Q => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, QN => 
                           n_1166);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_21_port, CK => clk
                           , RN => n11241, Q => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, QN => 
                           n_1167);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_20_port, CK => clk
                           , RN => n11243, Q => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, QN => 
                           n_1168);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_19_port, CK => clk
                           , RN => n11236, Q => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, QN => 
                           n_1169);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_18_port, CK => clk
                           , RN => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, QN => 
                           n_1170);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_17_port, CK => clk
                           , RN => n11242, Q => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, QN => 
                           n_1171);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_16_port, CK => clk
                           , RN => n11241, Q => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, QN => 
                           n_1172);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_15_port, CK => clk
                           , RN => n11243, Q => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, QN => 
                           n_1173);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_14_port, CK => clk
                           , RN => n11235, Q => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, QN => 
                           n_1174);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_13_port, CK => clk
                           , RN => n11240, Q => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, QN => 
                           n_1175);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_12_port, CK => clk
                           , RN => n11242, Q => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, QN => 
                           n_1176);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_11_port, CK => clk
                           , RN => n11241, Q => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, QN => 
                           n_1177);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_10_port, CK => clk
                           , RN => n11231, Q => n_1178, QN => n5132);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_9_port, CK => clk, RN
                           => n11241, Q => 
                           boothmul_pipelined_i_sum_out_5_9_port, QN => n_1179)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           n3093, CK => clk, RN => n11233, Q => 
                           boothmul_pipelined_i_sum_out_5_8_port, QN => n_1180)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_7_port, CK => clk, RN
                           => n11231, Q => 
                           boothmul_pipelined_i_sum_out_5_7_port, QN => n_1181)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_6_port, QN => n_1182)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_5_port, CK => clk, RN
                           => n11242, Q => 
                           boothmul_pipelined_i_sum_out_5_5_port, QN => n_1183)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_4_port, CK => clk, RN
                           => n11240, Q => 
                           boothmul_pipelined_i_sum_out_5_4_port, QN => n_1184)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_3_port, CK => clk, RN
                           => n11234, Q => 
                           boothmul_pipelined_i_sum_out_5_3_port, QN => n_1185)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_2_port, CK => clk, RN
                           => n11234, Q => 
                           boothmul_pipelined_i_sum_out_5_2_port, QN => n_1186)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_1_port, CK => clk, RN
                           => n11241, Q => 
                           boothmul_pipelined_i_sum_out_5_1_port, QN => n_1187)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_0_port, CK => clk, RN
                           => n11238, Q => 
                           boothmul_pipelined_i_sum_out_5_0_port, QN => n_1188)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_50_port, CK => 
                           clk, RN => n11233, Q => 
                           boothmul_pipelined_i_muxes_in_5_54_port, QN => n5128
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_51_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_5_55_port, QN => 
                           n_1189);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_52_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_5_56_port, QN => 
                           n_1190);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_53_port, CK => 
                           clk, RN => n11240, Q => 
                           boothmul_pipelined_i_muxes_in_5_57_port, QN => 
                           n_1191);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_54_port, CK => 
                           clk, RN => n11241, Q => 
                           boothmul_pipelined_i_muxes_in_5_58_port, QN => 
                           n_1192);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_55_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_5_59_port, QN => 
                           n_1193);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_56_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_5_60_port, QN => 
                           n_1194);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_57_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_5_61_port, QN => 
                           n_1195);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_58_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_5_62_port, QN => 
                           n_1196);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_59_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_5_63_port, QN => 
                           n_1197);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_60_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_5_64_port, QN => 
                           n_1198);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_61_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_5_65_port, QN => 
                           n_1199);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_62_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_5_66_port, QN => 
                           n_1200);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_63_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_5_67_port, QN => 
                           n_1201);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_64_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_5_68_port, QN => 
                           n_1202);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_175_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_5_189_port, QN => 
                           n_1203);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_176_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_5_190_port, QN => 
                           n_1204);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_177_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_5_191_port, QN => 
                           n_1205);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_178_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_5_192_port, QN => 
                           n_1206);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_179_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_5_193_port, QN => 
                           n_1207);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_180_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_5_194_port, QN => 
                           n_1208);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_181_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_5_195_port, QN => 
                           n_1209);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_182_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_5_196_port, QN => 
                           n_1210);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_183_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_5_197_port, QN => 
                           n_1211);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_184_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_5_198_port, QN => 
                           n_1212);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_185_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_5_199_port, QN => 
                           n_1213);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_186_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_5_200_port, QN => 
                           n_1214);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_187_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_5_201_port, QN => 
                           n_1215);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_188_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_5_202_port, QN => 
                           n_1216);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_189_port, CK => 
                           clk, RN => n11245, Q => 
                           boothmul_pipelined_i_muxes_in_5_203_port, QN => 
                           n_1217);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_190_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_5_204_port, QN => 
                           n_1218);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_65_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_5_205_port, QN => 
                           n5122);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_22_port, CK => clk
                           , RN => n11241, Q => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, QN => 
                           n_1219);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_21_port, CK => clk
                           , RN => n11244, Q => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, QN => 
                           n_1220);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_20_port, CK => clk
                           , RN => n11234, Q => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, QN => 
                           n_1221);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_19_port, CK => clk
                           , RN => n11232, Q => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, QN => 
                           n_1222);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_18_port, CK => clk
                           , RN => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, QN => 
                           n_1223);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_17_port, CK => clk
                           , RN => n11236, Q => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, QN => 
                           n_1224);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_16_port, CK => clk
                           , RN => n11244, Q => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, QN => 
                           n_1225);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_15_port, CK => clk
                           , RN => n11240, Q => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, QN => 
                           n_1226);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_14_port, CK => clk
                           , RN => n11244, Q => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, QN => 
                           n_1227);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_13_port, CK => clk
                           , RN => n11232, Q => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, QN => 
                           n_1228);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, QN => 
                           n_1229);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_11_port, CK => clk
                           , RN => n11235, Q => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, QN => 
                           n_1230);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_10_port, CK => clk
                           , RN => n11231, Q => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, QN => 
                           n_1231);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_9_port, CK => clk, RN
                           => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, QN => n_1232
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_8_port, CK => clk, RN
                           => n11244, Q => n_1233, QN => n5131);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_7_port, CK => clk, RN
                           => n11241, Q => 
                           boothmul_pipelined_i_sum_out_4_7_port, QN => n_1234)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           n3092, CK => clk, RN => n11242, Q => 
                           boothmul_pipelined_i_sum_out_4_6_port, QN => n_1235)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_5_port, CK => clk, RN
                           => n11237, Q => 
                           boothmul_pipelined_i_sum_out_4_5_port, QN => n_1236)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_4_port, CK => clk, RN
                           => n11239, Q => 
                           boothmul_pipelined_i_sum_out_4_4_port, QN => n_1237)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_3_port, CK => clk, RN
                           => n11244, Q => 
                           boothmul_pipelined_i_sum_out_4_3_port, QN => n_1238)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_2_port, CK => clk, RN
                           => n11237, Q => 
                           boothmul_pipelined_i_sum_out_4_2_port, QN => n_1239)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_1_port, CK => clk, RN
                           => n11240, Q => 
                           boothmul_pipelined_i_sum_out_4_1_port, QN => n_1240)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_0_port, CK => clk, RN
                           => n11240, Q => 
                           boothmul_pipelined_i_sum_out_4_0_port, QN => n_1241)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_46_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_4_50_port, QN => n5127
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_47_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_4_51_port, QN => 
                           n_1242);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_48_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_4_52_port, QN => 
                           n_1243);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_49_port, CK => 
                           clk, RN => n11233, Q => 
                           boothmul_pipelined_i_muxes_in_4_53_port, QN => 
                           n_1244);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_50_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_54_port, QN => 
                           n_1245);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_51_port, CK => 
                           clk, RN => n11241, Q => 
                           boothmul_pipelined_i_muxes_in_4_55_port, QN => 
                           n_1246);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_52_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_4_56_port, QN => 
                           n_1247);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_53_port, CK => 
                           clk, RN => n11241, Q => 
                           boothmul_pipelined_i_muxes_in_4_57_port, QN => 
                           n_1248);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_54_port, CK => 
                           clk, RN => n11233, Q => 
                           boothmul_pipelined_i_muxes_in_4_58_port, QN => 
                           n_1249);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_55_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port, QN => 
                           n_1250);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_56_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port, QN => 
                           n_1251);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_57_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port, QN => 
                           n_1252);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_58_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port, QN => 
                           n_1253);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_59_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port, QN => 
                           n_1254);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_60_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port, QN => 
                           n_1255);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_177_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_4_65_port, QN => n5121
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_161_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_4_175_port, QN => 
                           n_1256);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_162_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_4_176_port, QN => 
                           n_1257);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_163_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_4_177_port, QN => 
                           n_1258);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_164_port, CK => 
                           clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_4_178_port, QN => 
                           n_1259);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_165_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_4_179_port, QN => 
                           n_1260);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_166_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_4_180_port, QN => 
                           n_1261);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_167_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_4_181_port, QN => 
                           n_1262);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_168_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_182_port, QN => 
                           n_1263);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_169_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_4_183_port, QN => 
                           n_1264);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_170_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_4_184_port, QN => 
                           n_1265);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_171_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_4_185_port, QN => 
                           n_1266);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_172_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_4_186_port, QN => 
                           n_1267);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_173_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_4_187_port, QN => 
                           n_1268);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_174_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_4_188_port, QN => 
                           n_1269);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_175_port, CK => 
                           clk, RN => n11242, Q => 
                           boothmul_pipelined_i_muxes_in_4_189_port, QN => 
                           n_1270);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_176_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_4_190_port, QN => 
                           n_1271);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_20_port, CK => clk
                           , RN => n11238, Q => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, QN => 
                           n_1272);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_19_port, CK => clk
                           , RN => n11242, Q => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, QN => 
                           n_1273);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_18_port, CK => clk
                           , RN => n11231, Q => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, QN => 
                           n_1274);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_17_port, CK => clk
                           , RN => n11236, Q => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, QN => 
                           n_1275);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_16_port, CK => clk
                           , RN => n11239, Q => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, QN => 
                           n_1276);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_15_port, CK => clk
                           , RN => n11234, Q => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, QN => 
                           n_1277);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_14_port, CK => clk
                           , RN => n11238, Q => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, QN => 
                           n_1278);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_13_port, CK => clk
                           , RN => n11238, Q => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, QN => 
                           n_1279);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_12_port, CK => clk
                           , RN => n11235, Q => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, QN => 
                           n_1280);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_11_port, CK => clk
                           , RN => n11244, Q => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, QN => 
                           n_1281);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_10_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, QN => 
                           n_1282);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_9_port, CK => clk, RN
                           => n11233, Q => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, QN => n_1283
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_8_port, CK => clk, RN
                           => n11235, Q => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, QN => n_1284
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_7_port, CK => clk, RN
                           => n11233, Q => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, QN => n_1285
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_6_port, CK => clk, RN
                           => n11233, Q => n_1286, QN => n5124);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_5_port, CK => clk, RN
                           => n11244, Q => 
                           boothmul_pipelined_i_sum_out_3_5_port, QN => n_1287)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           n3091, CK => clk, RN => n11238, Q => 
                           boothmul_pipelined_i_sum_out_3_4_port, QN => n_1288)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_3_port, CK => clk, RN
                           => n11235, Q => 
                           boothmul_pipelined_i_sum_out_3_3_port, QN => n_1289)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_2_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_3_2_port, QN => n_1290)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_1_port, CK => clk, RN
                           => n11234, Q => 
                           boothmul_pipelined_i_sum_out_3_1_port, QN => n_1291)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_0_port, CK => clk, RN
                           => n11240, Q => 
                           boothmul_pipelined_i_sum_out_3_0_port, QN => n_1292)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_46_port, QN => n7164
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_3_47_port, QN => 
                           n_1293);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_3_48_port, QN => 
                           n_1294);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => n11241, Q => 
                           boothmul_pipelined_i_muxes_in_3_49_port, QN => 
                           n_1295);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => n11240, Q => 
                           boothmul_pipelined_i_muxes_in_3_50_port, QN => 
                           n_1296);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_3_51_port, QN => 
                           n_1297);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_3_52_port, QN => 
                           n_1298);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_3_53_port, QN => 
                           n_1299);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => n11233, Q => 
                           boothmul_pipelined_i_muxes_in_3_54_port, QN => 
                           n_1300);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_3_55_port, QN => 
                           n_1301);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_3_56_port, QN => 
                           n_1302);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_3_57_port, QN => 
                           n_1303);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_3_58_port, QN => 
                           n_1304);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => n11239, Q => 
                           boothmul_pipelined_i_muxes_in_3_59_port, QN => 
                           n_1305);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_3_60_port, QN => 
                           n_1306);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_119_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_3_161_port, QN => 
                           n_1307);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_3_162_port, QN => 
                           n_1308);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => n11231, Q => 
                           boothmul_pipelined_i_muxes_in_3_163_port, QN => 
                           n_1309);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => n11235, Q => 
                           boothmul_pipelined_i_muxes_in_3_164_port, QN => 
                           n_1310);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_3_165_port, QN => 
                           n_1311);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => n11234, Q => 
                           boothmul_pipelined_i_muxes_in_3_166_port, QN => 
                           n_1312);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_3_167_port, QN => 
                           n_1313);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_3_168_port, QN => 
                           n_1314);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => n11243, Q => 
                           boothmul_pipelined_i_muxes_in_3_169_port, QN => 
                           n_1315);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => n11244, Q => 
                           boothmul_pipelined_i_muxes_in_3_170_port, QN => 
                           n_1316);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_3_171_port, QN => 
                           n_1317);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_3_172_port, QN => 
                           n_1318);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_3_173_port, QN => 
                           n_1319);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => n11237, Q => 
                           boothmul_pipelined_i_muxes_in_3_174_port, QN => 
                           n_1320);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => n11238, Q => 
                           boothmul_pipelined_i_muxes_in_3_175_port, QN => 
                           n_1321);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => n11236, Q => 
                           boothmul_pipelined_i_muxes_in_3_176_port, QN => 
                           n_1322);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_18_port, CK => clk
                           , RN => n11232, Q => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, QN => 
                           n_1323);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_17_port, CK => clk
                           , RN => n11242, Q => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, QN => 
                           n_1324);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_16_port, CK => clk
                           , RN => n11235, Q => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, QN => 
                           n_1325);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_15_port, CK => clk
                           , RN => n11242, Q => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, QN => 
                           n_1326);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_14_port, CK => clk
                           , RN => n11239, Q => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, QN => 
                           n_1327);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_13_port, CK => clk
                           , RN => n11245, Q => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, QN => 
                           n_1328);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_12_port, CK => clk
                           , RN => n11239, Q => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, QN => 
                           n_1329);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_11_port, CK => clk
                           , RN => n11232, Q => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, QN => 
                           n_1330);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_10_port, CK => clk
                           , RN => n11231, Q => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, QN => 
                           n_1331);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_9_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, QN => n_1332
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_8_port, CK => clk, RN
                           => n11244, Q => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, QN => n_1333
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_7_port, CK => clk, RN
                           => n11242, Q => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, QN => n_1334
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_6_port, CK => clk, RN
                           => n11241, Q => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, QN => n_1335
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_5_port, CK => clk, RN
                           => n11233, Q => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, QN => n_1336
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_4_port, CK => clk, RN
                           => n11231, Q => n_1337, QN => n5130);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_3_port, CK => clk, RN
                           => n11232, Q => 
                           boothmul_pipelined_i_sum_out_2_3_port, QN => n_1338)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           n3086, CK => clk, RN => n11243, Q => 
                           boothmul_pipelined_i_sum_out_2_2_port, QN => n_1339)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           n2006, CK => clk, RN => n11245, Q => 
                           boothmul_pipelined_i_sum_out_2_1_port, QN => n_1340)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_0_port, CK => clk, RN
                           => n11242, Q => 
                           boothmul_pipelined_i_sum_out_2_0_port, QN => n_1341)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => n11232, Q => 
                           boothmul_pipelined_i_muxes_in_3_177_port, QN => 
                           n3077);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n13259, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n2007, B => n2008, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n2005, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n2004, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n2002, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n2000, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1998, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1993, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1990, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1988, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1986, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1984, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1982, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1980, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1978, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1976, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => n2003, 
                           CI => n3083, CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => boothmul_pipelined_i_sum_out_1_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => n2001, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_out_1_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => n1999, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_1_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => n1994, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_1_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => n1992, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_1_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => n1989, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_1_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => n1987, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_1_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => n1985, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_1_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => n1983, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_1_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => n1981, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_1_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => n1979, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_1_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => n1977, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_1_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_1_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_1_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_1_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1342, S => 
                           boothmul_pipelined_i_sum_out_1_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CI => n3085,
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_2_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_2_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_2_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_2_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_2_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_2_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_2_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_2_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_2_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_2_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_2_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_2_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_2_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_2_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_2_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CO => n_1343, S => 
                           boothmul_pipelined_i_sum_out_2_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3084,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_3_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_3_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_3_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_3_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_3_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_3_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_3_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_3_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_3_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_3_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_3_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_3_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_3_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_3_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_3_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n1991, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1344, S => 
                           boothmul_pipelined_i_sum_out_3_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CI => n3090,
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_4_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_4_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_4_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_4_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_4_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_4_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_4_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_4_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_4_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_4_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_4_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_4_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_4_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_4_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_4_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n1997, B => boothmul_pipelined_i_sum_B_in_4_24_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1345, S => 
                           boothmul_pipelined_i_sum_out_4_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CI => n3089
                           , CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_5_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_5_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_5_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_5_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_5_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_5_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_5_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_5_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_5_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_5_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_5_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_5_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_5_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_5_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_5_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n1996, B => boothmul_pipelined_i_sum_B_in_5_26_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1346, S => 
                           boothmul_pipelined_i_sum_out_5_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CI => n3088
                           , CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_6_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_6_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_6_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_6_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_6_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_6_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_6_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_6_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_6_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_6_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_6_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_6_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_6_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_out_6_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_out_6_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n1995, B => boothmul_pipelined_i_sum_B_in_6_28_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1347, S => 
                           boothmul_pipelined_i_sum_out_6_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CI => n3087
                           , CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_29_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1348, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n2009, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n2009, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n13259, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n2009, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n2009, Q => 
                           DATA2_I_26_port);
   U3 : CLKBUF_X1 port map( A => n11234, Z => n11231);
   U4 : CLKBUF_X1 port map( A => n11234, Z => n11232);
   U5 : CLKBUF_X1 port map( A => n11234, Z => n11233);
   U6 : CLKBUF_X1 port map( A => rst_BAR, Z => n11234);
   U7 : CLKBUF_X1 port map( A => n11238, Z => n11235);
   U8 : CLKBUF_X1 port map( A => n11231, Z => n11236);
   U9 : CLKBUF_X1 port map( A => n11232, Z => n11237);
   U10 : CLKBUF_X1 port map( A => n11232, Z => n11238);
   U11 : CLKBUF_X1 port map( A => n11232, Z => n11239);
   U12 : CLKBUF_X1 port map( A => n11232, Z => n11240);
   U13 : CLKBUF_X1 port map( A => n11233, Z => n11241);
   U14 : CLKBUF_X1 port map( A => n11233, Z => n11242);
   U15 : CLKBUF_X1 port map( A => n11233, Z => n11243);
   U16 : CLKBUF_X1 port map( A => n11233, Z => n11244);
   U17 : CLKBUF_X1 port map( A => n11233, Z => n11245);
   U18 : NOR2_X2 port map( A1 => n12926, A2 => n11404, ZN => n12917);
   U19 : NOR2_X4 port map( A1 => n11288, A2 => n12080, ZN => n12197);
   U20 : INV_X1 port map( A => n2009, ZN => n12927);
   U21 : CLKBUF_X1 port map( A => n12962, Z => n12952);
   U22 : INV_X1 port map( A => data1_mul_0_port, ZN => n2008);
   U23 : INV_X1 port map( A => data2_mul_1_port, ZN => n11246);
   U24 : NOR2_X1 port map( A1 => boothmul_pipelined_i_encoder_out_0_0_port, A2 
                           => n11246, ZN => n11257);
   U25 : CLKBUF_X1 port map( A => n11257, Z => n13234);
   U26 : NAND2_X1 port map( A1 => n11246, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n13237);
   U27 : INV_X1 port map( A => n13237, ZN => n11737);
   U28 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN =>
                           n12964);
   U29 : NOR2_X1 port map( A1 => n11246, A2 => n12964, ZN => n13235);
   U30 : CLKBUF_X1 port map( A => n13235, Z => n11260);
   U31 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, A2
                           => n13234, B1 => data1_mul_14_port, B2 => n11737, C1
                           => boothmul_pipelined_i_muxes_in_0_103_port, C2 => 
                           n11260, ZN => n11247);
   U32 : INV_X1 port map( A => n11247, ZN => n1977);
   U33 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, A2
                           => n13234, B1 => data1_mul_13_port, B2 => n11737, C1
                           => boothmul_pipelined_i_muxes_in_0_104_port, C2 => 
                           n13235, ZN => n11248);
   U34 : INV_X1 port map( A => n11248, ZN => n1979);
   U35 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, A2
                           => n13234, B1 => data1_mul_12_port, B2 => n11737, C1
                           => boothmul_pipelined_i_muxes_in_0_105_port, C2 => 
                           n11260, ZN => n11249);
   U36 : INV_X1 port map( A => n11249, ZN => n1981);
   U37 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, A2
                           => n13234, B1 => data1_mul_11_port, B2 => n11737, C1
                           => boothmul_pipelined_i_muxes_in_0_106_port, C2 => 
                           n13235, ZN => n11250);
   U38 : INV_X1 port map( A => n11250, ZN => n1983);
   U39 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, A2
                           => n11257, B1 => data1_mul_10_port, B2 => n11737, C1
                           => boothmul_pipelined_i_muxes_in_0_107_port, C2 => 
                           n11260, ZN => n11251);
   U40 : INV_X1 port map( A => n11251, ZN => n1985);
   U41 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, A2
                           => n11257, B1 => data1_mul_9_port, B2 => n11737, C1 
                           => boothmul_pipelined_i_muxes_in_0_108_port, C2 => 
                           n11260, ZN => n11252);
   U42 : INV_X1 port map( A => n11252, ZN => n1987);
   U43 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, A2
                           => n11257, B1 => data1_mul_8_port, B2 => n11737, C1 
                           => boothmul_pipelined_i_muxes_in_0_109_port, C2 => 
                           n11260, ZN => n11253);
   U44 : INV_X1 port map( A => n11253, ZN => n1989);
   U45 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, A2
                           => n11257, B1 => data1_mul_7_port, B2 => n11737, C1 
                           => boothmul_pipelined_i_muxes_in_0_110_port, C2 => 
                           n13235, ZN => n11254);
   U46 : INV_X1 port map( A => n11254, ZN => n1992);
   U47 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, A2
                           => n11257, B1 => data1_mul_6_port, B2 => n11737, C1 
                           => boothmul_pipelined_i_muxes_in_0_111_port, C2 => 
                           n11260, ZN => n11255);
   U48 : INV_X1 port map( A => n11255, ZN => n1994);
   U49 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, A2
                           => n11257, B1 => data1_mul_5_port, B2 => n11737, C1 
                           => boothmul_pipelined_i_muxes_in_0_112_port, C2 => 
                           n11260, ZN => n11256);
   U50 : INV_X1 port map( A => n11256, ZN => n1999);
   U51 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, A2
                           => n11257, B1 => data1_mul_4_port, B2 => n11737, C1 
                           => boothmul_pipelined_i_muxes_in_0_113_port, C2 => 
                           n13235, ZN => n11258);
   U52 : INV_X1 port map( A => n11258, ZN => n2001);
   U53 : AOI222_X1 port map( A1 => n13234, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           data1_mul_3_port, B2 => n11737, C1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, C2 => 
                           n13235, ZN => n11259);
   U54 : INV_X1 port map( A => n11259, ZN => n2003);
   U55 : AOI222_X1 port map( A1 => data1_mul_0_port, A2 => n13234, B1 => 
                           data1_mul_1_port, B2 => n11737, C1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, C2 => 
                           n11260, ZN => n11261);
   U56 : INV_X1 port map( A => n11261, ZN => n2006);
   U57 : CLKBUF_X1 port map( A => DATA1(10), Z => n13263);
   U58 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n11262);
   U59 : INV_X1 port map( A => FUNC(2), ZN => n11277);
   U60 : NAND2_X1 port map( A1 => n11262, A2 => n11277, ZN => n2009);
   U61 : CLKBUF_X1 port map( A => n2009, Z => n13259);
   U62 : CLKBUF_X1 port map( A => DATA1(2), Z => n13260);
   U63 : CLKBUF_X1 port map( A => DATA1(5), Z => n13261);
   U64 : CLKBUF_X1 port map( A => DATA1(8), Z => n13262);
   U65 : NOR3_X1 port map( A1 => FUNC(0), A2 => FUNC(1), A3 => n11277, ZN => 
                           n11276);
   U66 : INV_X1 port map( A => FUNC(3), ZN => n12926);
   U67 : NAND2_X1 port map( A1 => n11276, A2 => n12926, ZN => n553);
   U68 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n11275);
   U69 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n12556);
   U70 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => n12556
                           , ZN => n11405);
   U71 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => n11275
                           , ZN => n12588);
   U72 : NOR2_X1 port map( A1 => n11405, A2 => n12588, ZN => n11719);
   U73 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => n11273
                           );
   U74 : AND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n12634);
   U75 : INV_X1 port map( A => DATA1(8), ZN => n12696);
   U76 : XNOR2_X1 port map( A => DATA2_I_9_port, B => DATA1(9), ZN => n11820);
   U77 : INV_X1 port map( A => DATA2_I_8_port, ZN => n11263);
   U78 : NOR3_X1 port map( A1 => n12696, A2 => n11820, A3 => n11263, ZN => 
                           n12614);
   U79 : NAND2_X1 port map( A1 => n13263, A2 => DATA2_I_10_port, ZN => n11272);
   U80 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => n11272
                           , ZN => n11715);
   U81 : INV_X1 port map( A => n11715, ZN => n12633);
   U82 : OAI21_X1 port map( B1 => n12634, B2 => n12614, A => n12633, ZN => 
                           n11264);
   U83 : INV_X1 port map( A => n11264, ZN => n12613);
   U84 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => n13263, A => n12613, 
                           ZN => n12602);
   U85 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n11714);
   U86 : OAI21_X1 port map( B1 => n11273, B2 => n12602, A => n11714, ZN => 
                           n12587);
   U87 : NOR2_X1 port map( A1 => n11275, A2 => n11405, ZN => n11274);
   U88 : AOI21_X1 port map( B1 => n11719, B2 => n12587, A => n11274, ZN => 
                           n11713);
   U89 : NAND2_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, ZN => n11270)
                           ;
   U90 : OAI21_X1 port map( B1 => DATA1(7), B2 => DATA2_I_7_port, A => n11270, 
                           ZN => n11897);
   U91 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n11883)
                           ;
   U92 : NAND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n11267)
                           ;
   U93 : INV_X1 port map( A => n11267, ZN => n11881);
   U94 : XOR2_X1 port map( A => DATA2_I_3_port, B => DATA1(3), Z => n12059);
   U95 : NAND2_X1 port map( A1 => n13260, A2 => DATA2_I_2_port, ZN => n11878);
   U96 : OAI21_X1 port map( B1 => n13260, B2 => DATA2_I_2_port, A => n11878, ZN
                           => n12230);
   U97 : CLKBUF_X1 port map( A => DATA1(1), Z => n12398);
   U98 : NAND2_X1 port map( A1 => n12398, A2 => DATA2_I_1_port, ZN => n11876);
   U99 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n12639)
                           ;
   U100 : INV_X1 port map( A => n12639, ZN => n12401);
   U101 : NOR2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n12405)
                           ;
   U102 : OAI21_X1 port map( B1 => DATA1(1), B2 => DATA2_I_1_port, A => n11876,
                           ZN => n12404);
   U103 : NOR2_X1 port map( A1 => n12405, A2 => n12404, ZN => n12403);
   U104 : OAI21_X1 port map( B1 => n12401, B2 => cin, A => n12403, ZN => n11265
                           );
   U105 : OAI221_X1 port map( B1 => n12230, B2 => n11876, C1 => n12230, C2 => 
                           n11265, A => n11878, ZN => n11266);
   U106 : AND2_X1 port map( A1 => DATA1(3), A2 => DATA2_I_3_port, ZN => n11879)
                           ;
   U107 : AOI21_X1 port map( B1 => n12059, B2 => n11266, A => n11879, ZN => 
                           n11268);
   U108 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n11880
                           );
   U109 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n11880,
                           ZN => n12009);
   U110 : OAI21_X1 port map( B1 => DATA1(5), B2 => DATA2_I_5_port, A => n11267,
                           ZN => n11943);
   U111 : AOI221_X1 port map( B1 => n11268, B2 => n11880, C1 => n12009, C2 => 
                           n11880, A => n11943, ZN => n11269);
   U112 : XOR2_X1 port map( A => DATA2_I_6_port, B => DATA1(6), Z => n11885);
   U113 : OAI21_X1 port map( B1 => n11881, B2 => n11269, A => n11885, ZN => 
                           n11271);
   U114 : OAI221_X1 port map( B1 => n11897, B2 => n11883, C1 => n11897, C2 => 
                           n11271, A => n11270, ZN => n11717);
   U115 : NOR2_X1 port map( A1 => n13259, A2 => n11717, ZN => n12585);
   U116 : NAND2_X1 port map( A1 => n12927, A2 => n11717, ZN => n12533);
   U117 : INV_X1 port map( A => n12533, ZN => n12627);
   U118 : NOR2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n11818)
                           ;
   U119 : NOR2_X1 port map( A1 => n11818, A2 => n11820, ZN => n12629);
   U120 : OAI21_X1 port map( B1 => n12634, B2 => n12629, A => n12633, ZN => 
                           n12628);
   U121 : AND2_X1 port map( A1 => n11272, A2 => n12628, ZN => n12598);
   U122 : OAI21_X1 port map( B1 => n11273, B2 => n12598, A => n11714, ZN => 
                           n12579);
   U123 : AOI21_X1 port map( B1 => n11719, B2 => n12579, A => n11274, ZN => 
                           n12532);
   U124 : AOI22_X1 port map( A1 => n11713, A2 => n12585, B1 => n12627, B2 => 
                           n12532, ZN => n12557);
   U125 : AOI21_X1 port map( B1 => n11275, B2 => n11405, A => n12557, ZN => 
                           n11411);
   U126 : NAND2_X1 port map( A1 => FUNC(3), A2 => n11276, ZN => n12648);
   U127 : INV_X1 port map( A => n12648, ZN => n12520);
   U128 : INV_X1 port map( A => FUNC(0), ZN => n12737);
   U129 : NAND3_X1 port map( A1 => n11277, A2 => n12737, A3 => FUNC(1), ZN => 
                           n12641);
   U130 : INV_X1 port map( A => n12641, ZN => n12622);
   U131 : NAND2_X1 port map( A1 => n12926, A2 => n12622, ZN => n11935);
   U132 : INV_X1 port map( A => n11935, ZN => n12521);
   U133 : NOR2_X1 port map( A1 => n12520, A2 => n12521, ZN => n12616);
   U134 : INV_X1 port map( A => DATA2(13), ZN => n12946);
   U135 : INV_X1 port map( A => DATA1(13), ZN => n11803);
   U136 : NOR3_X1 port map( A1 => n12616, A2 => n12946, A3 => n11803, ZN => 
                           n11410);
   U137 : INV_X1 port map( A => DATA2(5), ZN => n12956);
   U138 : NAND4_X1 port map( A1 => n12956, A2 => n12737, A3 => FUNC(2), A4 => 
                           FUNC(1), ZN => n12159);
   U139 : INV_X1 port map( A => n12159, ZN => n11278);
   U140 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(4), ZN => n11611);
   U141 : INV_X1 port map( A => n11611, ZN => n11616);
   U142 : NAND2_X1 port map( A1 => DATA2(3), A2 => n11616, ZN => n11704);
   U143 : INV_X1 port map( A => DATA2(1), ZN => n12960);
   U144 : NOR2_X1 port map( A1 => n11704, A2 => n12960, ZN => n12911);
   U145 : NAND2_X1 port map( A1 => DATA2(0), A2 => n12911, ZN => n12160);
   U146 : NAND2_X1 port map( A1 => n11278, A2 => n12160, ZN => n11404);
   U147 : NOR2_X1 port map( A1 => FUNC(3), A2 => n11404, ZN => n12551);
   U148 : INV_X1 port map( A => n12551, ZN => n12610);
   U149 : NAND2_X1 port map( A1 => DATA2(0), A2 => DATA2(1), ZN => n11561);
   U150 : INV_X1 port map( A => n11561, ZN => n11608);
   U151 : NAND2_X1 port map( A1 => DATA2(3), A2 => n11608, ZN => n11412);
   U152 : OR2_X1 port map( A1 => DATA2(4), A2 => DATA2(5), ZN => n12135);
   U153 : NOR3_X1 port map( A1 => DATA2(2), A2 => n11412, A3 => n12135, ZN => 
                           n12570);
   U154 : INV_X1 port map( A => DATA2(3), ZN => n12958);
   U155 : INV_X1 port map( A => n12135, ZN => n12870);
   U156 : NAND2_X1 port map( A1 => n12958, A2 => n12870, ZN => n11288);
   U157 : NOR2_X1 port map( A1 => n11288, A2 => DATA2(2), ZN => n12105);
   U158 : CLKBUF_X1 port map( A => n12105, Z => n12186);
   U159 : NAND2_X1 port map( A1 => n11608, A2 => n12186, ZN => n12240);
   U160 : INV_X1 port map( A => n12240, ZN => n11853);
   U161 : CLKBUF_X1 port map( A => n11853, Z => n12018);
   U162 : NOR2_X1 port map( A1 => DATA2(0), A2 => DATA2(1), ZN => n11414);
   U163 : NAND2_X1 port map( A1 => n11414, A2 => n12105, ZN => n12220);
   U164 : INV_X1 port map( A => n12220, ZN => n12189);
   U165 : NAND2_X1 port map( A1 => n12189, A2 => DATA1(9), ZN => n11802);
   U166 : NAND2_X1 port map( A1 => DATA2(0), A2 => n12960, ZN => n11672);
   U167 : INV_X1 port map( A => n12186, ZN => n12017);
   U168 : NOR2_X1 port map( A1 => n11672, A2 => n12017, ZN => n12835);
   U169 : NAND2_X1 port map( A1 => n12835, A2 => DATA1(8), ZN => n11855);
   U170 : NOR2_X1 port map( A1 => n12960, A2 => DATA2(0), ZN => n11615);
   U171 : NAND2_X1 port map( A1 => n12105, A2 => n11615, ZN => n12241);
   U172 : INV_X1 port map( A => n12241, ZN => n12223);
   U173 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(7), ZN => n11948);
   U174 : NAND2_X1 port map( A1 => n13261, A2 => n12017, ZN => n12409);
   U175 : NAND4_X1 port map( A1 => n11802, A2 => n11855, A3 => n11948, A4 => 
                           n12409, ZN => n11279);
   U176 : AOI21_X1 port map( B1 => n12018, B2 => DATA1(6), A => n11279, ZN => 
                           n11290);
   U177 : OAI21_X1 port map( B1 => n11288, B2 => DATA2(1), A => n11752, ZN => 
                           n11954);
   U178 : CLKBUF_X1 port map( A => n12835, Z => n12408);
   U179 : INV_X1 port map( A => DATA1(7), ZN => n12693);
   U180 : NOR2_X1 port map( A1 => n12105, A2 => n12693, ZN => n11281);
   U181 : INV_X1 port map( A => DATA1(11), ZN => n12595);
   U182 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(9), ZN => n11856);
   U183 : NAND2_X1 port map( A1 => n11853, A2 => n13262, ZN => n11949);
   U184 : OAI211_X1 port map( C1 => n12220, C2 => n12595, A => n11856, B => 
                           n11949, ZN => n11280);
   U185 : AOI211_X1 port map( C1 => DATA1(10), C2 => n12408, A => n11281, B => 
                           n11280, ZN => n11299);
   U186 : INV_X1 port map( A => DATA2(0), ZN => n12961);
   U187 : INV_X1 port map( A => DATA2(2), ZN => n12959);
   U188 : OAI21_X1 port map( B1 => n12961, B2 => n12959, A => n11954, ZN => 
                           n12113);
   U189 : AOI22_X1 port map( A1 => n13263, A2 => n12189, B1 => DATA1(6), B2 => 
                           n12017, ZN => n11283);
   U190 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(9), ZN => n11282);
   U191 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(8), ZN => n11904);
   U192 : NAND2_X1 port map( A1 => n11853, A2 => DATA1(7), ZN => n11977);
   U193 : AND4_X1 port map( A1 => n11283, A2 => n11282, A3 => n11904, A4 => 
                           n11977, ZN => n11287);
   U194 : OR3_X1 port map( A1 => n12959, A2 => n11672, A3 => n11288, ZN => 
                           n12111);
   U195 : OAI222_X1 port map( A1 => n11290, A2 => n11954, B1 => n11299, B2 => 
                           n12113, C1 => n11287, C2 => n12111, ZN => n11574);
   U196 : INV_X1 port map( A => n11574, ZN => n11578);
   U197 : CLKBUF_X1 port map( A => n11954, Z => n12109);
   U198 : INV_X1 port map( A => n12109, ZN => n12192);
   U199 : OAI21_X1 port map( B1 => DATA2(0), B2 => n11288, A => n12192, ZN => 
                           n12080);
   U200 : INV_X1 port map( A => n12197, ZN => n12416);
   U201 : CLKBUF_X1 port map( A => n12416, Z => n12850);
   U202 : INV_X1 port map( A => n12135, ZN => n12034);
   U203 : INV_X1 port map( A => n11414, ZN => n11703);
   U204 : NOR2_X1 port map( A1 => n11703, A2 => DATA2(2), ZN => n11413);
   U205 : AND3_X1 port map( A1 => DATA2(3), A2 => n12034, A3 => n11413, ZN => 
                           n12117);
   U206 : CLKBUF_X1 port map( A => n12113, Z => n12002);
   U207 : INV_X1 port map( A => DATA1(6), ZN => n12691);
   U208 : NOR2_X1 port map( A1 => n12241, A2 => n12691, ZN => n11980);
   U209 : NAND2_X1 port map( A1 => n12189, A2 => n13262, ZN => n11827);
   U210 : NAND2_X1 port map( A1 => n12835, A2 => DATA1(7), ZN => n11903);
   U211 : NAND2_X1 port map( A1 => n11853, A2 => DATA1(5), ZN => n12185);
   U212 : NAND2_X1 port map( A1 => DATA1(4), A2 => n11752, ZN => n12836);
   U213 : NAND4_X1 port map( A1 => n11827, A2 => n11903, A3 => n12185, A4 => 
                           n12836, ZN => n11284);
   U214 : NOR2_X1 port map( A1 => n11980, A2 => n11284, ZN => n11292);
   U215 : OAI222_X1 port map( A1 => n12002, A2 => n11287, B1 => n12111, B2 => 
                           n11290, C1 => n12109, C2 => n11292, ZN => n11572);
   U216 : CLKBUF_X1 port map( A => n12080, Z => n12115);
   U217 : INV_X1 port map( A => n12835, ZN => n12396);
   U218 : NOR2_X1 port map( A1 => n12396, A2 => n12595, ZN => n11786);
   U219 : INV_X1 port map( A => DATA1(10), ZN => n12651);
   U220 : NOR2_X1 port map( A1 => n12241, A2 => n12651, ZN => n11829);
   U221 : NOR2_X1 port map( A1 => n12105, A2 => n12696, ZN => n11286);
   U222 : INV_X1 port map( A => DATA1(12), ZN => n12772);
   U223 : INV_X1 port map( A => DATA1(9), ZN => n11950);
   U224 : OAI22_X1 port map( A1 => n12772, A2 => n12220, B1 => n12240, B2 => 
                           n11950, ZN => n11285);
   U225 : NOR4_X1 port map( A1 => n11786, A2 => n11829, A3 => n11286, A4 => 
                           n11285, ZN => n11298);
   U226 : OAI222_X1 port map( A1 => n11287, A2 => n12109, B1 => n11298, B2 => 
                           n12113, C1 => n11299, C2 => n12111, ZN => n11573);
   U227 : AOI22_X1 port map( A1 => n12117, A2 => n11572, B1 => n12115, B2 => 
                           n11573, ZN => n11294);
   U228 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(2), ZN => n11312);
   U229 : OAI211_X1 port map( C1 => n12960, C2 => n12958, A => n11312, B => 
                           n12870, ZN => n12119);
   U230 : CLKBUF_X1 port map( A => n12119, Z => n12030);
   U231 : INV_X1 port map( A => n12030, ZN => n12853);
   U232 : NAND3_X1 port map( A1 => n11703, A2 => n11288, A3 => n12853, ZN => 
                           n12359);
   U233 : INV_X1 port map( A => n12359, ZN => n12857);
   U234 : NOR2_X1 port map( A1 => n12396, A2 => n12691, ZN => n11952);
   U235 : INV_X1 port map( A => DATA1(5), ZN => n12652);
   U236 : NOR2_X1 port map( A1 => n12241, A2 => n12652, ZN => n12019);
   U237 : INV_X1 port map( A => DATA1(3), ZN => n11306);
   U238 : NAND2_X1 port map( A1 => n11853, A2 => DATA1(4), ZN => n12410);
   U239 : CLKBUF_X1 port map( A => n12189, Z => n12834);
   U240 : NAND2_X1 port map( A1 => n12834, A2 => DATA1(7), ZN => n11854);
   U241 : OAI211_X1 port map( C1 => n12105, C2 => n11306, A => n12410, B => 
                           n11854, ZN => n11289);
   U242 : NOR3_X1 port map( A1 => n11952, A2 => n12019, A3 => n11289, ZN => 
                           n11305);
   U243 : OAI222_X1 port map( A1 => n12002, A2 => n11290, B1 => n12111, B2 => 
                           n11292, C1 => n11954, C2 => n11305, ZN => n11746);
   U244 : INV_X1 port map( A => DATA1(4), ZN => n12001);
   U245 : NOR2_X1 port map( A1 => n12241, A2 => n12001, ZN => n12188);
   U246 : INV_X1 port map( A => DATA1(2), ZN => n12224);
   U247 : NAND2_X1 port map( A1 => n11853, A2 => DATA1(3), ZN => n12837);
   U248 : NAND2_X1 port map( A1 => n12834, A2 => DATA1(6), ZN => n11902);
   U249 : OAI211_X1 port map( C1 => n12186, C2 => n12224, A => n12837, B => 
                           n11902, ZN => n11291);
   U250 : AOI211_X1 port map( C1 => DATA1(5), C2 => n12408, A => n12188, B => 
                           n11291, ZN => n11308);
   U251 : OAI222_X1 port map( A1 => n12002, A2 => n11292, B1 => n12111, B2 => 
                           n11305, C1 => n11954, C2 => n11308, ZN => n11843);
   U252 : AOI22_X1 port map( A1 => n12857, A2 => n11746, B1 => n12119, B2 => 
                           n11843, ZN => n11293);
   U253 : OAI211_X1 port map( C1 => n11578, C2 => n12850, A => n11294, B => 
                           n11293, ZN => n12568);
   U254 : AND3_X1 port map( A1 => n12034, A2 => n11412, A3 => n11312, ZN => 
                           n12617);
   U255 : INV_X1 port map( A => n11573, ZN => n11583);
   U256 : INV_X1 port map( A => n11572, ZN => n11295);
   U257 : CLKBUF_X1 port map( A => n12359, Z => n12026);
   U258 : OAI22_X1 port map( A1 => n11583, A2 => n12850, B1 => n11295, B2 => 
                           n12026, ZN => n11302);
   U259 : INV_X1 port map( A => n12115, ZN => n12415);
   U260 : INV_X1 port map( A => n12002, ZN => n12842);
   U261 : NOR2_X1 port map( A1 => n12241, A2 => n12595, ZN => n11805);
   U262 : NOR2_X1 port map( A1 => n12396, A2 => n12772, ZN => n11768);
   U263 : AOI211_X1 port map( C1 => DATA1(9), C2 => n11752, A => n11805, B => 
                           n11768, ZN => n11297);
   U264 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12189, ZN => n11296);
   U265 : OAI211_X1 port map( C1 => n12651, C2 => n12240, A => n11297, B => 
                           n11296, ZN => n11498);
   U266 : INV_X1 port map( A => n12111, ZN => n12193);
   U267 : INV_X1 port map( A => n11298, ZN => n11497);
   U268 : INV_X1 port map( A => n11299, ZN => n11300);
   U269 : AOI222_X1 port map( A1 => n12842, A2 => n11498, B1 => n12193, B2 => 
                           n11497, C1 => n12192, C2 => n11300, ZN => n11584);
   U270 : INV_X1 port map( A => n12117, ZN => n12361);
   U271 : OAI22_X1 port map( A1 => n12415, A2 => n11584, B1 => n11578, B2 => 
                           n12361, ZN => n11301);
   U272 : AOI211_X1 port map( C1 => n12030, C2 => n11746, A => n11302, B => 
                           n11301, ZN => n11692);
   U273 : INV_X1 port map( A => n11692, ZN => n11675);
   U274 : AOI22_X1 port map( A1 => n12570, A2 => n12568, B1 => n12617, B2 => 
                           n11675, ZN => n11325);
   U275 : OAI21_X1 port map( B1 => n12960, B2 => n11312, A => n12870, ZN => 
                           n12128);
   U276 : CLKBUF_X1 port map( A => n12128, Z => n11960);
   U277 : NOR3_X1 port map( A1 => n12961, A2 => n11312, A3 => n11960, ZN => 
                           n12425);
   U278 : INV_X1 port map( A => n11843, ZN => n11311);
   U279 : AOI22_X1 port map( A1 => n12197, A2 => n11746, B1 => n12080, B2 => 
                           n11572, ZN => n11310);
   U280 : NOR2_X1 port map( A1 => n12220, A2 => n12652, ZN => n11304);
   U281 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(4), ZN => n12020);
   U282 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(3), ZN => n12411);
   U283 : OAI211_X1 port map( C1 => n12240, C2 => n12224, A => n12020, B => 
                           n12411, ZN => n11303);
   U284 : AOI211_X1 port map( C1 => n12398, C2 => n11752, A => n11304, B => 
                           n11303, ZN => n11936);
   U285 : OAI222_X1 port map( A1 => n12113, A2 => n11305, B1 => n12111, B2 => 
                           n11308, C1 => n12109, C2 => n11936, ZN => n11890);
   U286 : NOR2_X1 port map( A1 => n12396, A2 => n11306, ZN => n12183);
   U287 : INV_X1 port map( A => DATA1(0), ZN => n12640);
   U288 : NAND2_X1 port map( A1 => n12223, A2 => n13260, ZN => n12838);
   U289 : NAND2_X1 port map( A1 => n12834, A2 => DATA1(4), ZN => n11978);
   U290 : OAI211_X1 port map( C1 => n12186, C2 => n12640, A => n12838, B => 
                           n11978, ZN => n11307);
   U291 : AOI211_X1 port map( C1 => n12018, C2 => DATA1(1), A => n12183, B => 
                           n11307, ZN => n12003);
   U292 : OAI222_X1 port map( A1 => n12002, A2 => n11308, B1 => n12111, B2 => 
                           n11936, C1 => n11954, C2 => n12003, ZN => n11926);
   U293 : AOI22_X1 port map( A1 => n12857, A2 => n11890, B1 => n12119, B2 => 
                           n11926, ZN => n11309);
   U294 : OAI211_X1 port map( C1 => n11311, C2 => n12361, A => n11310, B => 
                           n11309, ZN => n12619);
   U295 : NOR3_X1 port map( A1 => n12135, A2 => n11703, A3 => n11312, ZN => 
                           n12126);
   U296 : CLKBUF_X1 port map( A => n12126, Z => n12569);
   U297 : INV_X1 port map( A => n12115, ZN => n12849);
   U298 : AOI22_X1 port map( A1 => n12117, A2 => n11746, B1 => n12197, B2 => 
                           n11572, ZN => n11314);
   U299 : AOI22_X1 port map( A1 => n12857, A2 => n11843, B1 => n12119, B2 => 
                           n11890, ZN => n11313);
   U300 : OAI211_X1 port map( C1 => n12849, C2 => n11578, A => n11314, B => 
                           n11313, ZN => n12593);
   U301 : AOI22_X1 port map( A1 => n12425, A2 => n12619, B1 => n12569, B2 => 
                           n12593, ZN => n11324);
   U302 : NOR4_X1 port map( A1 => DATA2(8), A2 => DATA2(9), A3 => DATA2(6), A4 
                           => DATA2(7), ZN => n11322);
   U303 : INV_X1 port map( A => DATA2(12), ZN => n12947);
   U304 : INV_X1 port map( A => DATA2(10), ZN => n12949);
   U305 : INV_X1 port map( A => DATA2(11), ZN => n12948);
   U306 : NAND4_X1 port map( A1 => n12947, A2 => n12949, A3 => n12948, A4 => 
                           n12946, ZN => n11315);
   U307 : NOR4_X1 port map( A1 => DATA2(15), A2 => DATA2(14), A3 => n12220, A4 
                           => n11315, ZN => n11321);
   U308 : NOR4_X1 port map( A1 => DATA1(12), A2 => DATA1(13), A3 => DATA1(11), 
                           A4 => DATA1(14), ZN => n11319);
   U309 : NOR4_X1 port map( A1 => DATA1(15), A2 => n13263, A3 => DATA1(9), A4 
                           => n13262, ZN => n11318);
   U310 : NOR4_X1 port map( A1 => DATA1(7), A2 => DATA1(6), A3 => n13261, A4 =>
                           DATA1(4), ZN => n11317);
   U311 : NOR4_X1 port map( A1 => DATA1(3), A2 => n13260, A3 => n12398, A4 => 
                           DATA1(0), ZN => n11316);
   U312 : AND4_X1 port map( A1 => n11319, A2 => n11318, A3 => n11317, A4 => 
                           n11316, ZN => n11320);
   U313 : AOI211_X1 port map( C1 => n11322, C2 => n11321, A => n11320, B => 
                           n553, ZN => n12508);
   U314 : INV_X1 port map( A => n12508, ZN => n12546);
   U315 : INV_X1 port map( A => n12546, ZN => n12615);
   U316 : NOR2_X1 port map( A1 => n12946, A2 => DATA1(13), ZN => n12773);
   U317 : NOR2_X1 port map( A1 => n11803, A2 => DATA2(13), ZN => n12777);
   U318 : OR2_X1 port map( A1 => n12773, A2 => n12777, ZN => n12664);
   U319 : AOI22_X1 port map( A1 => dataout_mul_13_port, A2 => n12615, B1 => 
                           n12622, B2 => n12664, ZN => n11323);
   U320 : OAI221_X1 port map( B1 => n12610, B2 => n11325, C1 => n12610, C2 => 
                           n11324, A => n11323, ZN => n11409);
   U321 : OAI21_X1 port map( B1 => n12959, B2 => n11412, A => n12870, ZN => 
                           n12873);
   U322 : INV_X1 port map( A => n12873, ZN => n12550);
   U323 : NOR2_X1 port map( A1 => n12135, A2 => n12550, ZN => n12526);
   U324 : INV_X1 port map( A => n12526, ZN => n12875);
   U325 : CLKBUF_X1 port map( A => DATA1(25), Z => n12295);
   U326 : INV_X1 port map( A => n12105, ZN => n11752);
   U327 : AOI22_X1 port map( A1 => DATA1(24), A2 => n11853, B1 => n12295, B2 =>
                           n11752, ZN => n11326);
   U328 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(23), ZN => n11511);
   U329 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(22), ZN => n11463);
   U330 : NAND2_X1 port map( A1 => n12189, A2 => DATA1(21), ZN => n11420);
   U331 : NAND4_X1 port map( A1 => n11326, A2 => n11511, A3 => n11463, A4 => 
                           n11420, ZN => n11336);
   U332 : AOI22_X1 port map( A1 => DATA1(22), A2 => n11853, B1 => DATA1(23), B2
                           => n12017, ZN => n11327);
   U333 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(21), ZN => n11464);
   U334 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(20), ZN => n11421);
   U335 : NAND2_X1 port map( A1 => n12834, A2 => DATA1(19), ZN => n11416);
   U336 : NAND4_X1 port map( A1 => n11327, A2 => n11464, A3 => n11421, A4 => 
                           n11416, ZN => n11341);
   U337 : INV_X1 port map( A => n12002, ZN => n12267);
   U338 : CLKBUF_X1 port map( A => DATA1(24), Z => n12740);
   U339 : AOI22_X1 port map( A1 => DATA1(23), A2 => n11853, B1 => n12740, B2 =>
                           n11752, ZN => n11328);
   U340 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(22), ZN => n11483);
   U341 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(21), ZN => n11442);
   U342 : NAND2_X1 port map( A1 => n12834, A2 => DATA1(20), ZN => n11427);
   U343 : NAND4_X1 port map( A1 => n11328, A2 => n11483, A3 => n11442, A4 => 
                           n11427, ZN => n11334);
   U344 : INV_X1 port map( A => n12111, ZN => n12840);
   U345 : AOI222_X1 port map( A1 => n11336, A2 => n12192, B1 => n11341, B2 => 
                           n12267, C1 => n11334, C2 => n12840, ZN => n11357);
   U346 : INV_X1 port map( A => n11357, ZN => n11377);
   U347 : AOI22_X1 port map( A1 => DATA1(24), A2 => n12834, B1 => DATA1(28), B2
                           => n11752, ZN => n11329);
   U348 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(26), ZN => n11540);
   U349 : NAND2_X1 port map( A1 => n12018, A2 => DATA1(27), ZN => n12075);
   U350 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(25), ZN => n11506);
   U351 : NAND4_X1 port map( A1 => n11329, A2 => n11540, A3 => n12075, A4 => 
                           n11506, ZN => n11383);
   U352 : INV_X1 port map( A => n12109, ZN => n12844);
   U353 : AOI22_X1 port map( A1 => n12295, A2 => n12018, B1 => DATA1(26), B2 =>
                           n11752, ZN => n11330);
   U354 : NAND2_X1 port map( A1 => n12223, A2 => n12740, ZN => n11507);
   U355 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(23), ZN => n11482);
   U356 : NAND2_X1 port map( A1 => n12189, A2 => DATA1(22), ZN => n11441);
   U357 : NAND4_X1 port map( A1 => n11330, A2 => n11507, A3 => n11482, A4 => 
                           n11441, ZN => n11335);
   U358 : AOI22_X1 port map( A1 => DATA1(23), A2 => n12189, B1 => DATA1(27), B2
                           => n11752, ZN => n11331);
   U359 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(25), ZN => n11528);
   U360 : NAND2_X1 port map( A1 => n12408, A2 => n12740, ZN => n11510);
   U361 : NAND2_X1 port map( A1 => n12018, A2 => DATA1(26), ZN => n11642);
   U362 : NAND4_X1 port map( A1 => n11331, A2 => n11528, A3 => n11510, A4 => 
                           n11642, ZN => n11374);
   U363 : AOI222_X1 port map( A1 => n11383, A2 => n12844, B1 => n11335, B2 => 
                           n12267, C1 => n11374, C2 => n12840, ZN => n12358);
   U364 : AOI222_X1 port map( A1 => n11335, A2 => n12192, B1 => n11334, B2 => 
                           n12267, C1 => n11336, C2 => n12840, ZN => n11384);
   U365 : INV_X1 port map( A => n12117, ZN => n12846);
   U366 : OAI22_X1 port map( A1 => n12853, A2 => n12358, B1 => n11384, B2 => 
                           n12846, ZN => n11338);
   U367 : INV_X1 port map( A => DATA1(19), ZN => n12459);
   U368 : NOR2_X1 port map( A1 => n12396, A2 => n12459, ZN => n11426);
   U369 : INV_X1 port map( A => DATA1(22), ZN => n12801);
   U370 : NAND2_X1 port map( A1 => n11853, A2 => DATA1(21), ZN => n11484);
   U371 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(20), ZN => n11443);
   U372 : OAI211_X1 port map( C1 => n12186, C2 => n12801, A => n11484, B => 
                           n11443, ZN => n11332);
   U373 : AOI211_X1 port map( C1 => DATA1(18), C2 => n12834, A => n11426, B => 
                           n11332, ZN => n11333);
   U374 : INV_X1 port map( A => n11333, ZN => n11344);
   U375 : AOI222_X1 port map( A1 => n11334, A2 => n12192, B1 => n11344, B2 => 
                           n12267, C1 => n11341, C2 => n12840, ZN => n11358);
   U376 : AOI222_X1 port map( A1 => n11374, A2 => n12844, B1 => n11336, B2 => 
                           n12267, C1 => n11335, C2 => n12840, ZN => n11393);
   U377 : OAI22_X1 port map( A1 => n12415, A2 => n11358, B1 => n11393, B2 => 
                           n12359, ZN => n11337);
   U378 : AOI211_X1 port map( C1 => n12197, C2 => n11377, A => n11338, B => 
                           n11337, ZN => n12472);
   U379 : INV_X1 port map( A => n12472, ZN => n11390);
   U380 : INV_X1 port map( A => n12126, ZN => n12860);
   U381 : INV_X1 port map( A => DATA1(18), ZN => n12469);
   U382 : NOR2_X1 port map( A1 => n12396, A2 => n12469, ZN => n11415);
   U383 : INV_X1 port map( A => DATA1(21), ZN => n12369);
   U384 : NAND2_X1 port map( A1 => n11853, A2 => DATA1(20), ZN => n11465);
   U385 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(19), ZN => n11422);
   U386 : OAI211_X1 port map( C1 => n12186, C2 => n12369, A => n11465, B => 
                           n11422, ZN => n11339);
   U387 : AOI211_X1 port map( C1 => DATA1(17), C2 => n12189, A => n11415, B => 
                           n11339, ZN => n11340);
   U388 : INV_X1 port map( A => n11340, ZN => n11350);
   U389 : AOI222_X1 port map( A1 => n11341, A2 => n12192, B1 => n11350, B2 => 
                           n12842, C1 => n11344, C2 => n12840, ZN => n11367);
   U390 : INV_X1 port map( A => n11367, ZN => n11361);
   U391 : NOR2_X1 port map( A1 => n12240, A2 => n12459, ZN => n11445);
   U392 : INV_X1 port map( A => DATA1(20), ZN => n12388);
   U393 : NAND2_X1 port map( A1 => n12189, A2 => DATA1(16), ZN => n11437);
   U394 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(18), ZN => n11428);
   U395 : OAI211_X1 port map( C1 => n12186, C2 => n12388, A => n11437, B => 
                           n11428, ZN => n11342);
   U396 : AOI211_X1 port map( C1 => DATA1(17), C2 => n12408, A => n11445, B => 
                           n11342, ZN => n11343);
   U397 : INV_X1 port map( A => n11343, ZN => n11351);
   U398 : AOI222_X1 port map( A1 => n12842, A2 => n11351, B1 => n12193, B2 => 
                           n11350, C1 => n12192, C2 => n11344, ZN => n11364);
   U399 : OAI22_X1 port map( A1 => n12853, A2 => n11384, B1 => n12849, B2 => 
                           n11364, ZN => n11346);
   U400 : OAI22_X1 port map( A1 => n11358, A2 => n12361, B1 => n11357, B2 => 
                           n12359, ZN => n11345);
   U401 : AOI211_X1 port map( C1 => n12197, C2 => n11361, A => n11346, B => 
                           n11345, ZN => n11751);
   U402 : INV_X1 port map( A => n12617, ZN => n12858);
   U403 : AOI22_X1 port map( A1 => DATA1(14), A2 => n12189, B1 => DATA1(18), B2
                           => n11752, ZN => n11348);
   U404 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(16), ZN => n11430);
   U405 : NAND2_X1 port map( A1 => n12835, A2 => DATA1(15), ZN => n11438);
   U406 : INV_X1 port map( A => DATA1(17), ZN => n12491);
   U407 : NOR2_X1 port map( A1 => n12240, A2 => n12491, ZN => n11425);
   U408 : INV_X1 port map( A => n11425, ZN => n11347);
   U409 : NAND4_X1 port map( A1 => n11348, A2 => n11430, A3 => n11438, A4 => 
                           n11347, ZN => n11757);
   U410 : AOI22_X1 port map( A1 => DATA1(17), A2 => n12223, B1 => DATA1(19), B2
                           => n11752, ZN => n11349);
   U411 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(16), ZN => n11433);
   U412 : NAND2_X1 port map( A1 => n12834, A2 => DATA1(15), ZN => n11452);
   U413 : NAND2_X1 port map( A1 => n11853, A2 => DATA1(18), ZN => n11423);
   U414 : NAND4_X1 port map( A1 => n11349, A2 => n11433, A3 => n11452, A4 => 
                           n11423, ZN => n11366);
   U415 : AOI222_X1 port map( A1 => n11351, A2 => n12192, B1 => n11757, B2 => 
                           n12267, C1 => n11366, C2 => n12840, ZN => n11789);
   U416 : AOI222_X1 port map( A1 => n12842, A2 => n11366, B1 => n12840, B2 => 
                           n11351, C1 => n12192, C2 => n11350, ZN => n11764);
   U417 : OAI22_X1 port map( A1 => n12849, A2 => n11789, B1 => n11764, B2 => 
                           n12416, ZN => n11353);
   U418 : OAI22_X1 port map( A1 => n12853, A2 => n11358, B1 => n11364, B2 => 
                           n12846, ZN => n11352);
   U419 : AOI211_X1 port map( C1 => n12857, C2 => n11361, A => n11353, B => 
                           n11352, ZN => n11782);
   U420 : OAI22_X1 port map( A1 => n12860, A2 => n11751, B1 => n12858, B2 => 
                           n11782, ZN => n11363);
   U421 : INV_X1 port map( A => n12570, ZN => n12862);
   U422 : INV_X1 port map( A => n11358, ZN => n11356);
   U423 : OAI22_X1 port map( A1 => n11364, A2 => n12416, B1 => n11367, B2 => 
                           n12846, ZN => n11355);
   U424 : OAI22_X1 port map( A1 => n12853, A2 => n11357, B1 => n12849, B2 => 
                           n11764, ZN => n11354);
   U425 : AOI211_X1 port map( C1 => n12857, C2 => n11356, A => n11355, B => 
                           n11354, ZN => n11774);
   U426 : CLKBUF_X1 port map( A => n12425, Z => n12869);
   U427 : INV_X1 port map( A => n12869, ZN => n12473);
   U428 : OAI22_X1 port map( A1 => n12853, A2 => n11393, B1 => n11384, B2 => 
                           n12026, ZN => n11360);
   U429 : OAI22_X1 port map( A1 => n11358, A2 => n12416, B1 => n11357, B2 => 
                           n12846, ZN => n11359);
   U430 : AOI211_X1 port map( C1 => n12080, C2 => n11361, A => n11360, B => 
                           n11359, ZN => n11399);
   U431 : OAI22_X1 port map( A1 => n12862, A2 => n11774, B1 => n12473, B2 => 
                           n11399, ZN => n11362);
   U432 : AOI211_X1 port map( C1 => n12128, C2 => n11390, A => n11363, B => 
                           n11362, ZN => n11779);
   U433 : INV_X1 port map( A => n12550, ZN => n12506);
   U434 : INV_X1 port map( A => n12128, ZN => n12865);
   U435 : OAI22_X1 port map( A1 => n12865, A2 => n11399, B1 => n11751, B2 => 
                           n12473, ZN => n11371);
   U436 : INV_X1 port map( A => n11364, ZN => n11760);
   U437 : AOI22_X1 port map( A1 => n12189, A2 => DATA1(13), B1 => DATA1(17), B2
                           => n11752, ZN => n11365);
   U438 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(15), ZN => n11434);
   U439 : NAND2_X1 port map( A1 => n12018, A2 => DATA1(16), ZN => n11417);
   U440 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(14), ZN => n11453);
   U441 : NAND4_X1 port map( A1 => n11365, A2 => n11434, A3 => n11417, A4 => 
                           n11453, ZN => n11769);
   U442 : AOI222_X1 port map( A1 => n11366, A2 => n12192, B1 => n11769, B2 => 
                           n12267, C1 => n11757, C2 => n12840, ZN => n11807);
   U443 : OAI22_X1 port map( A1 => n12849, A2 => n11807, B1 => n11764, B2 => 
                           n12846, ZN => n11369);
   U444 : OAI22_X1 port map( A1 => n12853, A2 => n11367, B1 => n11789, B2 => 
                           n12416, ZN => n11368);
   U445 : AOI211_X1 port map( C1 => n12857, C2 => n11760, A => n11369, B => 
                           n11368, ZN => n11810);
   U446 : INV_X1 port map( A => n12617, ZN => n12471);
   U447 : OAI22_X1 port map( A1 => n11810, A2 => n12471, B1 => n11782, B2 => 
                           n12862, ZN => n11370);
   U448 : NOR2_X1 port map( A1 => n11371, A2 => n11370, ZN => n11777);
   U449 : OAI21_X1 port map( B1 => n11774, B2 => n12860, A => n11777, ZN => 
                           n11372);
   U450 : INV_X1 port map( A => n11372, ZN => n11778);
   U451 : AOI22_X1 port map( A1 => DATA1(25), A2 => n12834, B1 => DATA1(29), B2
                           => n12017, ZN => n11373);
   U452 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(26), ZN => n11527);
   U453 : NAND2_X1 port map( A1 => n12018, A2 => DATA1(28), ZN => n12103);
   U454 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(27), ZN => n11641);
   U455 : NAND4_X1 port map( A1 => n11373, A2 => n11527, A3 => n12103, A4 => 
                           n11641, ZN => n11395);
   U456 : AOI222_X1 port map( A1 => n11395, A2 => n12844, B1 => n11374, B2 => 
                           n12267, C1 => n11383, C2 => n12840, ZN => n12357);
   U457 : OAI22_X1 port map( A1 => n12853, A2 => n12357, B1 => n11393, B2 => 
                           n12846, ZN => n11376);
   U458 : OAI22_X1 port map( A1 => n11384, A2 => n12416, B1 => n12358, B2 => 
                           n12026, ZN => n11375);
   U459 : AOI211_X1 port map( C1 => n12115, C2 => n11377, A => n11376, B => 
                           n11375, ZN => n12470);
   U460 : OAI22_X1 port map( A1 => n12865, A2 => n12470, B1 => n12472, B2 => 
                           n12473, ZN => n11379);
   U461 : OAI22_X1 port map( A1 => n11774, A2 => n12471, B1 => n11751, B2 => 
                           n12862, ZN => n11378);
   U462 : NOR2_X1 port map( A1 => n11379, A2 => n11378, ZN => n11391);
   U463 : OAI222_X1 port map( A1 => n12875, A2 => n11779, B1 => n12506, B2 => 
                           n11778, C1 => n11391, C2 => n12034, ZN => n12575);
   U464 : INV_X1 port map( A => n11413, ZN => n11380);
   U465 : OAI21_X1 port map( B1 => n11380, B2 => DATA2(3), A => n12135, ZN => 
                           n12877);
   U466 : CLKBUF_X1 port map( A => n12877, Z => n12541);
   U467 : INV_X1 port map( A => DATA1(28), ZN => n12244);
   U468 : NOR2_X1 port map( A1 => n12241, A2 => n12244, ZN => n12074);
   U469 : INV_X1 port map( A => DATA1(30), ZN => n12825);
   U470 : NAND2_X1 port map( A1 => n12189, A2 => DATA1(26), ZN => n11505);
   U471 : NAND2_X1 port map( A1 => n12835, A2 => DATA1(27), ZN => n11539);
   U472 : OAI211_X1 port map( C1 => n12186, C2 => n12825, A => n11505, B => 
                           n11539, ZN => n11381);
   U473 : AOI211_X1 port map( C1 => DATA1(29), C2 => n12018, A => n12074, B => 
                           n11381, ZN => n11382);
   U474 : INV_X1 port map( A => n11382, ZN => n12282);
   U475 : AOI222_X1 port map( A1 => n12842, A2 => n11383, B1 => n12840, B2 => 
                           n11395, C1 => n12844, C2 => n12282, ZN => n12362);
   U476 : INV_X1 port map( A => n12362, ZN => n11387);
   U477 : OAI22_X1 port map( A1 => n12358, A2 => n12361, B1 => n12357, B2 => 
                           n12026, ZN => n11386);
   U478 : OAI22_X1 port map( A1 => n12849, A2 => n11384, B1 => n11393, B2 => 
                           n12850, ZN => n11385);
   U479 : AOI211_X1 port map( C1 => n12030, C2 => n11387, A => n11386, B => 
                           n11385, ZN => n12475);
   U480 : OAI22_X1 port map( A1 => n12865, A2 => n12475, B1 => n11399, B2 => 
                           n12862, ZN => n11389);
   U481 : OAI22_X1 port map( A1 => n11751, A2 => n12471, B1 => n12470, B2 => 
                           n12473, ZN => n11388);
   U482 : AOI211_X1 port map( C1 => n12569, C2 => n11390, A => n11389, B => 
                           n11388, ZN => n12507);
   U483 : OAI21_X1 port map( B1 => n12860, B2 => n11399, A => n11391, ZN => 
                           n11392);
   U484 : INV_X1 port map( A => n11392, ZN => n11403);
   U485 : INV_X1 port map( A => n12470, ZN => n11402);
   U486 : INV_X1 port map( A => n11393, ZN => n11398);
   U487 : OAI22_X1 port map( A1 => n12357, A2 => n12846, B1 => n12362, B2 => 
                           n12026, ZN => n11397);
   U488 : AOI22_X1 port map( A1 => DATA1(30), A2 => n11853, B1 => DATA1(31), B2
                           => n12017, ZN => n11394);
   U489 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(29), ZN => n12104);
   U490 : NAND2_X1 port map( A1 => n12835, A2 => DATA1(28), ZN => n11640);
   U491 : NAND2_X1 port map( A1 => n12189, A2 => DATA1(27), ZN => n11526);
   U492 : NAND4_X1 port map( A1 => n11394, A2 => n12104, A3 => n11640, A4 => 
                           n11526, ZN => n12281);
   U493 : AOI222_X1 port map( A1 => n12281, A2 => n12844, B1 => n11395, B2 => 
                           n12267, C1 => n12282, C2 => n12840, ZN => n12360);
   U494 : OAI22_X1 port map( A1 => n12853, A2 => n12360, B1 => n12358, B2 => 
                           n12850, ZN => n11396);
   U495 : AOI211_X1 port map( C1 => n12115, C2 => n11398, A => n11397, B => 
                           n11396, ZN => n12474);
   U496 : OAI22_X1 port map( A1 => n12865, A2 => n12474, B1 => n12472, B2 => 
                           n12862, ZN => n11401);
   U497 : OAI22_X1 port map( A1 => n11399, A2 => n12471, B1 => n12475, B2 => 
                           n12473, ZN => n11400);
   U498 : AOI211_X1 port map( C1 => n12569, C2 => n11402, A => n11401, B => 
                           n11400, ZN => n12505);
   U499 : OAI222_X1 port map( A1 => n12875, A2 => n12507, B1 => n12873, B2 => 
                           n11403, C1 => n12505, C2 => n12870, ZN => n12572);
   U500 : NOR2_X1 port map( A1 => n12958, A2 => n12870, ZN => n12829);
   U501 : NOR2_X1 port map( A1 => n11616, A2 => n12829, ZN => n12141);
   U502 : NAND3_X1 port map( A1 => n11615, A2 => n12141, A3 => n12135, ZN => 
                           n12482);
   U503 : INV_X1 port map( A => n12482, ZN => n12879);
   U504 : OAI222_X1 port map( A1 => n12875, A2 => n11403, B1 => n12873, B2 => 
                           n11779, C1 => n12507, C2 => n12034, ZN => n12571);
   U505 : NOR4_X1 port map( A1 => n12541, A2 => DATA2(2), A3 => DATA2(1), A4 =>
                           n12829, ZN => n12883);
   U506 : CLKBUF_X1 port map( A => n12883, Z => n12545);
   U507 : AOI222_X1 port map( A1 => n12575, A2 => n12541, B1 => n12572, B2 => 
                           n12879, C1 => n12571, C2 => n12545, ZN => n11407);
   U508 : INV_X1 port map( A => n12917, ZN => n12603);
   U509 : INV_X1 port map( A => n12588, ZN => n12586);
   U510 : NAND2_X1 port map( A1 => n12586, A2 => n12579, ZN => n12578);
   U511 : OAI211_X1 port map( C1 => n12587, C2 => n11717, A => n12927, B => 
                           n11405, ZN => n11406);
   U512 : OAI22_X1 port map( A1 => n11407, A2 => n12603, B1 => n12578, B2 => 
                           n11406, ZN => n11408);
   U513 : OR4_X1 port map( A1 => n11411, A2 => n11410, A3 => n11409, A4 => 
                           n11408, ZN => OUTALU(13));
   U514 : INV_X1 port map( A => DATA2(4), ZN => n12957);
   U515 : OAI21_X1 port map( B1 => n12957, B2 => n11412, A => n11704, ZN => 
                           n12914);
   U516 : INV_X1 port map( A => n12914, ZN => n12442);
   U517 : OAI211_X1 port map( C1 => DATA2(2), C2 => DATA2(1), A => DATA2(3), B 
                           => DATA2(4), ZN => n12897);
   U518 : CLKBUF_X1 port map( A => n12897, Z => n12215);
   U519 : NOR3_X1 port map( A1 => n12957, A2 => n12958, A3 => n11413, ZN => 
                           n12439);
   U520 : NAND2_X1 port map( A1 => n12215, A2 => n12439, ZN => n12896);
   U521 : INV_X1 port map( A => n12829, ZN => n12211);
   U522 : CLKBUF_X1 port map( A => n12141, Z => n12206);
   U523 : AOI21_X1 port map( B1 => n12211, B2 => n11414, A => n12206, ZN => 
                           n12626);
   U524 : INV_X1 port map( A => n12141, ZN => n12880);
   U525 : AOI21_X1 port map( B1 => DATA1(17), B2 => n12223, A => n11415, ZN => 
                           n11419);
   U526 : NAND2_X1 port map( A1 => DATA1(15), A2 => n12017, ZN => n11418);
   U527 : AND4_X1 port map( A1 => n11419, A2 => n11418, A3 => n11417, A4 => 
                           n11416, ZN => n11448);
   U528 : AND3_X1 port map( A1 => n11422, A2 => n11421, A3 => n11420, ZN => 
                           n11424);
   U529 : OAI211_X1 port map( C1 => n12186, C2 => n12491, A => n11424, B => 
                           n11423, ZN => n11469);
   U530 : INV_X1 port map( A => n11469, ZN => n11446);
   U531 : AOI211_X1 port map( C1 => DATA1(16), C2 => n11752, A => n11426, B => 
                           n11425, ZN => n11429);
   U532 : AND3_X1 port map( A1 => n11429, A2 => n11428, A3 => n11427, ZN => 
                           n11449);
   U533 : OAI222_X1 port map( A1 => n11448, A2 => n12109, B1 => n11446, B2 => 
                           n12113, C1 => n11449, C2 => n12111, ZN => n11519);
   U534 : INV_X1 port map( A => n11519, ZN => n11472);
   U535 : NOR2_X1 port map( A1 => n12220, A2 => n12469, ZN => n11432);
   U536 : INV_X1 port map( A => DATA1(14), ZN => n12548);
   U537 : NAND2_X1 port map( A1 => n12018, A2 => DATA1(15), ZN => n11753);
   U538 : OAI211_X1 port map( C1 => n12186, C2 => n12548, A => n11430, B => 
                           n11753, ZN => n11431);
   U539 : AOI211_X1 port map( C1 => DATA1(17), C2 => n12835, A => n11432, B => 
                           n11431, ZN => n11447);
   U540 : NAND2_X1 port map( A1 => n12018, A2 => DATA1(14), ZN => n11766);
   U541 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12017, ZN => n11435);
   U542 : NAND4_X1 port map( A1 => n11766, A2 => n11435, A3 => n11434, A4 => 
                           n11433, ZN => n11436);
   U543 : AOI21_X1 port map( B1 => n12834, B2 => DATA1(17), A => n11436, ZN => 
                           n11457);
   U544 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12018, ZN => n11784);
   U545 : NAND2_X1 port map( A1 => n12223, A2 => DATA1(14), ZN => n11755);
   U546 : AND3_X1 port map( A1 => n11755, A2 => n11438, A3 => n11437, ZN => 
                           n11439);
   U547 : OAI211_X1 port map( C1 => n12772, C2 => n12186, A => n11784, B => 
                           n11439, ZN => n11458);
   U548 : INV_X1 port map( A => n11458, ZN => n11440);
   U549 : OAI222_X1 port map( A1 => n12002, A2 => n11447, B1 => n12111, B2 => 
                           n11457, C1 => n12109, C2 => n11440, ZN => n11500);
   U550 : NAND3_X1 port map( A1 => n11443, A2 => n11442, A3 => n11441, ZN => 
                           n11444);
   U551 : AOI211_X1 port map( C1 => DATA1(18), C2 => n12017, A => n11445, B => 
                           n11444, ZN => n11468);
   U552 : OAI222_X1 port map( A1 => n12002, A2 => n11468, B1 => n12111, B2 => 
                           n11446, C1 => n11954, C2 => n11449, ZN => n11518);
   U553 : AOI22_X1 port map( A1 => n12030, A2 => n11500, B1 => n12115, B2 => 
                           n11518, ZN => n11451);
   U554 : OAI222_X1 port map( A1 => n12113, A2 => n11448, B1 => n12111, B2 => 
                           n11447, C1 => n12109, C2 => n11457, ZN => n11479);
   U555 : OAI222_X1 port map( A1 => n12002, A2 => n11449, B1 => n12111, B2 => 
                           n11448, C1 => n11954, C2 => n11447, ZN => n11488);
   U556 : AOI22_X1 port map( A1 => n12857, A2 => n11479, B1 => n12117, B2 => 
                           n11488, ZN => n11450);
   U557 : OAI211_X1 port map( C1 => n11472, C2 => n12850, A => n11451, B => 
                           n11450, ZN => n11555);
   U558 : NAND2_X1 port map( A1 => DATA1(13), A2 => n12223, ZN => n11765);
   U559 : AND3_X1 port map( A1 => n11765, A2 => n11453, A3 => n11452, ZN => 
                           n11454);
   U560 : NAND2_X1 port map( A1 => DATA1(12), A2 => n12018, ZN => n11801);
   U561 : OAI211_X1 port map( C1 => n12186, C2 => n12595, A => n11454, B => 
                           n11801, ZN => n11460);
   U562 : NAND2_X1 port map( A1 => DATA1(12), A2 => n12223, ZN => n11783);
   U563 : NAND2_X1 port map( A1 => DATA1(11), A2 => n12018, ZN => n11826);
   U564 : NAND2_X1 port map( A1 => n12835, A2 => DATA1(13), ZN => n11754);
   U565 : NAND2_X1 port map( A1 => n13263, A2 => n11752, ZN => n11455);
   U566 : AND4_X1 port map( A1 => n11783, A2 => n11826, A3 => n11754, A4 => 
                           n11455, ZN => n11456);
   U567 : OAI21_X1 port map( B1 => n12220, B2 => n12548, A => n11456, ZN => 
                           n11499);
   U568 : AOI222_X1 port map( A1 => n11498, A2 => n12844, B1 => n11460, B2 => 
                           n12267, C1 => n11499, C2 => n12840, ZN => n11585);
   U569 : AOI222_X1 port map( A1 => n11499, A2 => n12844, B1 => n11458, B2 => 
                           n12267, C1 => n11460, C2 => n12840, ZN => n11568);
   U570 : OAI22_X1 port map( A1 => n12853, A2 => n11585, B1 => n11568, B2 => 
                           n12359, ZN => n11462);
   U571 : INV_X1 port map( A => n11500, ZN => n11475);
   U572 : INV_X1 port map( A => n11457, ZN => n11459);
   U573 : AOI222_X1 port map( A1 => n11460, A2 => n12844, B1 => n11459, B2 => 
                           n12842, C1 => n11458, C2 => n12840, ZN => n11496);
   U574 : OAI22_X1 port map( A1 => n11475, A2 => n12850, B1 => n11496, B2 => 
                           n12361, ZN => n11461);
   U575 : AOI211_X1 port map( C1 => n12115, C2 => n11479, A => n11462, B => 
                           n11461, ZN => n11596);
   U576 : INV_X1 port map( A => DATA1(23), ZN => n12333);
   U577 : NAND2_X1 port map( A1 => DATA1(19), A2 => n12017, ZN => n11466);
   U578 : AND4_X1 port map( A1 => n11466, A2 => n11465, A3 => n11464, A4 => 
                           n11463, ZN => n11467);
   U579 : OAI21_X1 port map( B1 => n12220, B2 => n12333, A => n11467, ZN => 
                           n11513);
   U580 : INV_X1 port map( A => n11468, ZN => n11487);
   U581 : AOI222_X1 port map( A1 => n11469, A2 => n12844, B1 => n11513, B2 => 
                           n12267, C1 => n11487, C2 => n12840, ZN => n11531);
   U582 : OAI22_X1 port map( A1 => n12415, A2 => n11531, B1 => n11472, B2 => 
                           n12361, ZN => n11471);
   U583 : INV_X1 port map( A => n11488, ZN => n11476);
   U584 : INV_X1 port map( A => n11518, ZN => n11491);
   U585 : OAI22_X1 port map( A1 => n11476, A2 => n12026, B1 => n11491, B2 => 
                           n12416, ZN => n11470);
   U586 : AOI211_X1 port map( C1 => n12030, C2 => n11479, A => n11471, B => 
                           n11470, ZN => n11493);
   U587 : OAI22_X1 port map( A1 => n12865, A2 => n11596, B1 => n11493, B2 => 
                           n12858, ZN => n11481);
   U588 : OAI22_X1 port map( A1 => n12415, A2 => n11472, B1 => n11475, B2 => 
                           n12359, ZN => n11474);
   U589 : OAI22_X1 port map( A1 => n12853, A2 => n11496, B1 => n11476, B2 => 
                           n12416, ZN => n11473);
   U590 : AOI211_X1 port map( C1 => n12117, C2 => n11479, A => n11474, B => 
                           n11473, ZN => n11597);
   U591 : OAI22_X1 port map( A1 => n11475, A2 => n12846, B1 => n11496, B2 => 
                           n12026, ZN => n11478);
   U592 : OAI22_X1 port map( A1 => n12853, A2 => n11568, B1 => n12849, B2 => 
                           n11476, ZN => n11477);
   U593 : AOI211_X1 port map( C1 => n12197, C2 => n11479, A => n11478, B => 
                           n11477, ZN => n11598);
   U594 : OAI22_X1 port map( A1 => n11597, A2 => n12860, B1 => n11598, B2 => 
                           n12473, ZN => n11480);
   U595 : AOI211_X1 port map( C1 => n12570, C2 => n11555, A => n11481, B => 
                           n11480, ZN => n11602);
   U596 : INV_X1 port map( A => n11531, ZN => n11515);
   U597 : INV_X1 port map( A => DATA1(24), ZN => n12723);
   U598 : NAND2_X1 port map( A1 => DATA1(20), A2 => n11752, ZN => n11485);
   U599 : AND4_X1 port map( A1 => n11485, A2 => n11484, A3 => n11483, A4 => 
                           n11482, ZN => n11486);
   U600 : OAI21_X1 port map( B1 => n12220, B2 => n12723, A => n11486, ZN => 
                           n11514);
   U601 : AOI222_X1 port map( A1 => n12842, A2 => n11514, B1 => n12193, B2 => 
                           n11513, C1 => n12192, C2 => n11487, ZN => n11546);
   U602 : INV_X1 port map( A => n11546, ZN => n11520);
   U603 : AOI22_X1 port map( A1 => n12197, A2 => n11515, B1 => n12115, B2 => 
                           n11520, ZN => n11490);
   U604 : AOI22_X1 port map( A1 => n12857, A2 => n11519, B1 => n12119, B2 => 
                           n11488, ZN => n11489);
   U605 : OAI211_X1 port map( C1 => n11491, C2 => n12846, A => n11490, B => 
                           n11489, ZN => n11556);
   U606 : INV_X1 port map( A => n11597, ZN => n11492);
   U607 : INV_X1 port map( A => n11598, ZN => n11595);
   U608 : AOI22_X1 port map( A1 => n12869, A2 => n11492, B1 => n12128, B2 => 
                           n11595, ZN => n11495);
   U609 : INV_X1 port map( A => n11493, ZN => n11554);
   U610 : AOI22_X1 port map( A1 => n12570, A2 => n11554, B1 => n12569, B2 => 
                           n11555, ZN => n11494);
   U611 : NAND2_X1 port map( A1 => n11495, A2 => n11494, ZN => n11562);
   U612 : AOI21_X1 port map( B1 => n12617, B2 => n11556, A => n11562, ZN => 
                           n11560);
   U613 : INV_X1 port map( A => n11496, ZN => n11571);
   U614 : AOI222_X1 port map( A1 => n12842, A2 => n11499, B1 => n12193, B2 => 
                           n11498, C1 => n12192, C2 => n11497, ZN => n11582);
   U615 : INV_X1 port map( A => n11582, ZN => n11581);
   U616 : AOI22_X1 port map( A1 => n12197, A2 => n11571, B1 => n12119, B2 => 
                           n11581, ZN => n11502);
   U617 : INV_X1 port map( A => n11568, ZN => n11588);
   U618 : AOI22_X1 port map( A1 => n12117, A2 => n11588, B1 => n12115, B2 => 
                           n11500, ZN => n11501);
   U619 : OAI211_X1 port map( C1 => n11585, C2 => n12359, A => n11502, B => 
                           n11501, ZN => n11601);
   U620 : INV_X1 port map( A => n11555, ZN => n11525);
   U621 : OAI22_X1 port map( A1 => n11596, A2 => n12473, B1 => n11525, B2 => 
                           n12858, ZN => n11504);
   U622 : OAI22_X1 port map( A1 => n11597, A2 => n12862, B1 => n11598, B2 => 
                           n12860, ZN => n11503);
   U623 : AOI211_X1 port map( C1 => n12128, C2 => n11601, A => n11504, B => 
                           n11503, ZN => n11604);
   U624 : OAI222_X1 port map( A1 => n12875, A2 => n11602, B1 => n12873, B2 => 
                           n11560, C1 => n11604, C2 => n12034, ZN => n11637);
   U625 : INV_X1 port map( A => n12541, ZN => n12514);
   U626 : AOI22_X1 port map( A1 => DATA1(23), A2 => n11853, B1 => DATA1(22), B2
                           => n12017, ZN => n11508);
   U627 : NAND4_X1 port map( A1 => n11508, A2 => n11507, A3 => n11506, A4 => 
                           n11505, ZN => n11544);
   U628 : AOI22_X1 port map( A1 => DATA1(22), A2 => n12018, B1 => DATA1(21), B2
                           => n12017, ZN => n11512);
   U629 : NAND2_X1 port map( A1 => n12189, A2 => n12295, ZN => n11509);
   U630 : NAND4_X1 port map( A1 => n11512, A2 => n11511, A3 => n11510, A4 => 
                           n11509, ZN => n11530);
   U631 : AOI222_X1 port map( A1 => n11514, A2 => n12844, B1 => n11544, B2 => 
                           n12842, C1 => n11530, C2 => n12840, ZN => n12083);
   U632 : AOI222_X1 port map( A1 => n12842, A2 => n11530, B1 => n12193, B2 => 
                           n11514, C1 => n12192, C2 => n11513, ZN => n11547);
   U633 : INV_X1 port map( A => n11547, ZN => n11647);
   U634 : AOI22_X1 port map( A1 => n12857, A2 => n11515, B1 => n12197, B2 => 
                           n11647, ZN => n11517);
   U635 : AOI22_X1 port map( A1 => n12117, A2 => n11520, B1 => n12119, B2 => 
                           n11518, ZN => n11516);
   U636 : OAI211_X1 port map( C1 => n12415, C2 => n12083, A => n11517, B => 
                           n11516, ZN => n12084);
   U637 : AOI22_X1 port map( A1 => n12126, A2 => n11556, B1 => n12617, B2 => 
                           n12084, ZN => n11524);
   U638 : CLKBUF_X1 port map( A => n12570, Z => n12594);
   U639 : AOI22_X1 port map( A1 => n12857, A2 => n11518, B1 => n12115, B2 => 
                           n11647, ZN => n11522);
   U640 : AOI22_X1 port map( A1 => n12197, A2 => n11520, B1 => n12119, B2 => 
                           n11519, ZN => n11521);
   U641 : OAI211_X1 port map( C1 => n11531, C2 => n12846, A => n11522, B => 
                           n11521, ZN => n11650);
   U642 : AOI22_X1 port map( A1 => n12594, A2 => n11650, B1 => n12425, B2 => 
                           n11554, ZN => n11523);
   U643 : OAI211_X1 port map( C1 => n12865, C2 => n11525, A => n11524, B => 
                           n11523, ZN => n11564);
   U644 : INV_X1 port map( A => n12084, ZN => n11553);
   U645 : AOI22_X1 port map( A1 => n12740, A2 => n11853, B1 => DATA1(23), B2 =>
                           n12017, ZN => n11529);
   U646 : NAND4_X1 port map( A1 => n11529, A2 => n11528, A3 => n11527, A4 => 
                           n11526, ZN => n11543);
   U647 : AOI222_X1 port map( A1 => n11530, A2 => n12844, B1 => n11543, B2 => 
                           n12267, C1 => n11544, C2 => n12840, ZN => n11538);
   U648 : OAI22_X1 port map( A1 => n12415, A2 => n11538, B1 => n11546, B2 => 
                           n12359, ZN => n11533);
   U649 : OAI22_X1 port map( A1 => n12853, A2 => n11531, B1 => n12083, B2 => 
                           n12416, ZN => n11532);
   U650 : AOI211_X1 port map( C1 => n12117, C2 => n11647, A => n11533, B => 
                           n11532, ZN => n12087);
   U651 : AOI22_X1 port map( A1 => n12869, A2 => n11556, B1 => n11960, B2 => 
                           n11554, ZN => n11534);
   U652 : OAI21_X1 port map( B1 => n12087, B2 => n12471, A => n11534, ZN => 
                           n11535);
   U653 : INV_X1 port map( A => n11535, ZN => n11536);
   U654 : OAI21_X1 port map( B1 => n12862, B2 => n11553, A => n11536, ZN => 
                           n11653);
   U655 : AOI21_X1 port map( B1 => n11650, B2 => n12569, A => n11653, ZN => 
                           n11537);
   U656 : INV_X1 port map( A => n11537, ZN => n11563);
   U657 : INV_X1 port map( A => n12087, ZN => n12127);
   U658 : INV_X1 port map( A => n11538, ZN => n12118);
   U659 : NOR2_X1 port map( A1 => n12105, A2 => n12723, ZN => n11542);
   U660 : OAI211_X1 port map( C1 => n12220, C2 => n12244, A => n11540, B => 
                           n11539, ZN => n11541);
   U661 : AOI211_X1 port map( C1 => n12018, C2 => DATA1(25), A => n11542, B => 
                           n11541, ZN => n12078);
   U662 : INV_X1 port map( A => n11543, ZN => n11645);
   U663 : INV_X1 port map( A => n11544, ZN => n11545);
   U664 : OAI222_X1 port map( A1 => n12002, A2 => n12078, B1 => n12111, B2 => 
                           n11645, C1 => n12109, C2 => n11545, ZN => n12079);
   U665 : INV_X1 port map( A => n12079, ZN => n12123);
   U666 : OAI22_X1 port map( A1 => n12846, A2 => n12083, B1 => n12849, B2 => 
                           n12123, ZN => n11549);
   U667 : OAI22_X1 port map( A1 => n12359, A2 => n11547, B1 => n12853, B2 => 
                           n11546, ZN => n11548);
   U668 : AOI211_X1 port map( C1 => n12118, C2 => n12197, A => n11549, B => 
                           n11548, ZN => n11550);
   U669 : INV_X1 port map( A => n11550, ZN => n12129);
   U670 : AOI22_X1 port map( A1 => n12594, A2 => n12127, B1 => n12617, B2 => 
                           n12129, ZN => n11552);
   U671 : AOI22_X1 port map( A1 => n12869, A2 => n11650, B1 => n11960, B2 => 
                           n11556, ZN => n11551);
   U672 : OAI211_X1 port map( C1 => n11553, C2 => n12860, A => n11552, B => 
                           n11551, ZN => n12088);
   U673 : AOI222_X1 port map( A1 => n11564, A2 => n12135, B1 => n11563, B2 => 
                           n12526, C1 => n12088, C2 => n12550, ZN => n12139);
   U674 : AOI22_X1 port map( A1 => n12126, A2 => n11554, B1 => n12617, B2 => 
                           n11650, ZN => n11558);
   U675 : AOI22_X1 port map( A1 => n12570, A2 => n11556, B1 => n12869, B2 => 
                           n11555, ZN => n11557);
   U676 : OAI211_X1 port map( C1 => n12865, C2 => n11597, A => n11558, B => 
                           n11557, ZN => n11565);
   U677 : INV_X1 port map( A => n11565, ZN => n11559);
   U678 : OAI222_X1 port map( A1 => n11602, A2 => n12870, B1 => n11560, B2 => 
                           n12875, C1 => n11559, C2 => n12506, ZN => n11655);
   U679 : INV_X1 port map( A => n11655, ZN => n11620);
   U680 : NOR3_X1 port map( A1 => n12957, A2 => n11561, A3 => n12880, ZN => 
                           n12573);
   U681 : INV_X1 port map( A => n12573, ZN => n12886);
   U682 : OAI22_X1 port map( A1 => n12514, A2 => n12139, B1 => n11620, B2 => 
                           n12886, ZN => n11567);
   U683 : AOI222_X1 port map( A1 => n11562, A2 => n12135, B1 => n11565, B2 => 
                           n12526, C1 => n11564, C2 => n12550, ZN => n12089);
   U684 : AOI222_X1 port map( A1 => n11565, A2 => n12135, B1 => n11564, B2 => 
                           n12526, C1 => n11563, C2 => n12550, ZN => n12140);
   U685 : INV_X1 port map( A => n12883, ZN => n12495);
   U686 : OAI22_X1 port map( A1 => n12089, A2 => n12482, B1 => n12140, B2 => 
                           n12495, ZN => n11566);
   U687 : AOI211_X1 port map( C1 => n12880, C2 => n11637, A => n11567, B => 
                           n11566, ZN => n12071);
   U688 : OAI22_X1 port map( A1 => n12846, A2 => n11585, B1 => n12853, B2 => 
                           n11584, ZN => n11570);
   U689 : OAI22_X1 port map( A1 => n12026, A2 => n11582, B1 => n12416, B2 => 
                           n11568, ZN => n11569);
   U690 : AOI211_X1 port map( C1 => n12080, C2 => n11571, A => n11570, B => 
                           n11569, ZN => n11628);
   U691 : AOI22_X1 port map( A1 => n12117, A2 => n11573, B1 => n12119, B2 => 
                           n11572, ZN => n11576);
   U692 : AOI22_X1 port map( A1 => n12857, A2 => n11574, B1 => n12115, B2 => 
                           n11581, ZN => n11575);
   U693 : OAI211_X1 port map( C1 => n11584, C2 => n12850, A => n11576, B => 
                           n11575, ZN => n11689);
   U694 : INV_X1 port map( A => n11689, ZN => n11577);
   U695 : OAI22_X1 port map( A1 => n12862, A2 => n11628, B1 => n12865, B2 => 
                           n11577, ZN => n11590);
   U696 : OAI22_X1 port map( A1 => n12853, A2 => n11578, B1 => n11584, B2 => 
                           n12361, ZN => n11580);
   U697 : OAI22_X1 port map( A1 => n12415, A2 => n11585, B1 => n11583, B2 => 
                           n12026, ZN => n11579);
   U698 : AOI211_X1 port map( C1 => n12197, C2 => n11581, A => n11580, B => 
                           n11579, ZN => n11678);
   U699 : OAI22_X1 port map( A1 => n12853, A2 => n11583, B1 => n11582, B2 => 
                           n12361, ZN => n11587);
   U700 : OAI22_X1 port map( A1 => n11585, A2 => n12850, B1 => n11584, B2 => 
                           n12026, ZN => n11586);
   U701 : AOI211_X1 port map( C1 => n12115, C2 => n11588, A => n11587, B => 
                           n11586, ZN => n11681);
   U702 : OAI22_X1 port map( A1 => n12473, A2 => n11678, B1 => n12860, B2 => 
                           n11681, ZN => n11589);
   U703 : NOR2_X1 port map( A1 => n11590, A2 => n11589, ZN => n11625);
   U704 : OAI22_X1 port map( A1 => n12865, A2 => n11678, B1 => n11628, B2 => 
                           n12860, ZN => n11592);
   U705 : OAI22_X1 port map( A1 => n11596, A2 => n12858, B1 => n11681, B2 => 
                           n12473, ZN => n11591);
   U706 : AOI211_X1 port map( C1 => n12594, C2 => n11601, A => n11592, B => 
                           n11591, ZN => n11627);
   U707 : INV_X1 port map( A => n11601, ZN => n11626);
   U708 : OAI22_X1 port map( A1 => n12865, A2 => n11681, B1 => n11626, B2 => 
                           n12860, ZN => n11594);
   U709 : OAI22_X1 port map( A1 => n11596, A2 => n12862, B1 => n11628, B2 => 
                           n12473, ZN => n11593);
   U710 : AOI211_X1 port map( C1 => n12617, C2 => n11595, A => n11594, B => 
                           n11593, ZN => n11603);
   U711 : OAI222_X1 port map( A1 => n11625, A2 => n12034, B1 => n11627, B2 => 
                           n12875, C1 => n11603, C2 => n12506, ZN => n11624);
   U712 : INV_X1 port map( A => n11624, ZN => n11694);
   U713 : CLKBUF_X1 port map( A => n12573, Z => n12203);
   U714 : OAI22_X1 port map( A1 => n12860, A2 => n11596, B1 => n12865, B2 => 
                           n11628, ZN => n11600);
   U715 : OAI22_X1 port map( A1 => n12862, A2 => n11598, B1 => n12858, B2 => 
                           n11597, ZN => n11599);
   U716 : AOI211_X1 port map( C1 => n11601, C2 => n12425, A => n11600, B => 
                           n11599, ZN => n11605);
   U717 : OAI222_X1 port map( A1 => n12875, A2 => n11603, B1 => n12873, B2 => 
                           n11605, C1 => n11627, C2 => n12870, ZN => n11664);
   U718 : OAI222_X1 port map( A1 => n11605, A2 => n12034, B1 => n11604, B2 => 
                           n12875, C1 => n11602, C2 => n12506, ZN => n11633);
   U719 : INV_X1 port map( A => n11633, ZN => n11614);
   U720 : OAI222_X1 port map( A1 => n12875, A2 => n11605, B1 => n12873, B2 => 
                           n11604, C1 => n11603, C2 => n12034, ZN => n11617);
   U721 : INV_X1 port map( A => n11617, ZN => n11674);
   U722 : OAI22_X1 port map( A1 => n11614, A2 => n12495, B1 => n11674, B2 => 
                           n12482, ZN => n11606);
   U723 : AOI21_X1 port map( B1 => n12203, B2 => n11664, A => n11606, ZN => 
                           n11607);
   U724 : OAI21_X1 port map( B1 => n12206, B2 => n11694, A => n11607, ZN => 
                           n11636);
   U725 : NAND3_X1 port map( A1 => n12958, A2 => n11616, A3 => n11608, ZN => 
                           n12436);
   U726 : INV_X1 port map( A => n12436, ZN => n12891);
   U727 : AOI22_X1 port map( A1 => n12541, A2 => n11655, B1 => n12880, B2 => 
                           n11664, ZN => n11610);
   U728 : AOI22_X1 port map( A1 => n12883, A2 => n11637, B1 => n12203, B2 => 
                           n11617, ZN => n11609);
   U729 : OAI211_X1 port map( C1 => n11614, C2 => n12482, A => n11610, B => 
                           n11609, ZN => n11659);
   U730 : AOI22_X1 port map( A1 => n12829, A2 => n11636, B1 => n12891, B2 => 
                           n11659, ZN => n11622);
   U731 : NOR3_X1 port map( A1 => DATA2(3), A2 => n11611, A3 => n11672, ZN => 
                           n12831);
   U732 : INV_X1 port map( A => n12140, ZN => n11654);
   U733 : AOI22_X1 port map( A1 => n12879, A2 => n11655, B1 => n12877, B2 => 
                           n11654, ZN => n11613);
   U734 : INV_X1 port map( A => n12089, ZN => n11656);
   U735 : AOI22_X1 port map( A1 => n12545, A2 => n11656, B1 => n12203, B2 => 
                           n11637, ZN => n11612);
   U736 : OAI211_X1 port map( C1 => n12206, C2 => n11614, A => n11613, B => 
                           n11612, ZN => n12072);
   U737 : NAND3_X1 port map( A1 => n11616, A2 => n11615, A3 => n12211, ZN => 
                           n12894);
   U738 : INV_X1 port map( A => n12894, ZN => n12431);
   U739 : AOI22_X1 port map( A1 => n12879, A2 => n11637, B1 => n12880, B2 => 
                           n11617, ZN => n11619);
   U740 : AOI22_X1 port map( A1 => n12573, A2 => n11633, B1 => n12877, B2 => 
                           n11656, ZN => n11618);
   U741 : OAI211_X1 port map( C1 => n11620, C2 => n12495, A => n11619, B => 
                           n11618, ZN => n11660);
   U742 : AOI22_X1 port map( A1 => n12831, A2 => n12072, B1 => n12431, B2 => 
                           n11660, ZN => n11621);
   U743 : OAI211_X1 port map( C1 => n12626, C2 => n12071, A => n11622, B => 
                           n11621, ZN => n11623);
   U744 : INV_X1 port map( A => n11623, ZN => n12097);
   U745 : CLKBUF_X1 port map( A => n12626, Z => n12604);
   U746 : INV_X1 port map( A => n12604, ZN => n12889);
   U747 : AOI22_X1 port map( A1 => n12203, A2 => n11624, B1 => n12879, B2 => 
                           n11664, ZN => n11635);
   U748 : OAI21_X1 port map( B1 => n12858, B2 => n11626, A => n11625, ZN => 
                           n11667);
   U749 : INV_X1 port map( A => n11627, ZN => n11632);
   U750 : OAI22_X1 port map( A1 => n12865, A2 => n11692, B1 => n11678, B2 => 
                           n12860, ZN => n11630);
   U751 : OAI22_X1 port map( A1 => n11628, A2 => n12471, B1 => n11681, B2 => 
                           n12862, ZN => n11629);
   U752 : AOI211_X1 port map( C1 => n12869, C2 => n11689, A => n11630, B => 
                           n11629, ZN => n11631);
   U753 : INV_X1 port map( A => n11631, ZN => n11682);
   U754 : AOI222_X1 port map( A1 => n12526, A2 => n11667, B1 => n12550, B2 => 
                           n11632, C1 => n11682, C2 => n12135, ZN => n12456);
   U755 : INV_X1 port map( A => n12456, ZN => n11697);
   U756 : AOI22_X1 port map( A1 => n12541, A2 => n11633, B1 => n12880, B2 => 
                           n11697, ZN => n11634);
   U757 : OAI211_X1 port map( C1 => n11674, C2 => n12495, A => n11635, B => 
                           n11634, ZN => n11702);
   U758 : INV_X1 port map( A => n11702, ZN => n12332);
   U759 : INV_X1 port map( A => n11659, ZN => n11686);
   U760 : OAI22_X1 port map( A1 => n12332, A2 => n12211, B1 => n11686, B2 => 
                           n12894, ZN => n11639);
   U761 : AOI21_X1 port map( B1 => n12541, B2 => n11637, A => n11636, ZN => 
                           n11699);
   U762 : INV_X1 port map( A => n11660, ZN => n12094);
   U763 : INV_X1 port map( A => n12831, ZN => n12623);
   U764 : OAI22_X1 port map( A1 => n11699, A2 => n12436, B1 => n12094, B2 => 
                           n12623, ZN => n11638);
   U765 : AOI211_X1 port map( C1 => n12889, C2 => n12072, A => n11639, B => 
                           n11638, ZN => n11705);
   U766 : INV_X1 port map( A => n12083, ZN => n11646);
   U767 : NAND2_X1 port map( A1 => n12295, A2 => n12017, ZN => n11643);
   U768 : NAND4_X1 port map( A1 => n11643, A2 => n11642, A3 => n11641, A4 => 
                           n11640, ZN => n11644);
   U769 : AOI21_X1 port map( B1 => n12189, B2 => DATA1(29), A => n11644, ZN => 
                           n12108);
   U770 : OAI222_X1 port map( A1 => n12113, A2 => n12108, B1 => n12111, B2 => 
                           n12078, C1 => n11954, C2 => n11645, ZN => n12116);
   U771 : AOI22_X1 port map( A1 => n12857, A2 => n11646, B1 => n12080, B2 => 
                           n12116, ZN => n11649);
   U772 : AOI22_X1 port map( A1 => n12117, A2 => n12118, B1 => n12119, B2 => 
                           n11647, ZN => n11648);
   U773 : OAI211_X1 port map( C1 => n12123, C2 => n12850, A => n11649, B => 
                           n11648, ZN => n12125);
   U774 : AOI22_X1 port map( A1 => n12869, A2 => n12084, B1 => n12617, B2 => 
                           n12125, ZN => n11652);
   U775 : AOI22_X1 port map( A1 => n12594, A2 => n12129, B1 => n11960, B2 => 
                           n11650, ZN => n11651);
   U776 : OAI211_X1 port map( C1 => n12087, C2 => n12860, A => n11652, B => 
                           n11651, ZN => n12136);
   U777 : AOI222_X1 port map( A1 => n11653, A2 => n12135, B1 => n12088, B2 => 
                           n12526, C1 => n12136, C2 => n12550, ZN => n12137);
   U778 : INV_X1 port map( A => n12137, ZN => n12092);
   U779 : AOI22_X1 port map( A1 => n12879, A2 => n11654, B1 => n12877, B2 => 
                           n12092, ZN => n11658);
   U780 : AOI22_X1 port map( A1 => n12203, A2 => n11656, B1 => n12880, B2 => 
                           n11655, ZN => n11657);
   U781 : OAI211_X1 port map( C1 => n12139, C2 => n12495, A => n11658, B => 
                           n11657, ZN => n12093);
   U782 : AOI22_X1 port map( A1 => n12829, A2 => n11659, B1 => n12889, B2 => 
                           n12093, ZN => n11662);
   U783 : AOI22_X1 port map( A1 => n12891, A2 => n11660, B1 => n12431, B2 => 
                           n12072, ZN => n11661);
   U784 : OAI211_X1 port map( C1 => n12071, C2 => n12623, A => n11662, B => 
                           n11661, ZN => n11663);
   U785 : INV_X1 port map( A => n11663, ZN => n12151);
   U786 : OAI222_X1 port map( A1 => n12896, A2 => n12097, B1 => n12215, B2 => 
                           n11705, C1 => n12151, C2 => n12439, ZN => n12161);
   U787 : NAND2_X1 port map( A1 => n11704, A2 => n12914, ZN => n12446);
   U788 : INV_X1 port map( A => n12446, ZN => n12907);
   U789 : INV_X1 port map( A => n11664, ZN => n11683);
   U790 : OAI22_X1 port map( A1 => n11694, A2 => n12482, B1 => n11683, B2 => 
                           n12495, ZN => n11669);
   U791 : AOI22_X1 port map( A1 => n12869, A2 => n11675, B1 => n12569, B2 => 
                           n11689, ZN => n11666);
   U792 : NAND2_X1 port map( A1 => n12128, A2 => n12568, ZN => n11665);
   U793 : OAI211_X1 port map( C1 => n11678, C2 => n12862, A => n11666, B => 
                           n11665, ZN => n11679);
   U794 : AOI222_X1 port map( A1 => n11679, A2 => n12135, B1 => n11682, B2 => 
                           n12526, C1 => n11667, C2 => n12550, ZN => n12481);
   U795 : OAI22_X1 port map( A1 => n12141, A2 => n12481, B1 => n12456, B2 => 
                           n12886, ZN => n11668);
   U796 : NOR2_X1 port map( A1 => n11669, A2 => n11668, ZN => n11673);
   U797 : OAI22_X1 port map( A1 => n11699, A2 => n12894, B1 => n11673, B2 => 
                           n12211, ZN => n11671);
   U798 : OAI22_X1 port map( A1 => n12604, A2 => n12094, B1 => n11686, B2 => 
                           n12623, ZN => n11670);
   U799 : AOI211_X1 port map( C1 => n12891, C2 => n11702, A => n11671, B => 
                           n11670, ZN => n11706);
   U800 : CLKBUF_X1 port map( A => n12439, Z => n12213);
   U801 : OAI222_X1 port map( A1 => n12896, A2 => n11705, B1 => n12215, B2 => 
                           n11706, C1 => n12097, C2 => n12213, ZN => n12236);
   U802 : AOI22_X1 port map( A1 => n12442, A2 => n12161, B1 => n12907, B2 => 
                           n12236, ZN => n11708);
   U803 : NOR2_X1 port map( A1 => n11704, A2 => n11672, ZN => n12909);
   U804 : OAI21_X1 port map( B1 => n12514, B2 => n11674, A => n11673, ZN => 
                           n11698);
   U805 : OAI22_X1 port map( A1 => n11699, A2 => n12623, B1 => n12332, B2 => 
                           n12894, ZN => n11688);
   U806 : AOI22_X1 port map( A1 => n12126, A2 => n11675, B1 => n11960, B2 => 
                           n12593, ZN => n11677);
   U807 : AOI22_X1 port map( A1 => n12594, A2 => n11689, B1 => n12869, B2 => 
                           n12568, ZN => n11676);
   U808 : OAI211_X1 port map( C1 => n11678, C2 => n12471, A => n11677, B => 
                           n11676, ZN => n12527);
   U809 : INV_X1 port map( A => n11679, ZN => n11680);
   U810 : OAI21_X1 port map( B1 => n11681, B2 => n12471, A => n11680, ZN => 
                           n11693);
   U811 : AOI222_X1 port map( A1 => n12527, A2 => n12135, B1 => n11693, B2 => 
                           n12526, C1 => n11682, C2 => n12550, ZN => n12496);
   U812 : OAI22_X1 port map( A1 => n12206, A2 => n12496, B1 => n12481, B2 => 
                           n12886, ZN => n11685);
   U813 : OAI22_X1 port map( A1 => n12514, A2 => n11683, B1 => n11694, B2 => 
                           n12495, ZN => n11684);
   U814 : AOI211_X1 port map( C1 => n12879, C2 => n11697, A => n11685, B => 
                           n11684, ZN => n12373);
   U815 : OAI22_X1 port map( A1 => n12604, A2 => n11686, B1 => n12373, B2 => 
                           n12211, ZN => n11687);
   U816 : AOI211_X1 port map( C1 => n12891, C2 => n11698, A => n11688, B => 
                           n11687, ZN => n12303);
   U817 : AOI22_X1 port map( A1 => n12569, A2 => n12568, B1 => n11960, B2 => 
                           n12619, ZN => n11691);
   U818 : AOI22_X1 port map( A1 => n12425, A2 => n12593, B1 => n12617, B2 => 
                           n11689, ZN => n11690);
   U819 : OAI211_X1 port map( C1 => n11692, C2 => n12862, A => n11691, B => 
                           n11690, ZN => n12549);
   U820 : AOI222_X1 port map( A1 => n12549, A2 => n12135, B1 => n12527, B2 => 
                           n12526, C1 => n11693, C2 => n12550, ZN => n12513);
   U821 : OAI22_X1 port map( A1 => n12141, A2 => n12513, B1 => n12481, B2 => 
                           n12482, ZN => n11696);
   U822 : OAI22_X1 port map( A1 => n12514, A2 => n11694, B1 => n12496, B2 => 
                           n12886, ZN => n11695);
   U823 : AOI211_X1 port map( C1 => n12545, C2 => n11697, A => n11696, B => 
                           n11695, ZN => n12384);
   U824 : OAI22_X1 port map( A1 => n12384, A2 => n12211, B1 => n12373, B2 => 
                           n12436, ZN => n11701);
   U825 : INV_X1 port map( A => n11698, ZN => n12351);
   U826 : OAI22_X1 port map( A1 => n12604, A2 => n11699, B1 => n12351, B2 => 
                           n12894, ZN => n11700);
   U827 : AOI211_X1 port map( C1 => n12831, C2 => n11702, A => n11701, B => 
                           n11700, ZN => n12318);
   U828 : OAI222_X1 port map( A1 => n12896, A2 => n12303, B1 => n12897, B2 => 
                           n12318, C1 => n11706, C2 => n12213, ZN => n12289);
   U829 : NOR2_X1 port map( A1 => n11704, A2 => n11703, ZN => n12905);
   U830 : OAI222_X1 port map( A1 => n12896, A2 => n11706, B1 => n12215, B2 => 
                           n12303, C1 => n11705, C2 => n12213, ZN => n12263);
   U831 : AOI22_X1 port map( A1 => n12909, A2 => n12289, B1 => n12905, B2 => 
                           n12263, ZN => n11707);
   U832 : AOI21_X1 port map( B1 => n11708, B2 => n11707, A => n12610, ZN => 
                           n11735);
   U833 : INV_X1 port map( A => DATA1(29), ZN => n12073);
   U834 : NOR2_X1 port map( A1 => n12220, A2 => n12073, ZN => n11709);
   U835 : NOR2_X1 port map( A1 => n12396, A2 => n12825, ZN => n12107);
   U836 : AOI211_X1 port map( C1 => DATA1(31), C2 => n12223, A => n11709, B => 
                           n12107, ZN => n11712);
   U837 : NAND2_X1 port map( A1 => DATA2(29), A2 => n12073, ZN => n12819);
   U838 : NOR2_X1 port map( A1 => n12073, A2 => DATA2(29), ZN => n12731);
   U839 : INV_X1 port map( A => n12731, ZN => n12816);
   U840 : NAND2_X1 port map( A1 => n12819, A2 => n12816, ZN => n12656);
   U841 : AOI22_X1 port map( A1 => dataout_mul_29_port, A2 => n12615, B1 => 
                           n12622, B2 => n12656, ZN => n11711);
   U842 : INV_X1 port map( A => n12616, ZN => n12580);
   U843 : NAND3_X1 port map( A1 => DATA2(29), A2 => DATA1(29), A3 => n12580, ZN
                           => n11710);
   U844 : OAI211_X1 port map( C1 => n11712, C2 => n12603, A => n11711, B => 
                           n11710, ZN => n11734);
   U845 : NAND2_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, ZN => 
                           n11725);
   U846 : OAI21_X1 port map( B1 => DATA1(23), B2 => DATA2_I_23_port, A => 
                           n11725, ZN => n12346);
   U847 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n12347);
   U848 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n12328);
   U849 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => 
                           n12328, ZN => n11723);
   U850 : NAND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n12330);
   U851 : OAI21_X1 port map( B1 => DATA1(21), B2 => DATA2_I_21_port, A => 
                           n12330, ZN => n12380);
   U852 : XOR2_X1 port map( A => DATA2_I_18_port, B => DATA1(18), Z => n12490);
   U853 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n12511);
   U854 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n12325);
   U855 : OAI21_X1 port map( B1 => DATA1(17), B2 => DATA2_I_17_port, A => 
                           n12325, ZN => n12503);
   U856 : NOR2_X1 port map( A1 => n12511, A2 => n12503, ZN => n12323);
   U857 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n12326);
   U858 : AOI21_X1 port map( B1 => DATA2_I_19_port, B2 => DATA1(19), A => 
                           n12326, ZN => n12452);
   U859 : NAND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n11720);
   U860 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => 
                           n11720, ZN => n12535);
   U861 : XOR2_X1 port map( A => DATA2_I_14_port, B => DATA1(14), Z => n12559);
   U862 : NAND2_X1 port map( A1 => n11713, A2 => n12556, ZN => n12553);
   U863 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n12559, B2 => n12553, ZN => n12528);
   U864 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => DATA1(8), A => n11818,
                           ZN => n11852);
   U865 : INV_X1 port map( A => n12559, ZN => n11716);
   U866 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => 
                           n11714, ZN => n12601);
   U867 : NOR4_X1 port map( A1 => n11716, A2 => n11820, A3 => n11715, A4 => 
                           n12601, ZN => n11718);
   U868 : NAND4_X1 port map( A1 => n11719, A2 => n11852, A3 => n11718, A4 => 
                           n11717, ZN => n11721);
   U869 : OAI221_X1 port map( B1 => n12535, B2 => n12528, C1 => n12535, C2 => 
                           n11721, A => n11720, ZN => n12331);
   U870 : NAND4_X1 port map( A1 => n12490, A2 => n12323, A3 => n12452, A4 => 
                           n12331, ZN => n11722);
   U871 : NOR3_X1 port map( A1 => n11723, A2 => n12380, A3 => n11722, ZN => 
                           n11724);
   U872 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n12510);
   U873 : OAI21_X1 port map( B1 => n12510, B2 => n12503, A => n12325, ZN => 
                           n12484);
   U874 : AOI22_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, B1 => 
                           n12490, B2 => n12484, ZN => n12454);
   U875 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n12327);
   U876 : AOI21_X1 port map( B1 => n12454, B2 => n12327, A => n12326, ZN => 
                           n12383);
   U877 : INV_X1 port map( A => n11723, ZN => n12395);
   U878 : AOI22_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, B1 => 
                           n12383, B2 => n12395, ZN => n12375);
   U879 : OAI21_X1 port map( B1 => n12375, B2 => n12380, A => n12330, ZN => 
                           n12343);
   U880 : XOR2_X1 port map( A => DATA2_I_22_port, B => DATA1(22), Z => n12341);
   U881 : OAI21_X1 port map( B1 => n11724, B2 => n12343, A => n12341, ZN => 
                           n11726);
   U882 : OAI221_X1 port map( B1 => n12346, B2 => n12347, C1 => n12346, C2 => 
                           n11726, A => n11725, ZN => n11727);
   U883 : NOR2_X1 port map( A1 => n13259, A2 => n11727, ZN => n12313);
   U884 : AND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n11729);
   U885 : XOR2_X1 port map( A => DATA2_I_26_port, B => DATA1(26), Z => n12293);
   U886 : NAND2_X1 port map( A1 => n12295, A2 => DATA2_I_25_port, ZN => n12280)
                           ;
   U887 : XOR2_X1 port map( A => DATA2_I_25_port, B => n12295, Z => n12305);
   U888 : NAND3_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, A3 => 
                           n12305, ZN => n12294);
   U889 : NAND2_X1 port map( A1 => n12280, A2 => n12294, ZN => n12277);
   U890 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, B1 => 
                           n12293, B2 => n12277, ZN => n12237);
   U891 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n12250);
   U892 : XOR2_X1 port map( A => DATA2_I_28_port, B => DATA1(28), Z => n12254);
   U893 : OAI21_X1 port map( B1 => DATA1(27), B2 => DATA2_I_27_port, A => 
                           n12254, ZN => n11728);
   U894 : AOI21_X1 port map( B1 => n12237, B2 => n12250, A => n11728, ZN => 
                           n12252);
   U895 : XOR2_X1 port map( A => DATA2_I_29_port, B => DATA1(29), Z => n11731);
   U896 : OAI21_X1 port map( B1 => n11729, B2 => n12252, A => n11731, ZN => 
                           n12066);
   U897 : NAND2_X1 port map( A1 => n11727, A2 => n12927, ZN => n12321);
   U898 : INV_X1 port map( A => n12321, ZN => n12298);
   U899 : INV_X1 port map( A => DATA2_I_24_port, ZN => n12310);
   U900 : NAND2_X1 port map( A1 => n12723, A2 => n12310, ZN => n12322);
   U901 : NAND2_X1 port map( A1 => n12305, A2 => n12322, ZN => n12278);
   U902 : NAND2_X1 port map( A1 => n12280, A2 => n12278, ZN => n12276);
   U903 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, B1 => 
                           n12293, B2 => n12276, ZN => n12238);
   U904 : AOI21_X1 port map( B1 => n12238, B2 => n12250, A => n11728, ZN => 
                           n12251);
   U905 : OAI21_X1 port map( B1 => n11729, B2 => n12251, A => n11731, ZN => 
                           n12065);
   U906 : AOI22_X1 port map( A1 => n12313, A2 => n12066, B1 => n12298, B2 => 
                           n12065, ZN => n12062);
   U907 : NOR2_X1 port map( A1 => n11729, A2 => n11731, ZN => n11732);
   U908 : AOI22_X1 port map( A1 => n12313, A2 => n12252, B1 => n12298, B2 => 
                           n12251, ZN => n11730);
   U909 : OAI22_X1 port map( A1 => n12062, A2 => n11732, B1 => n11731, B2 => 
                           n11730, ZN => n11733);
   U910 : OR3_X1 port map( A1 => n11735, A2 => n11734, A3 => n11733, ZN => 
                           OUTALU(29));
   U911 : INV_X1 port map( A => data1_mul_15_port, ZN => n1976);
   U912 : INV_X1 port map( A => data1_mul_14_port, ZN => n1978);
   U913 : INV_X1 port map( A => data1_mul_13_port, ZN => n1980);
   U914 : INV_X1 port map( A => data1_mul_12_port, ZN => n1982);
   U915 : INV_X1 port map( A => data1_mul_11_port, ZN => n1984);
   U916 : INV_X1 port map( A => data1_mul_10_port, ZN => n1986);
   U917 : INV_X1 port map( A => data1_mul_9_port, ZN => n1988);
   U918 : INV_X1 port map( A => data1_mul_8_port, ZN => n1990);
   U919 : INV_X1 port map( A => data1_mul_7_port, ZN => n1993);
   U920 : INV_X1 port map( A => data1_mul_6_port, ZN => n1998);
   U921 : INV_X1 port map( A => data1_mul_5_port, ZN => n2000);
   U922 : INV_X1 port map( A => data1_mul_4_port, ZN => n2002);
   U923 : INV_X1 port map( A => data1_mul_3_port, ZN => n2004);
   U924 : INV_X1 port map( A => data1_mul_2_port, ZN => n2005);
   U925 : INV_X1 port map( A => data1_mul_1_port, ZN => n2007);
   U926 : XOR2_X1 port map( A => n1976, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => boothmul_pipelined_i_muxes_in_0_119_port);
   U927 : AOI22_X1 port map( A1 => n13235, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n13234, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n11736);
   U928 : OAI21_X1 port map( B1 => n13237, B2 => n1976, A => n11736, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U929 : AOI222_X1 port map( A1 => n11737, A2 => data1_mul_2_port, B1 => 
                           n13235, B2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, C1 => 
                           n13234, C2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n11739);
   U930 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n13005);
   U931 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n13005, ZN => n12965);
   U932 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n12965, ZN => n11738
                           );
   U933 : NOR2_X1 port map( A1 => n11739, A2 => n11738, ZN => n3083);
   U934 : AOI21_X1 port map( B1 => n11739, B2 => n11738, A => n3083, ZN => 
                           n3086);
   U935 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n11740);
   U936 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n11740, ZN => n13007);
   U937 : NOR3_X1 port map( A1 => n5130, A2 => n13007, A3 => n2008, ZN => n3085
                           );
   U938 : OR2_X1 port map( A1 => n2008, A2 => n13007, ZN => n11741);
   U939 : AOI21_X1 port map( B1 => n5130, B2 => n11741, A => n3085, ZN => n3091
                           );
   U940 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n11742);
   U941 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, A
                           => n11742, ZN => n13048);
   U942 : NOR3_X1 port map( A1 => n3077, A2 => n5124, A3 => n13048, ZN => n3084
                           );
   U943 : AOI221_X1 port map( B1 => n3077, B2 => n5124, C1 => n13048, C2 => 
                           n5124, A => n3084, ZN => n3092);
   U944 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n11743);
   U945 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, A
                           => n11743, ZN => n13084);
   U946 : NOR3_X1 port map( A1 => n5121, A2 => n5131, A3 => n13084, ZN => n3090
                           );
   U947 : AOI221_X1 port map( B1 => n5121, B2 => n5131, C1 => n13084, C2 => 
                           n5131, A => n3090, ZN => n3093);
   U948 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n11744);
   U949 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           A => n11744, ZN => n13120);
   U950 : NOR3_X1 port map( A1 => n5122, A2 => n5132, A3 => n13120, ZN => n3089
                           );
   U951 : AOI221_X1 port map( B1 => n5122, B2 => n5132, C1 => n13120, C2 => 
                           n5132, A => n3089, ZN => n3094);
   U952 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n11745);
   U953 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           A => n11745, ZN => n13156);
   U954 : NOR3_X1 port map( A1 => n5123, A2 => n5133, A3 => n13156, ZN => n3088
                           );
   U955 : AOI221_X1 port map( B1 => n5123, B2 => n5133, C1 => n13156, C2 => 
                           n5133, A => n3088, ZN => n3095);
   U956 : INV_X1 port map( A => DATA2(9), ZN => n12950);
   U957 : NAND2_X1 port map( A1 => n12950, A2 => DATA1(9), ZN => n12766);
   U958 : INV_X1 port map( A => n12766, ZN => n12697);
   U959 : NAND2_X1 port map( A1 => n11950, A2 => DATA2(9), ZN => n12699);
   U960 : INV_X1 port map( A => n12699, ZN => n12760);
   U961 : NOR2_X1 port map( A1 => n12697, A2 => n12760, ZN => n12670);
   U962 : INV_X1 port map( A => n12546, ZN => n12649);
   U963 : NOR3_X1 port map( A1 => n12616, A2 => n12950, A3 => n11950, ZN => 
                           n11750);
   U964 : AOI22_X1 port map( A1 => n12117, A2 => n11890, B1 => n12197, B2 => 
                           n11843, ZN => n11748);
   U965 : AOI22_X1 port map( A1 => n12857, A2 => n11926, B1 => n12115, B2 => 
                           n11746, ZN => n11747);
   U966 : AOI21_X1 port map( B1 => n11748, B2 => n11747, A => n12610, ZN => 
                           n11749);
   U967 : AOI211_X1 port map( C1 => dataout_mul_9_port, C2 => n12649, A => 
                           n11750, B => n11749, ZN => n11825);
   U968 : INV_X1 port map( A => n11751, ZN => n11763);
   U969 : AOI22_X1 port map( A1 => n12834, A2 => DATA1(12), B1 => DATA1(16), B2
                           => n11752, ZN => n11756);
   U970 : NAND4_X1 port map( A1 => n11756, A2 => n11755, A3 => n11754, A4 => 
                           n11753, ZN => n11787);
   U971 : AOI222_X1 port map( A1 => n11757, A2 => n12192, B1 => n11787, B2 => 
                           n12267, C1 => n11769, C2 => n12840, ZN => n11834);
   U972 : OAI22_X1 port map( A1 => n12849, A2 => n11834, B1 => n11807, B2 => 
                           n12850, ZN => n11759);
   U973 : OAI22_X1 port map( A1 => n11789, A2 => n12361, B1 => n11764, B2 => 
                           n12026, ZN => n11758);
   U974 : AOI211_X1 port map( C1 => n12030, C2 => n11760, A => n11759, B => 
                           n11758, ZN => n11835);
   U975 : OAI22_X1 port map( A1 => n12860, A2 => n11782, B1 => n12858, B2 => 
                           n11835, ZN => n11762);
   U976 : OAI22_X1 port map( A1 => n12862, A2 => n11810, B1 => n12473, B2 => 
                           n11774, ZN => n11761);
   U977 : AOI211_X1 port map( C1 => n11960, C2 => n11763, A => n11762, B => 
                           n11761, ZN => n11797);
   U978 : INV_X1 port map( A => n11835, ZN => n11796);
   U979 : INV_X1 port map( A => n11764, ZN => n11773);
   U980 : INV_X1 port map( A => DATA1(15), ZN => n12531);
   U981 : OAI211_X1 port map( C1 => n12186, C2 => n12531, A => n11766, B => 
                           n11765, ZN => n11767);
   U982 : AOI211_X1 port map( C1 => DATA1(11), C2 => n12189, A => n11768, B => 
                           n11767, ZN => n11806);
   U983 : INV_X1 port map( A => n11806, ZN => n11770);
   U984 : AOI222_X1 port map( A1 => n12842, A2 => n11770, B1 => n12840, B2 => 
                           n11787, C1 => n12844, C2 => n11769, ZN => n11861);
   U985 : OAI22_X1 port map( A1 => n12849, A2 => n11861, B1 => n11834, B2 => 
                           n12850, ZN => n11772);
   U986 : OAI22_X1 port map( A1 => n11807, A2 => n12361, B1 => n11789, B2 => 
                           n12026, ZN => n11771);
   U987 : AOI211_X1 port map( C1 => n12030, C2 => n11773, A => n11772, B => 
                           n11771, ZN => n11864);
   U988 : OAI22_X1 port map( A1 => n11864, A2 => n12471, B1 => n11810, B2 => 
                           n12860, ZN => n11776);
   U989 : OAI22_X1 port map( A1 => n12865, A2 => n11774, B1 => n11782, B2 => 
                           n12473, ZN => n11775);
   U990 : AOI211_X1 port map( C1 => n12594, C2 => n11796, A => n11776, B => 
                           n11775, ZN => n11814);
   U991 : OAI222_X1 port map( A1 => n12875, A2 => n11797, B1 => n12506, B2 => 
                           n11814, C1 => n11777, C2 => n12870, ZN => n11868);
   U992 : INV_X1 port map( A => n11868, ZN => n11839);
   U993 : OAI222_X1 port map( A1 => n11779, A2 => n12034, B1 => n11778, B2 => 
                           n12875, C1 => n11797, C2 => n12506, ZN => n12574);
   U994 : AOI22_X1 port map( A1 => n12545, A2 => n12574, B1 => n12880, B2 => 
                           n12572, ZN => n11781);
   U995 : AOI22_X1 port map( A1 => n12203, A2 => n12571, B1 => n12879, B2 => 
                           n12575, ZN => n11780);
   U996 : OAI211_X1 port map( C1 => n12514, C2 => n11839, A => n11781, B => 
                           n11780, ZN => n11875);
   U997 : INV_X1 port map( A => n11875, ZN => n12624);
   U998 : OAI22_X1 port map( A1 => n12865, A2 => n11782, B1 => n11810, B2 => 
                           n12473, ZN => n11794);
   U999 : INV_X1 port map( A => n11807, ZN => n11792);
   U1000 : OAI22_X1 port map( A1 => n11834, A2 => n12361, B1 => n11861, B2 => 
                           n12416, ZN => n11791);
   U1001 : OAI211_X1 port map( C1 => n12186, C2 => n12548, A => n11784, B => 
                           n11783, ZN => n11785);
   U1002 : AOI211_X1 port map( C1 => DATA1(10), C2 => n12834, A => n11786, B =>
                           n11785, ZN => n11830);
   U1003 : INV_X1 port map( A => n11787, ZN => n11788);
   U1004 : OAI222_X1 port map( A1 => n12111, A2 => n11806, B1 => n12002, B2 => 
                           n11830, C1 => n11954, C2 => n11788, ZN => n11907);
   U1005 : INV_X1 port map( A => n11907, ZN => n11860);
   U1006 : OAI22_X1 port map( A1 => n12853, A2 => n11789, B1 => n11860, B2 => 
                           n12849, ZN => n11790);
   U1007 : AOI211_X1 port map( C1 => n12857, C2 => n11792, A => n11791, B => 
                           n11790, ZN => n11913);
   U1008 : OAI22_X1 port map( A1 => n11913, A2 => n12471, B1 => n11864, B2 => 
                           n12862, ZN => n11793);
   U1009 : NOR2_X1 port map( A1 => n11794, A2 => n11793, ZN => n11838);
   U1010 : INV_X1 port map( A => n11838, ZN => n11795);
   U1011 : AOI21_X1 port map( B1 => n12569, B2 => n11796, A => n11795, ZN => 
                           n11815);
   U1012 : OAI222_X1 port map( A1 => n11797, A2 => n12034, B1 => n11814, B2 => 
                           n12875, C1 => n11815, C2 => n12506, ZN => n11869);
   U1013 : INV_X1 port map( A => n11869, ZN => n11919);
   U1014 : INV_X1 port map( A => n12574, ZN => n11840);
   U1015 : AOI22_X1 port map( A1 => n12573, A2 => n12575, B1 => n12880, B2 => 
                           n12571, ZN => n11798);
   U1016 : OAI21_X1 port map( B1 => n11840, B2 => n12482, A => n11798, ZN => 
                           n11799);
   U1017 : AOI21_X1 port map( B1 => n12545, B2 => n11868, A => n11799, ZN => 
                           n11901);
   U1018 : OAI21_X1 port map( B1 => n12514, B2 => n11919, A => n11901, ZN => 
                           n11800);
   U1019 : INV_X1 port map( A => n11800, ZN => n12625);
   U1020 : INV_X1 port map( A => n11864, ZN => n11813);
   U1021 : OAI211_X1 port map( C1 => n12105, C2 => n11803, A => n11802, B => 
                           n11801, ZN => n11804);
   U1022 : AOI211_X1 port map( C1 => n13263, C2 => n12408, A => n11805, B => 
                           n11804, ZN => n11858);
   U1023 : OAI222_X1 port map( A1 => n12111, A2 => n11830, B1 => n12002, B2 => 
                           n11858, C1 => n11954, C2 => n11806, ZN => n11955);
   U1024 : INV_X1 port map( A => n11955, ZN => n11910);
   U1025 : OAI22_X1 port map( A1 => n11910, A2 => n12849, B1 => n11861, B2 => 
                           n12361, ZN => n11809);
   U1026 : OAI22_X1 port map( A1 => n12853, A2 => n11807, B1 => n11834, B2 => 
                           n12359, ZN => n11808);
   U1027 : AOI211_X1 port map( C1 => n12197, C2 => n11907, A => n11809, B => 
                           n11808, ZN => n11912);
   U1028 : OAI22_X1 port map( A1 => n11912, A2 => n12471, B1 => n11913, B2 => 
                           n12862, ZN => n11812);
   U1029 : OAI22_X1 port map( A1 => n12865, A2 => n11810, B1 => n11835, B2 => 
                           n12473, ZN => n11811);
   U1030 : AOI211_X1 port map( C1 => n12569, C2 => n11813, A => n11812, B => 
                           n11811, ZN => n11867);
   U1031 : OAI222_X1 port map( A1 => n12875, A2 => n11815, B1 => n12873, B2 => 
                           n11867, C1 => n11814, C2 => n12034, ZN => n11965);
   U1032 : AOI22_X1 port map( A1 => n12573, A2 => n12574, B1 => n12877, B2 => 
                           n11965, ZN => n11817);
   U1033 : AOI22_X1 port map( A1 => n12879, A2 => n11868, B1 => n12880, B2 => 
                           n12575, ZN => n11816);
   U1034 : OAI211_X1 port map( C1 => n11919, C2 => n12495, A => n11817, B => 
                           n11816, ZN => n11970);
   U1035 : INV_X1 port map( A => n11970, ZN => n11922);
   U1036 : OAI222_X1 port map( A1 => n12894, A2 => n12624, B1 => n12623, B2 => 
                           n12625, C1 => n11922, C2 => n12626, ZN => n11823);
   U1037 : AOI211_X1 port map( C1 => n11818, C2 => n11820, A => n12629, B => 
                           n12533, ZN => n11822);
   U1038 : NAND2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => 
                           n11819);
   U1039 : INV_X1 port map( A => n12585, ZN => n12612);
   U1040 : AOI211_X1 port map( C1 => n11820, C2 => n11819, A => n12614, B => 
                           n12612, ZN => n11821);
   U1041 : AOI211_X1 port map( C1 => n12917, C2 => n11823, A => n11822, B => 
                           n11821, ZN => n11824);
   U1042 : OAI211_X1 port map( C1 => n12670, C2 => n12641, A => n11825, B => 
                           n11824, ZN => OUTALU(9));
   U1043 : INV_X1 port map( A => n11852, ZN => n11851);
   U1044 : OAI22_X1 port map( A1 => n11922, A2 => n12623, B1 => n12625, B2 => 
                           n12894, ZN => n11849);
   U1045 : INV_X1 port map( A => n11912, ZN => n11959);
   U1046 : INV_X1 port map( A => n11861, ZN => n11831);
   U1047 : OAI211_X1 port map( C1 => n12186, C2 => n12772, A => n11827, B => 
                           n11826, ZN => n11828);
   U1048 : AOI211_X1 port map( C1 => DATA1(9), C2 => n12408, A => n11829, B => 
                           n11828, ZN => n11906);
   U1049 : OAI222_X1 port map( A1 => n12002, A2 => n11906, B1 => n12111, B2 => 
                           n11858, C1 => n12109, C2 => n11830, ZN => n11982);
   U1050 : AOI22_X1 port map( A1 => n12857, A2 => n11831, B1 => n11982, B2 => 
                           n12080, ZN => n11833);
   U1051 : AOI22_X1 port map( A1 => n12117, A2 => n11907, B1 => n12197, B2 => 
                           n11955, ZN => n11832);
   U1052 : OAI211_X1 port map( C1 => n12853, C2 => n11834, A => n11833, B => 
                           n11832, ZN => n11986);
   U1053 : INV_X1 port map( A => n11986, ZN => n11911);
   U1054 : OAI22_X1 port map( A1 => n11911, A2 => n12858, B1 => n11913, B2 => 
                           n12860, ZN => n11837);
   U1055 : OAI22_X1 port map( A1 => n12865, A2 => n11835, B1 => n11864, B2 => 
                           n12473, ZN => n11836);
   U1056 : AOI211_X1 port map( C1 => n12594, C2 => n11959, A => n11837, B => 
                           n11836, ZN => n11916);
   U1057 : OAI222_X1 port map( A1 => n12875, A2 => n11867, B1 => n12873, B2 => 
                           n11916, C1 => n11838, C2 => n12034, ZN => n11976);
   U1058 : INV_X1 port map( A => n11976, ZN => n11917);
   U1059 : OAI22_X1 port map( A1 => n12514, A2 => n11917, B1 => n11919, B2 => 
                           n12482, ZN => n11842);
   U1060 : OAI22_X1 port map( A1 => n12206, A2 => n11840, B1 => n11839, B2 => 
                           n12886, ZN => n11841);
   U1061 : AOI211_X1 port map( C1 => n12545, C2 => n11965, A => n11842, B => 
                           n11841, ZN => n11993);
   U1062 : OAI22_X1 port map( A1 => n12604, A2 => n11993, B1 => n12624, B2 => 
                           n12436, ZN => n11848);
   U1063 : AOI222_X1 port map( A1 => n11843, A2 => n12080, B1 => n11890, B2 => 
                           n12197, C1 => n11926, C2 => n12117, ZN => n11846);
   U1064 : INV_X1 port map( A => DATA2(8), ZN => n12951);
   U1065 : NAND2_X1 port map( A1 => n12951, A2 => n13262, ZN => n12762);
   U1066 : OAI21_X1 port map( B1 => n12951, B2 => n13262, A => n12762, ZN => 
                           n12671);
   U1067 : AOI22_X1 port map( A1 => dataout_mul_8_port, A2 => n12615, B1 => 
                           n12622, B2 => n12671, ZN => n11845);
   U1068 : NAND3_X1 port map( A1 => DATA2(8), A2 => n13262, A3 => n12580, ZN =>
                           n11844);
   U1069 : OAI211_X1 port map( C1 => n11846, C2 => n12610, A => n11845, B => 
                           n11844, ZN => n11847);
   U1070 : AOI221_X1 port map( B1 => n11849, B2 => n12917, C1 => n11848, C2 => 
                           n12917, A => n11847, ZN => n11850);
   U1071 : OAI221_X1 port map( B1 => n11852, B2 => n12533, C1 => n11851, C2 => 
                           n12612, A => n11850, ZN => OUTALU(8));
   U1072 : AOI22_X1 port map( A1 => DATA1(10), A2 => n11853, B1 => DATA1(11), 
                           B2 => n12017, ZN => n11857);
   U1073 : AND4_X1 port map( A1 => n11857, A2 => n11856, A3 => n11855, A4 => 
                           n11854, ZN => n11953);
   U1074 : OAI222_X1 port map( A1 => n11858, A2 => n12109, B1 => n11953, B2 => 
                           n12002, C1 => n11906, C2 => n12111, ZN => n12029);
   U1075 : INV_X1 port map( A => n12029, ZN => n11859);
   U1076 : OAI22_X1 port map( A1 => n12415, A2 => n11859, B1 => n11910, B2 => 
                           n12361, ZN => n11863);
   U1077 : OAI22_X1 port map( A1 => n12853, A2 => n11861, B1 => n11860, B2 => 
                           n12026, ZN => n11862);
   U1078 : AOI211_X1 port map( C1 => n12197, C2 => n11982, A => n11863, B => 
                           n11862, ZN => n12014);
   U1079 : OAI22_X1 port map( A1 => n12014, A2 => n12471, B1 => n11912, B2 => 
                           n12860, ZN => n11866);
   U1080 : OAI22_X1 port map( A1 => n12865, A2 => n11864, B1 => n11913, B2 => 
                           n12473, ZN => n11865);
   U1081 : AOI211_X1 port map( C1 => n12594, C2 => n11986, A => n11866, B => 
                           n11865, ZN => n11964);
   U1082 : OAI222_X1 port map( A1 => n12875, A2 => n11916, B1 => n12873, B2 => 
                           n11964, C1 => n11867, C2 => n12034, ZN => n12036);
   U1083 : INV_X1 port map( A => n11965, ZN => n11918);
   U1084 : AOI22_X1 port map( A1 => n12573, A2 => n11869, B1 => n12880, B2 => 
                           n11868, ZN => n11870);
   U1085 : OAI21_X1 port map( B1 => n11918, B2 => n12482, A => n11870, ZN => 
                           n11871);
   U1086 : AOI21_X1 port map( B1 => n12541, B2 => n12036, A => n11871, ZN => 
                           n12040);
   U1087 : OAI21_X1 port map( B1 => n12495, B2 => n11917, A => n12040, ZN => 
                           n11872);
   U1088 : INV_X1 port map( A => n11872, ZN => n11994);
   U1089 : OAI22_X1 port map( A1 => n12604, A2 => n11994, B1 => n11993, B2 => 
                           n12623, ZN => n11874);
   U1090 : OAI22_X1 port map( A1 => n11922, A2 => n12894, B1 => n12625, B2 => 
                           n12436, ZN => n11873);
   U1091 : AOI211_X1 port map( C1 => n12829, C2 => n11875, A => n11874, B => 
                           n11873, ZN => n11971);
   U1092 : INV_X1 port map( A => n12439, ZN => n12902);
   U1093 : NAND2_X1 port map( A1 => n12902, A2 => n12917, ZN => n11899);
   U1094 : NOR2_X1 port map( A1 => n13259, A2 => cin, ZN => n12216);
   U1095 : INV_X1 port map( A => n12216, ZN => n12643);
   U1096 : INV_X1 port map( A => n12404, ZN => n12400);
   U1097 : INV_X1 port map( A => n11876, ZN => n11877);
   U1098 : AOI21_X1 port map( B1 => n12401, B2 => n12400, A => n11877, ZN => 
                           n12219);
   U1099 : OAI21_X1 port map( B1 => n12219, B2 => n12230, A => n11878, ZN => 
                           n12046);
   U1100 : AOI21_X1 port map( B1 => n12046, B2 => n12059, A => n11879, ZN => 
                           n12000);
   U1101 : OAI21_X1 port map( B1 => n12000, B2 => n12009, A => n11880, ZN => 
                           n11941);
   U1102 : INV_X1 port map( A => n11943, ZN => n11946);
   U1103 : AOI21_X1 port map( B1 => n11941, B2 => n11946, A => n11881, ZN => 
                           n11884);
   U1104 : NAND2_X1 port map( A1 => n12927, A2 => cin, ZN => n12402);
   U1105 : NOR2_X1 port map( A1 => n11877, A2 => n12403, ZN => n12218);
   U1106 : OAI21_X1 port map( B1 => n12218, B2 => n12230, A => n11878, ZN => 
                           n12045);
   U1107 : AOI21_X1 port map( B1 => n12045, B2 => n12059, A => n11879, ZN => 
                           n11999);
   U1108 : OAI21_X1 port map( B1 => n11999, B2 => n12009, A => n11880, ZN => 
                           n11940);
   U1109 : AOI21_X1 port map( B1 => n11940, B2 => n11946, A => n11881, ZN => 
                           n11888);
   U1110 : OAI22_X1 port map( A1 => n12643, A2 => n11884, B1 => n12402, B2 => 
                           n11888, ZN => n11882);
   U1111 : INV_X1 port map( A => n11882, ZN => n11929);
   U1112 : INV_X1 port map( A => n11885, ZN => n11928);
   U1113 : OAI22_X1 port map( A1 => n11929, A2 => n11928, B1 => n13259, B2 => 
                           n11883, ZN => n11896);
   U1114 : INV_X1 port map( A => n11883, ZN => n11889);
   U1115 : INV_X1 port map( A => n12402, ZN => n12646);
   U1116 : INV_X1 port map( A => n11884, ZN => n11886);
   U1117 : OAI21_X1 port map( B1 => n12643, B2 => n11886, A => n11885, ZN => 
                           n11887);
   U1118 : AOI21_X1 port map( B1 => n12646, B2 => n11888, A => n11887, ZN => 
                           n11927);
   U1119 : NOR4_X1 port map( A1 => n11889, A2 => n11927, A3 => n13259, A4 => 
                           n11897, ZN => n11895);
   U1120 : AOI22_X1 port map( A1 => n12197, A2 => n11926, B1 => n12115, B2 => 
                           n11890, ZN => n11893);
   U1121 : NAND2_X1 port map( A1 => DATA2(7), A2 => n12693, ZN => n12757);
   U1122 : OAI21_X1 port map( B1 => DATA2(7), B2 => n12693, A => n12757, ZN => 
                           n12653);
   U1123 : AOI22_X1 port map( A1 => dataout_mul_7_port, A2 => n12615, B1 => 
                           n12622, B2 => n12653, ZN => n11892);
   U1124 : NAND3_X1 port map( A1 => DATA2(7), A2 => DATA1(7), A3 => n12580, ZN 
                           => n11891);
   U1125 : OAI211_X1 port map( C1 => n11893, C2 => n12610, A => n11892, B => 
                           n11891, ZN => n11894);
   U1126 : AOI211_X1 port map( C1 => n11897, C2 => n11896, A => n11895, B => 
                           n11894, ZN => n11898);
   U1127 : OAI21_X1 port map( B1 => n11971, B2 => n11899, A => n11898, ZN => 
                           OUTALU(7));
   U1128 : INV_X1 port map( A => DATA2(6), ZN => n12955);
   U1129 : NAND2_X1 port map( A1 => DATA1(6), A2 => n12955, ZN => n12692);
   U1130 : OAI221_X1 port map( B1 => DATA1(6), B2 => n12641, C1 => n12691, C2 
                           => n12648, A => n11935, ZN => n11900);
   U1131 : AOI22_X1 port map( A1 => DATA2(6), A2 => n11900, B1 => n12508, B2 =>
                           dataout_mul_6_port, ZN => n11934);
   U1132 : INV_X1 port map( A => n11993, ZN => n11925);
   U1133 : OAI22_X1 port map( A1 => n11994, A2 => n12623, B1 => n11901, B2 => 
                           n12211, ZN => n11924);
   U1134 : INV_X1 port map( A => n12014, ZN => n11958);
   U1135 : AOI22_X1 port map( A1 => DATA1(9), A2 => n12018, B1 => n13263, B2 =>
                           n12017, ZN => n11905);
   U1136 : AND4_X1 port map( A1 => n11905, A2 => n11904, A3 => n11903, A4 => 
                           n11902, ZN => n11981);
   U1137 : OAI222_X1 port map( A1 => n11906, A2 => n12109, B1 => n11981, B2 => 
                           n12113, C1 => n11953, C2 => n12111, ZN => n11947);
   U1138 : AOI22_X1 port map( A1 => n12080, A2 => n11947, B1 => n12029, B2 => 
                           n12197, ZN => n11909);
   U1139 : AOI22_X1 port map( A1 => n11982, A2 => n12117, B1 => n12030, B2 => 
                           n11907, ZN => n11908);
   U1140 : OAI211_X1 port map( C1 => n12359, C2 => n11910, A => n11909, B => 
                           n11908, ZN => n11985);
   U1141 : INV_X1 port map( A => n11985, ZN => n12198);
   U1142 : OAI22_X1 port map( A1 => n11911, A2 => n12860, B1 => n12198, B2 => 
                           n12471, ZN => n11915);
   U1143 : OAI22_X1 port map( A1 => n12865, A2 => n11913, B1 => n11912, B2 => 
                           n12473, ZN => n11914);
   U1144 : AOI211_X1 port map( C1 => n12594, C2 => n11958, A => n11915, B => 
                           n11914, ZN => n11990);
   U1145 : OAI222_X1 port map( A1 => n12875, A2 => n11964, B1 => n12873, B2 => 
                           n11990, C1 => n11916, C2 => n12034, ZN => n12037);
   U1146 : INV_X1 port map( A => n12037, ZN => n12207);
   U1147 : OAI22_X1 port map( A1 => n12514, A2 => n12207, B1 => n11917, B2 => 
                           n12482, ZN => n11921);
   U1148 : OAI22_X1 port map( A1 => n12141, A2 => n11919, B1 => n11918, B2 => 
                           n12886, ZN => n11920);
   U1149 : AOI211_X1 port map( C1 => n12545, C2 => n12036, A => n11921, B => 
                           n11920, ZN => n12212);
   U1150 : OAI22_X1 port map( A1 => n12212, A2 => n12626, B1 => n11922, B2 => 
                           n12436, ZN => n11923);
   U1151 : AOI211_X1 port map( C1 => n12431, C2 => n11925, A => n11924, B => 
                           n11923, ZN => n11997);
   U1152 : OAI22_X1 port map( A1 => n12439, A2 => n11997, B1 => n11971, B2 => 
                           n12896, ZN => n11932);
   U1153 : CLKBUF_X1 port map( A => n12551, Z => n12618);
   U1154 : AND3_X1 port map( A1 => n12115, A2 => n11926, A3 => n12618, ZN => 
                           n11931);
   U1155 : AOI21_X1 port map( B1 => n11929, B2 => n11928, A => n11927, ZN => 
                           n11930);
   U1156 : AOI211_X1 port map( C1 => n12917, C2 => n11932, A => n11931, B => 
                           n11930, ZN => n11933);
   U1157 : OAI211_X1 port map( C1 => n12692, C2 => n12641, A => n11934, B => 
                           n11933, ZN => OUTALU(6));
   U1158 : OAI221_X1 port map( B1 => n13261, B2 => n12641, C1 => n12652, C2 => 
                           n12648, A => n11935, ZN => n11938);
   U1159 : OAI22_X1 port map( A1 => n11936, A2 => n12113, B1 => n12003, B2 => 
                           n12111, ZN => n11937);
   U1160 : AOI22_X1 port map( A1 => DATA2(5), A2 => n11938, B1 => n12618, B2 =>
                           n11937, ZN => n11975);
   U1161 : NAND2_X1 port map( A1 => n12956, A2 => n13261, ZN => n12690);
   U1162 : INV_X1 port map( A => n12690, ZN => n11939);
   U1163 : AOI22_X1 port map( A1 => n11939, A2 => n12622, B1 => n12508, B2 => 
                           dataout_mul_5_port, ZN => n11974);
   U1164 : OAI22_X1 port map( A1 => n12643, A2 => n11941, B1 => n12402, B2 => 
                           n11940, ZN => n11945);
   U1165 : AOI22_X1 port map( A1 => n11941, A2 => n12216, B1 => n11940, B2 => 
                           n12646, ZN => n11942);
   U1166 : INV_X1 port map( A => n11942, ZN => n11944);
   U1167 : AOI22_X1 port map( A1 => n11946, A2 => n11945, B1 => n11944, B2 => 
                           n11943, ZN => n11973);
   U1168 : INV_X1 port map( A => n11947, ZN => n12194);
   U1169 : OAI211_X1 port map( C1 => n12105, C2 => n11950, A => n11949, B => 
                           n11948, ZN => n11951);
   U1170 : AOI211_X1 port map( C1 => n12834, C2 => DATA1(5), A => n11952, B => 
                           n11951, ZN => n12016);
   U1171 : OAI222_X1 port map( A1 => n12002, A2 => n12016, B1 => n12111, B2 => 
                           n11981, C1 => n11954, C2 => n11953, ZN => n12025);
   U1172 : AOI22_X1 port map( A1 => n12117, A2 => n12029, B1 => n12115, B2 => 
                           n12025, ZN => n11957);
   U1173 : AOI22_X1 port map( A1 => n12857, A2 => n11982, B1 => n12030, B2 => 
                           n11955, ZN => n11956);
   U1174 : OAI211_X1 port map( C1 => n12194, C2 => n12850, A => n11957, B => 
                           n11956, ZN => n12015);
   U1175 : AOI22_X1 port map( A1 => n12569, A2 => n11958, B1 => n12617, B2 => 
                           n12015, ZN => n11962);
   U1176 : AOI22_X1 port map( A1 => n12869, A2 => n11986, B1 => n11960, B2 => 
                           n11959, ZN => n11961);
   U1177 : OAI211_X1 port map( C1 => n12198, C2 => n12862, A => n11962, B => 
                           n11961, ZN => n11963);
   U1178 : INV_X1 port map( A => n11963, ZN => n12035);
   U1179 : OAI222_X1 port map( A1 => n11964, A2 => n12870, B1 => n11990, B2 => 
                           n12875, C1 => n12035, C2 => n12506, ZN => n12427);
   U1180 : AOI22_X1 port map( A1 => n12879, A2 => n12036, B1 => n12541, B2 => 
                           n12427, ZN => n11967);
   U1181 : AOI22_X1 port map( A1 => n12203, A2 => n11976, B1 => n12880, B2 => 
                           n11965, ZN => n11966);
   U1182 : OAI211_X1 port map( C1 => n12207, C2 => n12495, A => n11967, B => 
                           n11966, ZN => n12432);
   U1183 : INV_X1 port map( A => n12432, ZN => n12041);
   U1184 : OAI22_X1 port map( A1 => n12041, A2 => n12626, B1 => n11994, B2 => 
                           n12894, ZN => n11969);
   U1185 : OAI22_X1 port map( A1 => n12212, A2 => n12623, B1 => n11993, B2 => 
                           n12436, ZN => n11968);
   U1186 : AOI211_X1 port map( C1 => n12829, C2 => n11970, A => n11969, B => 
                           n11968, ZN => n12044);
   U1187 : OAI222_X1 port map( A1 => n12896, A2 => n11997, B1 => n12215, B2 => 
                           n11971, C1 => n12044, C2 => n12213, ZN => n12443);
   U1188 : NAND3_X1 port map( A1 => n12917, A2 => n12442, A3 => n12443, ZN => 
                           n11972);
   U1189 : NAND4_X1 port map( A1 => n11975, A2 => n11974, A3 => n11973, A4 => 
                           n11972, ZN => OUTALU(5));
   U1190 : AOI22_X1 port map( A1 => n12203, A2 => n12036, B1 => n12880, B2 => 
                           n11976, ZN => n11992);
   U1191 : OAI211_X1 port map( C1 => n12186, C2 => n12696, A => n11978, B => 
                           n11977, ZN => n11979);
   U1192 : AOI211_X1 port map( C1 => n13261, C2 => n12835, A => n11980, B => 
                           n11979, ZN => n12023);
   U1193 : OAI222_X1 port map( A1 => n12002, A2 => n12023, B1 => n12111, B2 => 
                           n12016, C1 => n12109, C2 => n11981, ZN => n12420);
   U1194 : AOI22_X1 port map( A1 => n12857, A2 => n12029, B1 => n12115, B2 => 
                           n12420, ZN => n11984);
   U1195 : AOI22_X1 port map( A1 => n12197, A2 => n12025, B1 => n12030, B2 => 
                           n11982, ZN => n11983);
   U1196 : OAI211_X1 port map( C1 => n12194, C2 => n12361, A => n11984, B => 
                           n11983, ZN => n12424);
   U1197 : AOI22_X1 port map( A1 => n12617, A2 => n12424, B1 => n12569, B2 => 
                           n11985, ZN => n11988);
   U1198 : AOI22_X1 port map( A1 => n12594, A2 => n12015, B1 => n11986, B2 => 
                           n12128, ZN => n11987);
   U1199 : OAI211_X1 port map( C1 => n12014, C2 => n12473, A => n11988, B => 
                           n11987, ZN => n11989);
   U1200 : INV_X1 port map( A => n11989, ZN => n12202);
   U1201 : OAI222_X1 port map( A1 => n11990, A2 => n12870, B1 => n12035, B2 => 
                           n12875, C1 => n12202, C2 => n12506, ZN => n12881);
   U1202 : AOI22_X1 port map( A1 => n12879, A2 => n12037, B1 => n12877, B2 => 
                           n12881, ZN => n11991);
   U1203 : NAND2_X1 port map( A1 => n11992, A2 => n11991, ZN => n12828);
   U1204 : AOI21_X1 port map( B1 => n12545, B2 => n12427, A => n12828, ZN => 
                           n12437);
   U1205 : OAI22_X1 port map( A1 => n12437, A2 => n12626, B1 => n11993, B2 => 
                           n12211, ZN => n11996);
   U1206 : OAI22_X1 port map( A1 => n12212, A2 => n12894, B1 => n11994, B2 => 
                           n12436, ZN => n11995);
   U1207 : AOI211_X1 port map( C1 => n12831, C2 => n12432, A => n11996, B => 
                           n11995, ZN => n12214);
   U1208 : OAI222_X1 port map( A1 => n12896, A2 => n12044, B1 => n12897, B2 => 
                           n11997, C1 => n12214, C2 => n12213, ZN => n12910);
   U1209 : AOI22_X1 port map( A1 => n12442, A2 => n12910, B1 => n12907, B2 => 
                           n12443, ZN => n12013);
   U1210 : INV_X1 port map( A => n12009, ZN => n12011);
   U1211 : AOI22_X1 port map( A1 => n12216, A2 => n12000, B1 => n12646, B2 => 
                           n11999, ZN => n11998);
   U1212 : INV_X1 port map( A => n11998, ZN => n12010);
   U1213 : OAI22_X1 port map( A1 => n12000, A2 => n12643, B1 => n11999, B2 => 
                           n12402, ZN => n12008);
   U1214 : NAND2_X1 port map( A1 => n12957, A2 => DATA1(4), ZN => n12685);
   U1215 : NOR2_X1 port map( A1 => n12957, A2 => DATA1(4), ZN => n12748);
   U1216 : INV_X1 port map( A => n12748, ZN => n12688);
   U1217 : NOR3_X1 port map( A1 => n12616, A2 => n12001, A3 => n12957, ZN => 
                           n12005);
   U1218 : NOR3_X1 port map( A1 => n12003, A2 => n12610, A3 => n12002, ZN => 
                           n12004);
   U1219 : AOI211_X1 port map( C1 => dataout_mul_4_port, C2 => n12615, A => 
                           n12005, B => n12004, ZN => n12006);
   U1220 : OAI221_X1 port map( B1 => n12641, B2 => n12685, C1 => n12641, C2 => 
                           n12688, A => n12006, ZN => n12007);
   U1221 : AOI221_X1 port map( B1 => n12011, B2 => n12010, C1 => n12009, C2 => 
                           n12008, A => n12007, ZN => n12012);
   U1222 : OAI21_X1 port map( B1 => n12013, B2 => n12603, A => n12012, ZN => 
                           OUTALU(4));
   U1223 : INV_X1 port map( A => n12881, ZN => n12430);
   U1224 : INV_X1 port map( A => n12424, ZN => n12864);
   U1225 : OAI22_X1 port map( A1 => n12865, A2 => n12014, B1 => n12198, B2 => 
                           n12473, ZN => n12032);
   U1226 : INV_X1 port map( A => n12015, ZN => n12421);
   U1227 : INV_X1 port map( A => n12016, ZN => n12024);
   U1228 : AOI22_X1 port map( A1 => DATA1(6), A2 => n12018, B1 => DATA1(7), B2 
                           => n12017, ZN => n12022);
   U1229 : INV_X1 port map( A => n12019, ZN => n12021);
   U1230 : NAND2_X1 port map( A1 => n12189, A2 => DATA1(3), ZN => n12048);
   U1231 : NAND4_X1 port map( A1 => n12022, A2 => n12021, A3 => n12020, A4 => 
                           n12048, ZN => n12413);
   U1232 : INV_X1 port map( A => n12023, ZN => n12191);
   U1233 : AOI222_X1 port map( A1 => n12024, A2 => n12844, B1 => n12413, B2 => 
                           n12267, C1 => n12191, C2 => n12840, ZN => n12414);
   U1234 : INV_X1 port map( A => n12025, ZN => n12417);
   U1235 : OAI22_X1 port map( A1 => n12415, A2 => n12414, B1 => n12417, B2 => 
                           n12361, ZN => n12028);
   U1236 : INV_X1 port map( A => n12420, ZN => n12852);
   U1237 : OAI22_X1 port map( A1 => n12194, A2 => n12026, B1 => n12852, B2 => 
                           n12416, ZN => n12027);
   U1238 : AOI211_X1 port map( C1 => n12030, C2 => n12029, A => n12028, B => 
                           n12027, ZN => n12833);
   U1239 : OAI22_X1 port map( A1 => n12421, A2 => n12860, B1 => n12833, B2 => 
                           n12858, ZN => n12031);
   U1240 : NOR2_X1 port map( A1 => n12032, A2 => n12031, ZN => n12426);
   U1241 : OAI21_X1 port map( B1 => n12864, B2 => n12862, A => n12426, ZN => 
                           n12033);
   U1242 : INV_X1 port map( A => n12033, ZN => n12201);
   U1243 : OAI222_X1 port map( A1 => n12035, A2 => n12034, B1 => n12202, B2 => 
                           n12875, C1 => n12201, C2 => n12506, ZN => n12832);
   U1244 : AOI22_X1 port map( A1 => n12879, A2 => n12427, B1 => n12877, B2 => 
                           n12832, ZN => n12039);
   U1245 : AOI22_X1 port map( A1 => n12203, A2 => n12037, B1 => n12880, B2 => 
                           n12036, ZN => n12038);
   U1246 : OAI211_X1 port map( C1 => n12430, C2 => n12495, A => n12039, B => 
                           n12038, ZN => n12890);
   U1247 : OAI22_X1 port map( A1 => n12437, A2 => n12623, B1 => n12040, B2 => 
                           n12211, ZN => n12043);
   U1248 : OAI22_X1 port map( A1 => n12041, A2 => n12894, B1 => n12212, B2 => 
                           n12436, ZN => n12042);
   U1249 : AOI211_X1 port map( C1 => n12890, C2 => n12889, A => n12043, B => 
                           n12042, ZN => n12440);
   U1250 : OAI222_X1 port map( A1 => n12896, A2 => n12214, B1 => n12897, B2 => 
                           n12044, C1 => n12440, C2 => n12213, ZN => n12908);
   U1251 : AOI222_X1 port map( A1 => n12908, A2 => n12442, B1 => n12443, B2 => 
                           n12905, C1 => n12910, C2 => n12907, ZN => n12061);
   U1252 : OAI22_X1 port map( A1 => n12643, A2 => n12046, B1 => n12402, B2 => 
                           n12045, ZN => n12058);
   U1253 : INV_X1 port map( A => n12059, ZN => n12057);
   U1254 : AOI22_X1 port map( A1 => n12046, A2 => n12216, B1 => n12045, B2 => 
                           n12646, ZN => n12047);
   U1255 : INV_X1 port map( A => n12047, ZN => n12056);
   U1256 : NAND2_X1 port map( A1 => n12408, A2 => DATA1(2), ZN => n12049);
   U1257 : OAI211_X1 port map( C1 => n12240, C2 => n12640, A => n12049, B => 
                           n12048, ZN => n12050);
   U1258 : AOI21_X1 port map( B1 => n12223, B2 => n12398, A => n12050, ZN => 
                           n12054);
   U1259 : NOR2_X1 port map( A1 => n12958, A2 => DATA1(3), ZN => n12749);
   U1260 : INV_X1 port map( A => n12749, ZN => n12051);
   U1261 : NAND2_X1 port map( A1 => DATA1(3), A2 => n12958, ZN => n12750);
   U1262 : NAND2_X1 port map( A1 => n12051, A2 => n12750, ZN => n12655);
   U1263 : AOI22_X1 port map( A1 => dataout_mul_3_port, A2 => n12615, B1 => 
                           n12622, B2 => n12655, ZN => n12053);
   U1264 : NAND3_X1 port map( A1 => DATA1(3), A2 => DATA2(3), A3 => n12580, ZN 
                           => n12052);
   U1265 : OAI211_X1 port map( C1 => n12054, C2 => n12610, A => n12053, B => 
                           n12052, ZN => n12055);
   U1266 : AOI221_X1 port map( B1 => n12059, B2 => n12058, C1 => n12057, C2 => 
                           n12056, A => n12055, ZN => n12060);
   U1267 : OAI21_X1 port map( B1 => n12061, B2 => n12603, A => n12060, ZN => 
                           OUTALU(3));
   U1268 : INV_X1 port map( A => DATA2(31), ZN => n12928);
   U1269 : NAND2_X1 port map( A1 => n12928, A2 => DATA1(31), ZN => n12827);
   U1270 : INV_X1 port map( A => n12827, ZN => n12733);
   U1271 : INV_X1 port map( A => DATA1(31), ZN => n12239);
   U1272 : NAND2_X1 port map( A1 => n12239, A2 => DATA2(31), ZN => n12824);
   U1273 : INV_X1 port map( A => n12824, ZN => n12736);
   U1274 : NOR2_X1 port map( A1 => n12733, A2 => n12736, ZN => n12678);
   U1275 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n12063);
   U1276 : AND2_X1 port map( A1 => DATA1(29), A2 => DATA2_I_29_port, ZN => 
                           n12178);
   U1277 : XOR2_X1 port map( A => DATA2_I_30_port, B => DATA1(30), Z => n12182)
                           ;
   U1278 : OAI22_X1 port map( A1 => n12178, A2 => n12062, B1 => n12182, B2 => 
                           n13259, ZN => n12177);
   U1279 : NAND2_X1 port map( A1 => n12063, A2 => n12177, ZN => n12156);
   U1280 : INV_X1 port map( A => DATA2_I_31_port, ZN => n12157);
   U1281 : AOI22_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, B1 => 
                           n12178, B2 => n12182, ZN => n12064);
   U1282 : INV_X1 port map( A => n12064, ZN => n12067);
   U1283 : INV_X1 port map( A => n12313, ZN => n12262);
   U1284 : OAI22_X1 port map( A1 => n12262, A2 => n12066, B1 => n12321, B2 => 
                           n12065, ZN => n12170);
   U1285 : AOI22_X1 port map( A1 => n12067, A2 => n12927, B1 => n12170, B2 => 
                           n12182, ZN => n12158);
   U1286 : OAI22_X1 port map( A1 => n12928, A2 => n12616, B1 => n12157, B2 => 
                           n12158, ZN => n12068);
   U1287 : INV_X1 port map( A => n12068, ZN => n12069);
   U1288 : NAND2_X1 port map( A1 => n12834, A2 => n12917, ZN => n12171);
   U1289 : OAI211_X1 port map( C1 => DATA2_I_31_port, C2 => n12156, A => n12069
                           , B => n12171, ZN => n12070);
   U1290 : AOI22_X1 port map( A1 => DATA1(31), A2 => n12070, B1 => n12508, B2 
                           => dataout_mul_31_port, ZN => n12169);
   U1291 : INV_X1 port map( A => n12071, ZN => n12149);
   U1292 : INV_X1 port map( A => n12072, ZN => n12145);
   U1293 : INV_X1 port map( A => DATA1(26), ZN => n12283);
   U1294 : NOR2_X1 port map( A1 => n12396, A2 => n12073, ZN => n12243);
   U1295 : AOI211_X1 port map( C1 => n12834, C2 => DATA1(30), A => n12074, B =>
                           n12243, ZN => n12076);
   U1296 : OAI211_X1 port map( C1 => n12186, C2 => n12283, A => n12076, B => 
                           n12075, ZN => n12077);
   U1297 : INV_X1 port map( A => n12077, ZN => n12110);
   U1298 : OAI222_X1 port map( A1 => n12078, A2 => n12109, B1 => n12110, B2 => 
                           n12113, C1 => n12108, C2 => n12111, ZN => n12120);
   U1299 : AOI22_X1 port map( A1 => n12080, A2 => n12120, B1 => n12079, B2 => 
                           n12117, ZN => n12082);
   U1300 : AOI22_X1 port map( A1 => n12118, A2 => n12857, B1 => n12116, B2 => 
                           n12197, ZN => n12081);
   U1301 : OAI211_X1 port map( C1 => n12853, C2 => n12083, A => n12082, B => 
                           n12081, ZN => n12102);
   U1302 : AOI22_X1 port map( A1 => n12129, A2 => n12126, B1 => n12102, B2 => 
                           n12617, ZN => n12086);
   U1303 : AOI22_X1 port map( A1 => n12128, A2 => n12084, B1 => n12125, B2 => 
                           n12594, ZN => n12085);
   U1304 : OAI211_X1 port map( C1 => n12473, C2 => n12087, A => n12086, B => 
                           n12085, ZN => n12134);
   U1305 : AOI222_X1 port map( A1 => n12526, A2 => n12136, B1 => n12550, B2 => 
                           n12134, C1 => n12088, C2 => n12135, ZN => n12101);
   U1306 : OAI22_X1 port map( A1 => n12482, A2 => n12139, B1 => n12514, B2 => 
                           n12101, ZN => n12091);
   U1307 : OAI22_X1 port map( A1 => n12886, A2 => n12140, B1 => n12206, B2 => 
                           n12089, ZN => n12090);
   U1308 : AOI211_X1 port map( C1 => n12092, C2 => n12545, A => n12091, B => 
                           n12090, ZN => n12099);
   U1309 : OAI22_X1 port map( A1 => n12436, A2 => n12145, B1 => n12626, B2 => 
                           n12099, ZN => n12096);
   U1310 : INV_X1 port map( A => n12093, ZN => n12100);
   U1311 : OAI22_X1 port map( A1 => n12623, A2 => n12100, B1 => n12211, B2 => 
                           n12094, ZN => n12095);
   U1312 : AOI211_X1 port map( C1 => n12149, C2 => n12431, A => n12096, B => 
                           n12095, ZN => n12152);
   U1313 : OAI222_X1 port map( A1 => n12152, A2 => n12213, B1 => n12151, B2 => 
                           n12896, C1 => n12097, C2 => n12215, ZN => n12098);
   U1314 : INV_X1 port map( A => n12098, ZN => n12164);
   U1315 : OAI22_X1 port map( A1 => n12100, A2 => n12894, B1 => n12099, B2 => 
                           n12623, ZN => n12148);
   U1316 : INV_X1 port map( A => n12101, ZN => n12144);
   U1317 : INV_X1 port map( A => n12102, ZN => n12132);
   U1318 : INV_X1 port map( A => DATA1(27), ZN => n12264);
   U1319 : OAI211_X1 port map( C1 => n12105, C2 => n12264, A => n12104, B => 
                           n12103, ZN => n12106);
   U1320 : AOI211_X1 port map( C1 => DATA1(31), C2 => n12189, A => n12107, B =>
                           n12106, ZN => n12112);
   U1321 : OAI222_X1 port map( A1 => n12113, A2 => n12112, B1 => n12111, B2 => 
                           n12110, C1 => n12109, C2 => n12108, ZN => n12114);
   U1322 : AOI22_X1 port map( A1 => n12117, A2 => n12116, B1 => n12115, B2 => 
                           n12114, ZN => n12122);
   U1323 : AOI22_X1 port map( A1 => n12197, A2 => n12120, B1 => n12119, B2 => 
                           n12118, ZN => n12121);
   U1324 : OAI211_X1 port map( C1 => n12123, C2 => n12359, A => n12122, B => 
                           n12121, ZN => n12124);
   U1325 : AOI22_X1 port map( A1 => n12126, A2 => n12125, B1 => n12617, B2 => 
                           n12124, ZN => n12131);
   U1326 : AOI22_X1 port map( A1 => n12425, A2 => n12129, B1 => n12128, B2 => 
                           n12127, ZN => n12130);
   U1327 : OAI211_X1 port map( C1 => n12132, C2 => n12862, A => n12131, B => 
                           n12130, ZN => n12133);
   U1328 : AOI222_X1 port map( A1 => n12136, A2 => n12135, B1 => n12134, B2 => 
                           n12526, C1 => n12133, C2 => n12550, ZN => n12138);
   U1329 : OAI22_X1 port map( A1 => n12514, A2 => n12138, B1 => n12137, B2 => 
                           n12482, ZN => n12143);
   U1330 : OAI22_X1 port map( A1 => n12141, A2 => n12140, B1 => n12139, B2 => 
                           n12886, ZN => n12142);
   U1331 : AOI211_X1 port map( C1 => n12545, C2 => n12144, A => n12143, B => 
                           n12142, ZN => n12146);
   U1332 : OAI22_X1 port map( A1 => n12604, A2 => n12146, B1 => n12145, B2 => 
                           n12211, ZN => n12147);
   U1333 : AOI211_X1 port map( C1 => n12891, C2 => n12149, A => n12148, B => 
                           n12147, ZN => n12150);
   U1334 : OAI222_X1 port map( A1 => n12896, A2 => n12152, B1 => n12897, B2 => 
                           n12151, C1 => n12150, C2 => n12213, ZN => n12153);
   U1335 : AOI22_X1 port map( A1 => n12442, A2 => n12153, B1 => n12911, B2 => 
                           n12263, ZN => n12155);
   U1336 : AOI22_X1 port map( A1 => n12909, A2 => n12236, B1 => n12905, B2 => 
                           n12161, ZN => n12154);
   U1337 : OAI211_X1 port map( C1 => n12164, C2 => n12446, A => n12155, B => 
                           n12154, ZN => n12167);
   U1338 : AOI221_X1 port map( B1 => n12158, B2 => n12157, C1 => n12156, C2 => 
                           DATA2_I_31_port, A => DATA1(31), ZN => n12166);
   U1339 : NOR2_X1 port map( A1 => n12160, A2 => n12159, ZN => n12921);
   U1340 : AOI22_X1 port map( A1 => n12909, A2 => n12263, B1 => n12907, B2 => 
                           n12161, ZN => n12163);
   U1341 : AOI22_X1 port map( A1 => n12911, A2 => n12289, B1 => n12905, B2 => 
                           n12236, ZN => n12162);
   U1342 : OAI211_X1 port map( C1 => n12164, C2 => n12914, A => n12163, B => 
                           n12162, ZN => n12176);
   U1343 : AND3_X1 port map( A1 => n12921, A2 => n12926, A3 => n12176, ZN => 
                           n12165);
   U1344 : AOI211_X1 port map( C1 => n12551, C2 => n12167, A => n12166, B => 
                           n12165, ZN => n12168);
   U1345 : OAI211_X1 port map( C1 => n12678, C2 => n12641, A => n12169, B => 
                           n12168, ZN => OUTALU(31));
   U1346 : INV_X1 port map( A => n12170, ZN => n12181);
   U1347 : INV_X1 port map( A => DATA2(30), ZN => n12929);
   U1348 : OAI22_X1 port map( A1 => n12825, A2 => DATA2(30), B1 => n12929, B2 
                           => DATA1(30), ZN => n12730);
   U1349 : INV_X1 port map( A => n12730, ZN => n12820);
   U1350 : OAI21_X1 port map( B1 => n12616, B2 => n12929, A => n12171, ZN => 
                           n12172);
   U1351 : AOI22_X1 port map( A1 => DATA1(30), A2 => n12172, B1 => n12508, B2 
                           => dataout_mul_30_port, ZN => n12174);
   U1352 : NAND3_X1 port map( A1 => n12835, A2 => n12917, A3 => DATA1(31), ZN 
                           => n12173);
   U1353 : OAI211_X1 port map( C1 => n12820, C2 => n12641, A => n12174, B => 
                           n12173, ZN => n12175);
   U1354 : AOI21_X1 port map( B1 => n12618, B2 => n12176, A => n12175, ZN => 
                           n12180);
   U1355 : OAI21_X1 port map( B1 => n12178, B2 => n12182, A => n12177, ZN => 
                           n12179);
   U1356 : OAI211_X1 port map( C1 => n12182, C2 => n12181, A => n12180, B => 
                           n12179, ZN => OUTALU(30));
   U1357 : AOI22_X1 port map( A1 => n12905, A2 => n12910, B1 => n12907, B2 => 
                           n12908, ZN => n12235);
   U1358 : AOI22_X1 port map( A1 => n12881, A2 => n12879, B1 => n12832, B2 => 
                           n12545, ZN => n12205);
   U1359 : INV_X1 port map( A => n12414, ZN => n12856);
   U1360 : INV_X1 port map( A => n12183, ZN => n12184);
   U1361 : OAI211_X1 port map( C1 => n12186, C2 => n12691, A => n12185, B => 
                           n12184, ZN => n12187);
   U1362 : AOI211_X1 port map( C1 => n12189, C2 => DATA1(2), A => n12188, B => 
                           n12187, ZN => n12190);
   U1363 : INV_X1 port map( A => n12190, ZN => n12845);
   U1364 : AOI222_X1 port map( A1 => n12842, A2 => n12845, B1 => n12193, B2 => 
                           n12413, C1 => n12192, C2 => n12191, ZN => n12847);
   U1365 : OAI22_X1 port map( A1 => n12846, A2 => n12852, B1 => n12849, B2 => 
                           n12847, ZN => n12196);
   U1366 : OAI22_X1 port map( A1 => n12359, A2 => n12417, B1 => n12853, B2 => 
                           n12194, ZN => n12195);
   U1367 : AOI211_X1 port map( C1 => n12856, C2 => n12197, A => n12196, B => 
                           n12195, ZN => n12861);
   U1368 : OAI22_X1 port map( A1 => n12473, A2 => n12421, B1 => n12858, B2 => 
                           n12861, ZN => n12200);
   U1369 : OAI22_X1 port map( A1 => n12862, A2 => n12833, B1 => n12198, B2 => 
                           n12865, ZN => n12199);
   U1370 : AOI211_X1 port map( C1 => n12424, C2 => n12569, A => n12200, B => 
                           n12199, ZN => n12871);
   U1371 : OAI222_X1 port map( A1 => n12202, A2 => n12870, B1 => n12201, B2 => 
                           n12875, C1 => n12871, C2 => n12506, ZN => n12878);
   U1372 : AOI22_X1 port map( A1 => n12541, A2 => n12878, B1 => n12427, B2 => 
                           n12203, ZN => n12204);
   U1373 : OAI211_X1 port map( C1 => n12207, C2 => n12206, A => n12205, B => 
                           n12204, ZN => n12433);
   U1374 : INV_X1 port map( A => n12433, ZN => n12895);
   U1375 : OAI22_X1 port map( A1 => n12894, A2 => n12437, B1 => n12626, B2 => 
                           n12895, ZN => n12208);
   U1376 : INV_X1 port map( A => n12208, ZN => n12210);
   U1377 : AOI22_X1 port map( A1 => n12831, A2 => n12890, B1 => n12891, B2 => 
                           n12432, ZN => n12209);
   U1378 : OAI211_X1 port map( C1 => n12212, C2 => n12211, A => n12210, B => 
                           n12209, ZN => n12899);
   U1379 : INV_X1 port map( A => n12899, ZN => n12441);
   U1380 : OAI222_X1 port map( A1 => n12896, A2 => n12440, B1 => n12215, B2 => 
                           n12214, C1 => n12213, C2 => n12441, ZN => n12904);
   U1381 : AOI22_X1 port map( A1 => n12442, A2 => n12904, B1 => n12909, B2 => 
                           n12443, ZN => n12234);
   U1382 : INV_X1 port map( A => n12230, ZN => n12232);
   U1383 : AOI22_X1 port map( A1 => n12216, A2 => n12219, B1 => n12646, B2 => 
                           n12218, ZN => n12217);
   U1384 : INV_X1 port map( A => n12217, ZN => n12231);
   U1385 : OAI22_X1 port map( A1 => n12219, A2 => n12643, B1 => n12218, B2 => 
                           n12402, ZN => n12229);
   U1386 : NOR2_X1 port map( A1 => n12220, A2 => n12224, ZN => n12222);
   U1387 : AND2_X1 port map( A1 => n12408, A2 => n12398, ZN => n12221);
   U1388 : AOI211_X1 port map( C1 => n12223, C2 => DATA1(0), A => n12222, B => 
                           n12221, ZN => n12227);
   U1389 : OAI22_X1 port map( A1 => n12959, A2 => DATA1(2), B1 => n12224, B2 =>
                           DATA2(2), ZN => n12742);
   U1390 : AOI22_X1 port map( A1 => dataout_mul_2_port, A2 => n12615, B1 => 
                           n12622, B2 => n12742, ZN => n12226);
   U1391 : NAND3_X1 port map( A1 => n13260, A2 => DATA2(2), A3 => n12580, ZN =>
                           n12225);
   U1392 : OAI211_X1 port map( C1 => n12227, C2 => n12610, A => n12226, B => 
                           n12225, ZN => n12228);
   U1393 : AOI221_X1 port map( B1 => n12232, B2 => n12231, C1 => n12230, C2 => 
                           n12229, A => n12228, ZN => n12233);
   U1394 : OAI221_X1 port map( B1 => n12603, B2 => n12235, C1 => n12603, C2 => 
                           n12234, A => n12233, ZN => OUTALU(2));
   U1395 : AOI222_X1 port map( A1 => n12236, A2 => n12442, B1 => n12289, B2 => 
                           n12905, C1 => n12263, C2 => n12907, ZN => n12257);
   U1396 : NOR2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n12258);
   U1397 : INV_X1 port map( A => n12237, ZN => n12261);
   U1398 : INV_X1 port map( A => n12238, ZN => n12260);
   U1399 : AOI22_X1 port map( A1 => n12313, A2 => n12261, B1 => n12298, B2 => 
                           n12260, ZN => n12275);
   U1400 : NOR3_X1 port map( A1 => n12258, A2 => n12254, A3 => n12275, ZN => 
                           n12249);
   U1401 : OAI22_X1 port map( A1 => n12241, A2 => n12825, B1 => n12240, B2 => 
                           n12239, ZN => n12242);
   U1402 : AOI211_X1 port map( C1 => DATA1(28), C2 => n12834, A => n12243, B =>
                           n12242, ZN => n12247);
   U1403 : NOR2_X1 port map( A1 => DATA2(28), A2 => n12244, ZN => n12822);
   U1404 : INV_X1 port map( A => DATA2(28), ZN => n12931);
   U1405 : NOR2_X1 port map( A1 => n12931, A2 => DATA1(28), ZN => n12727);
   U1406 : OAI21_X1 port map( B1 => n12822, B2 => n12727, A => n12622, ZN => 
                           n12246);
   U1407 : NAND3_X1 port map( A1 => DATA2(28), A2 => DATA1(28), A3 => n12580, 
                           ZN => n12245);
   U1408 : OAI211_X1 port map( C1 => n12247, C2 => n12603, A => n12246, B => 
                           n12245, ZN => n12248);
   U1409 : AOI211_X1 port map( C1 => n12649, C2 => dataout_mul_28_port, A => 
                           n12249, B => n12248, ZN => n12256);
   U1410 : INV_X1 port map( A => n12250, ZN => n12259);
   U1411 : OAI22_X1 port map( A1 => n12252, A2 => n12262, B1 => n12251, B2 => 
                           n12321, ZN => n12253);
   U1412 : OAI21_X1 port map( B1 => n12259, B2 => n12254, A => n12253, ZN => 
                           n12255);
   U1413 : OAI211_X1 port map( C1 => n12257, C2 => n12610, A => n12256, B => 
                           n12255, ZN => OUTALU(28));
   U1414 : NOR2_X1 port map( A1 => n12259, A2 => n12258, ZN => n12274);
   U1415 : OAI22_X1 port map( A1 => n12262, A2 => n12261, B1 => n12321, B2 => 
                           n12260, ZN => n12272);
   U1416 : AOI22_X1 port map( A1 => n12442, A2 => n12263, B1 => n12907, B2 => 
                           n12289, ZN => n12270);
   U1417 : INV_X1 port map( A => DATA2(27), ZN => n12932);
   U1418 : NAND2_X1 port map( A1 => n12932, A2 => DATA1(27), ZN => n12668);
   U1419 : NAND2_X1 port map( A1 => DATA2(27), A2 => n12264, ZN => n12815);
   U1420 : AOI21_X1 port map( B1 => n12668, B2 => n12815, A => n12641, ZN => 
                           n12266);
   U1421 : NOR3_X1 port map( A1 => n12616, A2 => n12932, A3 => n12264, ZN => 
                           n12265);
   U1422 : AOI211_X1 port map( C1 => n12649, C2 => dataout_mul_27_port, A => 
                           n12266, B => n12265, ZN => n12269);
   U1423 : NAND3_X1 port map( A1 => n12917, A2 => n12267, A3 => n12281, ZN => 
                           n12268);
   U1424 : OAI211_X1 port map( C1 => n12270, C2 => n12610, A => n12269, B => 
                           n12268, ZN => n12271);
   U1425 : AOI21_X1 port map( B1 => n12274, B2 => n12272, A => n12271, ZN => 
                           n12273);
   U1426 : OAI21_X1 port map( B1 => n12275, B2 => n12274, A => n12273, ZN => 
                           OUTALU(27));
   U1427 : AOI22_X1 port map( A1 => n12313, A2 => n12277, B1 => n12298, B2 => 
                           n12276, ZN => n12292);
   U1428 : AOI22_X1 port map( A1 => n12313, A2 => n12294, B1 => n12298, B2 => 
                           n12278, ZN => n12279);
   U1429 : INV_X1 port map( A => n12279, ZN => n12304);
   U1430 : AND2_X1 port map( A1 => n12280, A2 => n12304, ZN => n12288);
   U1431 : AOI22_X1 port map( A1 => n12842, A2 => n12282, B1 => n12840, B2 => 
                           n12281, ZN => n12286);
   U1432 : NOR2_X1 port map( A1 => n12283, A2 => DATA2(26), ZN => n12810);
   U1433 : INV_X1 port map( A => n12810, ZN => n12724);
   U1434 : NAND2_X1 port map( A1 => DATA2(26), A2 => n12283, ZN => n12813);
   U1435 : NAND2_X1 port map( A1 => n12724, A2 => n12813, ZN => n12654);
   U1436 : AOI22_X1 port map( A1 => dataout_mul_26_port, A2 => n12615, B1 => 
                           n12622, B2 => n12654, ZN => n12285);
   U1437 : NAND3_X1 port map( A1 => DATA2(26), A2 => DATA1(26), A3 => n12580, 
                           ZN => n12284);
   U1438 : OAI211_X1 port map( C1 => n12286, C2 => n12603, A => n12285, B => 
                           n12284, ZN => n12287);
   U1439 : AOI21_X1 port map( B1 => n12288, B2 => n12293, A => n12287, ZN => 
                           n12291);
   U1440 : NAND3_X1 port map( A1 => n12551, A2 => n12442, A3 => n12289, ZN => 
                           n12290);
   U1441 : OAI211_X1 port map( C1 => n12293, C2 => n12292, A => n12291, B => 
                           n12290, ZN => OUTALU(26));
   U1442 : NAND2_X1 port map( A1 => n12740, A2 => DATA2_I_24_port, ZN => n12312
                           );
   U1443 : NAND2_X1 port map( A1 => n12313, A2 => n12294, ZN => n12309);
   U1444 : NOR3_X1 port map( A1 => n12415, A2 => n12360, A3 => n12603, ZN => 
                           n12302);
   U1445 : INV_X1 port map( A => DATA2(25), ZN => n12934);
   U1446 : NOR2_X1 port map( A1 => n12295, A2 => n12934, ZN => n12809);
   U1447 : NAND2_X1 port map( A1 => n12934, A2 => DATA1(25), ZN => n12806);
   U1448 : INV_X1 port map( A => n12806, ZN => n12296);
   U1449 : NOR2_X1 port map( A1 => n12809, A2 => n12296, ZN => n12658);
   U1450 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n12580, 
                           ZN => n12300);
   U1451 : INV_X1 port map( A => n12305, ZN => n12297);
   U1452 : NAND3_X1 port map( A1 => n12298, A2 => n12297, A3 => n12322, ZN => 
                           n12299);
   U1453 : OAI211_X1 port map( C1 => n12658, C2 => n12641, A => n12300, B => 
                           n12299, ZN => n12301);
   U1454 : AOI211_X1 port map( C1 => dataout_mul_25_port, C2 => n12649, A => 
                           n12302, B => n12301, ZN => n12308);
   U1455 : OAI22_X1 port map( A1 => n12439, A2 => n12303, B1 => n12318, B2 => 
                           n12896, ZN => n12306);
   U1456 : AOI22_X1 port map( A1 => n12618, A2 => n12306, B1 => n12305, B2 => 
                           n12304, ZN => n12307);
   U1457 : OAI211_X1 port map( C1 => n12312, C2 => n12309, A => n12308, B => 
                           n12307, ZN => OUTALU(25));
   U1458 : INV_X1 port map( A => DATA2(24), ZN => n12935);
   U1459 : OAI22_X1 port map( A1 => n12935, A2 => n12648, B1 => n12310, B2 => 
                           n12321, ZN => n12317);
   U1460 : OAI22_X1 port map( A1 => n12723, A2 => DATA2(24), B1 => n12935, B2 
                           => n12740, ZN => n12720);
   U1461 : INV_X1 port map( A => n12720, ZN => n12803);
   U1462 : OAI22_X1 port map( A1 => n12415, A2 => n12362, B1 => n12360, B2 => 
                           n12850, ZN => n12311);
   U1463 : AOI22_X1 port map( A1 => n12917, A2 => n12311, B1 => n12649, B2 => 
                           dataout_mul_24_port, ZN => n12315);
   U1464 : NAND3_X1 port map( A1 => n12313, A2 => n12312, A3 => n12322, ZN => 
                           n12314);
   U1465 : OAI211_X1 port map( C1 => n12803, C2 => n12641, A => n12315, B => 
                           n12314, ZN => n12316);
   U1466 : AOI221_X1 port map( B1 => n12521, B2 => DATA1(24), C1 => n12317, C2 
                           => DATA1(24), A => n12316, ZN => n12320);
   U1467 : OR3_X1 port map( A1 => n12610, A2 => n12439, A3 => n12318, ZN => 
                           n12319);
   U1468 : OAI211_X1 port map( C1 => n12322, C2 => n12321, A => n12320, B => 
                           n12319, ZN => OUTALU(24));
   U1469 : NAND2_X1 port map( A1 => n12331, A2 => n12927, ZN => n12498);
   U1470 : INV_X1 port map( A => n12498, ZN => n12519);
   U1471 : INV_X1 port map( A => n12323, ZN => n12324);
   U1472 : NAND2_X1 port map( A1 => n12325, A2 => n12324, ZN => n12483);
   U1473 : AOI22_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, B1 => 
                           n12490, B2 => n12483, ZN => n12453);
   U1474 : AOI21_X1 port map( B1 => n12453, B2 => n12327, A => n12326, ZN => 
                           n12382);
   U1475 : INV_X1 port map( A => n12328, ZN => n12329);
   U1476 : AOI21_X1 port map( B1 => n12395, B2 => n12382, A => n12329, ZN => 
                           n12374);
   U1477 : OAI21_X1 port map( B1 => n12374, B2 => n12380, A => n12330, ZN => 
                           n12342);
   U1478 : NOR2_X1 port map( A1 => n13259, A2 => n12331, ZN => n12517);
   U1479 : AOI22_X1 port map( A1 => n12519, A2 => n12342, B1 => n12517, B2 => 
                           n12343, ZN => n12354);
   U1480 : NAND2_X1 port map( A1 => n12341, A2 => n12346, ZN => n12350);
   U1481 : OAI22_X1 port map( A1 => n12626, A2 => n12332, B1 => n12351, B2 => 
                           n12623, ZN => n12340);
   U1482 : OAI22_X1 port map( A1 => n12384, A2 => n12436, B1 => n12373, B2 => 
                           n12894, ZN => n12339);
   U1483 : NAND2_X1 port map( A1 => n12333, A2 => DATA2(23), ZN => n12802);
   U1484 : INV_X1 port map( A => n12802, ZN => n12334);
   U1485 : NOR2_X1 port map( A1 => DATA2(23), A2 => n12333, ZN => n12805);
   U1486 : NOR2_X1 port map( A1 => n12334, A2 => n12805, ZN => n12669);
   U1487 : OAI222_X1 port map( A1 => n12416, A2 => n12362, B1 => n12846, B2 => 
                           n12360, C1 => n12357, C2 => n12415, ZN => n12335);
   U1488 : AOI22_X1 port map( A1 => n12917, A2 => n12335, B1 => n12615, B2 => 
                           dataout_mul_23_port, ZN => n12337);
   U1489 : NAND3_X1 port map( A1 => DATA2(23), A2 => DATA1(23), A3 => n12580, 
                           ZN => n12336);
   U1490 : OAI211_X1 port map( C1 => n12669, C2 => n12641, A => n12337, B => 
                           n12336, ZN => n12338);
   U1491 : AOI221_X1 port map( B1 => n12340, B2 => n12618, C1 => n12339, C2 => 
                           n12551, A => n12338, ZN => n12349);
   U1492 : INV_X1 port map( A => n12341, ZN => n12353);
   U1493 : INV_X1 port map( A => n12517, ZN => n12497);
   U1494 : OAI22_X1 port map( A1 => n12343, A2 => n12497, B1 => n12498, B2 => 
                           n12342, ZN => n12344);
   U1495 : NOR2_X1 port map( A1 => n12353, A2 => n12344, ZN => n12352);
   U1496 : OAI21_X1 port map( B1 => n12352, B2 => n12346, A => n12347, ZN => 
                           n12345);
   U1497 : OAI211_X1 port map( C1 => n12347, C2 => n12346, A => n12927, B => 
                           n12345, ZN => n12348);
   U1498 : OAI211_X1 port map( C1 => n12354, C2 => n12350, A => n12349, B => 
                           n12348, ZN => OUTALU(23));
   U1499 : INV_X1 port map( A => DATA2(22), ZN => n12937);
   U1500 : OAI22_X1 port map( A1 => n12801, A2 => DATA2(22), B1 => n12937, B2 
                           => DATA1(22), ZN => n12715);
   U1501 : AOI22_X1 port map( A1 => dataout_mul_22_port, A2 => n12615, B1 => 
                           n12622, B2 => n12715, ZN => n12368);
   U1502 : OAI222_X1 port map( A1 => n12894, A2 => n12384, B1 => n12623, B2 => 
                           n12373, C1 => n12351, C2 => n12604, ZN => n12356);
   U1503 : AOI21_X1 port map( B1 => n12354, B2 => n12353, A => n12352, ZN => 
                           n12355);
   U1504 : AOI21_X1 port map( B1 => n12551, B2 => n12356, A => n12355, ZN => 
                           n12367);
   U1505 : OAI22_X1 port map( A1 => n12415, A2 => n12358, B1 => n12357, B2 => 
                           n12416, ZN => n12364);
   U1506 : OAI22_X1 port map( A1 => n12362, A2 => n12361, B1 => n12360, B2 => 
                           n12359, ZN => n12363);
   U1507 : OAI21_X1 port map( B1 => n12364, B2 => n12363, A => n12917, ZN => 
                           n12366);
   U1508 : NAND3_X1 port map( A1 => DATA2(22), A2 => DATA1(22), A3 => n12580, 
                           ZN => n12365);
   U1509 : NAND4_X1 port map( A1 => n12368, A2 => n12367, A3 => n12366, A4 => 
                           n12365, ZN => OUTALU(22));
   U1510 : AOI22_X1 port map( A1 => n12375, A2 => n12517, B1 => n12519, B2 => 
                           n12374, ZN => n12381);
   U1511 : NOR3_X1 port map( A1 => n12474, A2 => n12603, A3 => n12858, ZN => 
                           n12372);
   U1512 : NAND2_X1 port map( A1 => n12369, A2 => DATA2(21), ZN => n12796);
   U1513 : INV_X1 port map( A => n12796, ZN => n12712);
   U1514 : INV_X1 port map( A => DATA2(21), ZN => n12938);
   U1515 : NAND2_X1 port map( A1 => n12938, A2 => DATA1(21), ZN => n12793);
   U1516 : INV_X1 port map( A => n12793, ZN => n12716);
   U1517 : NOR2_X1 port map( A1 => n12712, A2 => n12716, ZN => n12679);
   U1518 : AOI21_X1 port map( B1 => n12520, B2 => DATA2(21), A => n12521, ZN =>
                           n12370);
   U1519 : OAI22_X1 port map( A1 => n12679, A2 => n12641, B1 => n12370, B2 => 
                           n12369, ZN => n12371);
   U1520 : AOI211_X1 port map( C1 => dataout_mul_21_port, C2 => n12649, A => 
                           n12372, B => n12371, ZN => n12379);
   U1521 : OAI22_X1 port map( A1 => n12626, A2 => n12373, B1 => n12384, B2 => 
                           n12623, ZN => n12377);
   U1522 : OAI22_X1 port map( A1 => n12375, A2 => n12497, B1 => n12374, B2 => 
                           n12498, ZN => n12376);
   U1523 : AOI22_X1 port map( A1 => n12551, A2 => n12377, B1 => n12380, B2 => 
                           n12376, ZN => n12378);
   U1524 : OAI211_X1 port map( C1 => n12381, C2 => n12380, A => n12379, B => 
                           n12378, ZN => OUTALU(21));
   U1525 : AOI22_X1 port map( A1 => n12383, A2 => n12517, B1 => n12519, B2 => 
                           n12382, ZN => n12394);
   U1526 : OAI22_X1 port map( A1 => n12383, A2 => n12497, B1 => n12382, B2 => 
                           n12498, ZN => n12392);
   U1527 : NOR3_X1 port map( A1 => n12604, A2 => n12384, A3 => n12610, ZN => 
                           n12391);
   U1528 : AOI21_X1 port map( B1 => n12520, B2 => DATA2(20), A => n12521, ZN =>
                           n12389);
   U1529 : OAI22_X1 port map( A1 => n12475, A2 => n12471, B1 => n12474, B2 => 
                           n12862, ZN => n12385);
   U1530 : AOI22_X1 port map( A1 => n12917, A2 => n12385, B1 => n12649, B2 => 
                           dataout_mul_20_port, ZN => n12387);
   U1531 : NOR2_X1 port map( A1 => DATA2(20), A2 => n12388, ZN => n12799);
   U1532 : INV_X1 port map( A => DATA2(20), ZN => n12939);
   U1533 : NOR2_X1 port map( A1 => n12939, A2 => DATA1(20), ZN => n12660);
   U1534 : OAI21_X1 port map( B1 => n12799, B2 => n12660, A => n12622, ZN => 
                           n12386);
   U1535 : OAI211_X1 port map( C1 => n12389, C2 => n12388, A => n12387, B => 
                           n12386, ZN => n12390);
   U1536 : AOI211_X1 port map( C1 => n12395, C2 => n12392, A => n12391, B => 
                           n12390, ZN => n12393);
   U1537 : OAI21_X1 port map( B1 => n12395, B2 => n12394, A => n12393, ZN => 
                           OUTALU(20));
   U1538 : NOR2_X1 port map( A1 => n12396, A2 => n12640, ZN => n12397);
   U1539 : AOI22_X1 port map( A1 => n12615, A2 => dataout_mul_1_port, B1 => 
                           n12618, B2 => n12397, ZN => n12451);
   U1540 : NOR2_X1 port map( A1 => n12960, A2 => n12398, ZN => n12745);
   U1541 : INV_X1 port map( A => n12745, ZN => n12399);
   U1542 : NAND2_X1 port map( A1 => n12398, A2 => n12960, ZN => n12743);
   U1543 : NAND2_X1 port map( A1 => n12399, A2 => n12743, ZN => n12682);
   U1544 : AOI221_X1 port map( B1 => n12401, B2 => n12400, C1 => n12639, C2 => 
                           n12404, A => n12643, ZN => n12407);
   U1545 : AOI211_X1 port map( C1 => n12405, C2 => n12404, A => n12403, B => 
                           n12402, ZN => n12406);
   U1546 : AOI211_X1 port map( C1 => n12622, C2 => n12682, A => n12407, B => 
                           n12406, ZN => n12450);
   U1547 : AOI21_X1 port map( B1 => n12618, B2 => n12834, A => n12521, ZN => 
                           n12647);
   U1548 : OAI21_X1 port map( B1 => n12960, B2 => n12648, A => n12647, ZN => 
                           n12448);
   U1549 : INV_X1 port map( A => n12904, ZN => n12447);
   U1550 : AOI22_X1 port map( A1 => n12408, A2 => DATA1(2), B1 => n12834, B2 =>
                           DATA1(1), ZN => n12412);
   U1551 : NAND4_X1 port map( A1 => n12412, A2 => n12411, A3 => n12410, A4 => 
                           n12409, ZN => n12841);
   U1552 : AOI222_X1 port map( A1 => n12413, A2 => n12844, B1 => n12841, B2 => 
                           n12842, C1 => n12845, C2 => n12840, ZN => n12851);
   U1553 : OAI22_X1 port map( A1 => n12415, A2 => n12851, B1 => n12414, B2 => 
                           n12846, ZN => n12419);
   U1554 : OAI22_X1 port map( A1 => n12853, A2 => n12417, B1 => n12847, B2 => 
                           n12416, ZN => n12418);
   U1555 : AOI211_X1 port map( C1 => n12857, C2 => n12420, A => n12419, B => 
                           n12418, ZN => n12863);
   U1556 : OAI22_X1 port map( A1 => n12833, A2 => n12860, B1 => n12863, B2 => 
                           n12858, ZN => n12423);
   U1557 : OAI22_X1 port map( A1 => n12865, A2 => n12421, B1 => n12861, B2 => 
                           n12862, ZN => n12422);
   U1558 : AOI211_X1 port map( C1 => n12425, C2 => n12424, A => n12423, B => 
                           n12422, ZN => n12874);
   U1559 : OAI222_X1 port map( A1 => n12875, A2 => n12871, B1 => n12873, B2 => 
                           n12874, C1 => n12426, C2 => n12870, ZN => n12882);
   U1560 : AOI22_X1 port map( A1 => n12879, A2 => n12832, B1 => n12877, B2 => 
                           n12882, ZN => n12429);
   U1561 : AOI22_X1 port map( A1 => n12545, A2 => n12878, B1 => n12880, B2 => 
                           n12427, ZN => n12428);
   U1562 : OAI211_X1 port map( C1 => n12430, C2 => n12886, A => n12429, B => 
                           n12428, ZN => n12830);
   U1563 : AOI22_X1 port map( A1 => n12431, A2 => n12890, B1 => n12889, B2 => 
                           n12830, ZN => n12435);
   U1564 : AOI22_X1 port map( A1 => n12831, A2 => n12433, B1 => n12829, B2 => 
                           n12432, ZN => n12434);
   U1565 : OAI211_X1 port map( C1 => n12437, C2 => n12436, A => n12435, B => 
                           n12434, ZN => n12901);
   U1566 : INV_X1 port map( A => n12901, ZN => n12438);
   U1567 : OAI222_X1 port map( A1 => n12896, A2 => n12441, B1 => n12897, B2 => 
                           n12440, C1 => n12439, C2 => n12438, ZN => n12906);
   U1568 : AOI22_X1 port map( A1 => n12442, A2 => n12906, B1 => n12909, B2 => 
                           n12910, ZN => n12445);
   U1569 : AOI22_X1 port map( A1 => n12911, A2 => n12443, B1 => n12905, B2 => 
                           n12908, ZN => n12444);
   U1570 : OAI211_X1 port map( C1 => n12447, C2 => n12446, A => n12445, B => 
                           n12444, ZN => n12920);
   U1571 : AOI22_X1 port map( A1 => DATA1(1), A2 => n12448, B1 => n12917, B2 =>
                           n12920, ZN => n12449);
   U1572 : NAND3_X1 port map( A1 => n12451, A2 => n12450, A3 => n12449, ZN => 
                           OUTALU(1));
   U1573 : AOI22_X1 port map( A1 => n12454, A2 => n12517, B1 => n12519, B2 => 
                           n12453, ZN => n12468);
   U1574 : INV_X1 port map( A => n12452, ZN => n12467);
   U1575 : OAI22_X1 port map( A1 => n12454, A2 => n12497, B1 => n12453, B2 => 
                           n12498, ZN => n12465);
   U1576 : OAI222_X1 port map( A1 => n12860, A2 => n12474, B1 => n12858, B2 => 
                           n12470, C1 => n12862, C2 => n12475, ZN => n12455);
   U1577 : AOI22_X1 port map( A1 => n12917, A2 => n12455, B1 => n12649, B2 => 
                           dataout_mul_19_port, ZN => n12463);
   U1578 : OAI22_X1 port map( A1 => n12514, A2 => n12456, B1 => n12481, B2 => 
                           n12495, ZN => n12458);
   U1579 : OAI22_X1 port map( A1 => n12496, A2 => n12482, B1 => n12513, B2 => 
                           n12886, ZN => n12457);
   U1580 : OAI21_X1 port map( B1 => n12458, B2 => n12457, A => n12551, ZN => 
                           n12462);
   U1581 : NAND3_X1 port map( A1 => DATA2(19), A2 => DATA1(19), A3 => n12580, 
                           ZN => n12461);
   U1582 : NOR2_X1 port map( A1 => DATA2(19), A2 => n12459, ZN => n12789);
   U1583 : INV_X1 port map( A => DATA2(19), ZN => n12940);
   U1584 : NOR2_X1 port map( A1 => n12940, A2 => DATA1(19), ZN => n12659);
   U1585 : OAI21_X1 port map( B1 => n12789, B2 => n12659, A => n12622, ZN => 
                           n12460);
   U1586 : NAND4_X1 port map( A1 => n12463, A2 => n12462, A3 => n12461, A4 => 
                           n12460, ZN => n12464);
   U1587 : AOI21_X1 port map( B1 => n12465, B2 => n12467, A => n12464, ZN => 
                           n12466);
   U1588 : OAI21_X1 port map( B1 => n12468, B2 => n12467, A => n12466, ZN => 
                           OUTALU(19));
   U1589 : AOI22_X1 port map( A1 => n12519, A2 => n12483, B1 => n12517, B2 => 
                           n12484, ZN => n12489);
   U1590 : INV_X1 port map( A => DATA2(18), ZN => n12941);
   U1591 : NOR3_X1 port map( A1 => n12616, A2 => n12941, A3 => n12469, ZN => 
                           n12480);
   U1592 : NAND2_X1 port map( A1 => n12941, A2 => DATA1(18), ZN => n12788);
   U1593 : NAND2_X1 port map( A1 => DATA2(18), A2 => n12469, ZN => n12792);
   U1594 : OAI22_X1 port map( A1 => n12472, A2 => n12471, B1 => n12470, B2 => 
                           n12862, ZN => n12477);
   U1595 : OAI22_X1 port map( A1 => n12475, A2 => n12860, B1 => n12474, B2 => 
                           n12473, ZN => n12476);
   U1596 : OAI21_X1 port map( B1 => n12477, B2 => n12476, A => n12917, ZN => 
                           n12478);
   U1597 : OAI221_X1 port map( B1 => n12641, B2 => n12788, C1 => n12641, C2 => 
                           n12792, A => n12478, ZN => n12479);
   U1598 : AOI211_X1 port map( C1 => n12649, C2 => dataout_mul_18_port, A => 
                           n12480, B => n12479, ZN => n12488);
   U1599 : OAI222_X1 port map( A1 => n12482, A2 => n12513, B1 => n12495, B2 => 
                           n12496, C1 => n12481, C2 => n12514, ZN => n12486);
   U1600 : OAI22_X1 port map( A1 => n12484, A2 => n12497, B1 => n12498, B2 => 
                           n12483, ZN => n12485);
   U1601 : AOI22_X1 port map( A1 => n12618, A2 => n12486, B1 => n12490, B2 => 
                           n12485, ZN => n12487);
   U1602 : OAI211_X1 port map( C1 => n12490, C2 => n12489, A => n12488, B => 
                           n12487, ZN => OUTALU(18));
   U1603 : AOI22_X1 port map( A1 => n12519, A2 => n12511, B1 => n12517, B2 => 
                           n12510, ZN => n12504);
   U1604 : NOR3_X1 port map( A1 => n12505, A2 => n12603, A3 => n12506, ZN => 
                           n12494);
   U1605 : NAND2_X1 port map( A1 => n12491, A2 => DATA2(17), ZN => n12741);
   U1606 : INV_X1 port map( A => DATA2(17), ZN => n12942);
   U1607 : NAND2_X1 port map( A1 => n12942, A2 => DATA1(17), ZN => n12785);
   U1608 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n12580, 
                           ZN => n12492);
   U1609 : OAI221_X1 port map( B1 => n12641, B2 => n12741, C1 => n12641, C2 => 
                           n12785, A => n12492, ZN => n12493);
   U1610 : AOI211_X1 port map( C1 => dataout_mul_17_port, C2 => n12649, A => 
                           n12494, B => n12493, ZN => n12502);
   U1611 : OAI22_X1 port map( A1 => n12514, A2 => n12496, B1 => n12513, B2 => 
                           n12495, ZN => n12500);
   U1612 : OAI22_X1 port map( A1 => n12511, A2 => n12498, B1 => n12510, B2 => 
                           n12497, ZN => n12499);
   U1613 : AOI22_X1 port map( A1 => n12618, A2 => n12500, B1 => n12503, B2 => 
                           n12499, ZN => n12501);
   U1614 : OAI211_X1 port map( C1 => n12504, C2 => n12503, A => n12502, B => 
                           n12501, ZN => OUTALU(17));
   U1615 : OAI22_X1 port map( A1 => n12507, A2 => n12506, B1 => n12505, B2 => 
                           n12875, ZN => n12509);
   U1616 : AOI22_X1 port map( A1 => n12917, A2 => n12509, B1 => n12508, B2 => 
                           dataout_mul_16_port, ZN => n12525);
   U1617 : INV_X1 port map( A => n12510, ZN => n12512);
   U1618 : NOR2_X1 port map( A1 => n12512, A2 => n12511, ZN => n12516);
   U1619 : INV_X1 port map( A => n12516, ZN => n12518);
   U1620 : NOR3_X1 port map( A1 => n12514, A2 => n12513, A3 => n12610, ZN => 
                           n12515);
   U1621 : AOI221_X1 port map( B1 => n12519, B2 => n12518, C1 => n12517, C2 => 
                           n12516, A => n12515, ZN => n12524);
   U1622 : INV_X1 port map( A => DATA2(16), ZN => n12943);
   U1623 : AND2_X1 port map( A1 => n12943, A2 => DATA1(16), ZN => n12784);
   U1624 : NOR2_X1 port map( A1 => DATA1(16), A2 => n12943, ZN => n12665);
   U1625 : OAI21_X1 port map( B1 => n12784, B2 => n12665, A => n12622, ZN => 
                           n12523);
   U1626 : OAI211_X1 port map( C1 => n12521, C2 => n12520, A => DATA2(16), B =>
                           DATA1(16), ZN => n12522);
   U1627 : NAND4_X1 port map( A1 => n12525, A2 => n12524, A3 => n12523, A4 => 
                           n12522, ZN => OUTALU(16));
   U1628 : AOI22_X1 port map( A1 => n12550, A2 => n12527, B1 => n12526, B2 => 
                           n12549, ZN => n12544);
   U1629 : INV_X1 port map( A => n12535, ZN => n12530);
   U1630 : INV_X1 port map( A => n12528, ZN => n12529);
   U1631 : AOI221_X1 port map( B1 => n12530, B2 => n12529, C1 => n12535, C2 => 
                           n12528, A => n12612, ZN => n12540);
   U1632 : NAND2_X1 port map( A1 => n12531, A2 => DATA2(15), ZN => n12783);
   U1633 : INV_X1 port map( A => DATA2(15), ZN => n12944);
   U1634 : OAI221_X1 port map( B1 => DATA2(15), B2 => n12622, C1 => n12944, C2 
                           => n12580, A => DATA1(15), ZN => n12538);
   U1635 : NAND2_X1 port map( A1 => n12532, A2 => n12556, ZN => n12554);
   U1636 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n12559, B2 => n12554, ZN => n12536);
   U1637 : AOI21_X1 port map( B1 => n12536, B2 => n12535, A => n12533, ZN => 
                           n12534);
   U1638 : OAI21_X1 port map( B1 => n12536, B2 => n12535, A => n12534, ZN => 
                           n12537);
   U1639 : OAI211_X1 port map( C1 => n12641, C2 => n12783, A => n12538, B => 
                           n12537, ZN => n12539);
   U1640 : AOI211_X1 port map( C1 => n12649, C2 => dataout_mul_15_port, A => 
                           n12540, B => n12539, ZN => n12543);
   U1641 : NAND3_X1 port map( A1 => n12917, A2 => n12541, A3 => n12572, ZN => 
                           n12542);
   U1642 : OAI211_X1 port map( C1 => n12544, C2 => n12610, A => n12543, B => 
                           n12542, ZN => OUTALU(15));
   U1643 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           ZN => n13191);
   U1644 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A => n13191, ZN => n13192);
   U1645 : NOR3_X1 port map( A1 => n5126, A2 => n5134, A3 => n13192, ZN => 
                           n3087);
   U1646 : AOI22_X1 port map( A1 => n12545, A2 => n12572, B1 => n12877, B2 => 
                           n12571, ZN => n12567);
   U1647 : OR2_X1 port map( A1 => n5134, A2 => n13192, ZN => n12547);
   U1648 : AOI211_X1 port map( C1 => n5126, C2 => n12547, A => n3087, B => 
                           n12546, ZN => n12565);
   U1649 : INV_X1 port map( A => DATA2(14), ZN => n12945);
   U1650 : NOR3_X1 port map( A1 => n12616, A2 => n12945, A3 => n12548, ZN => 
                           n12564);
   U1651 : NAND2_X1 port map( A1 => n12548, A2 => DATA2(14), ZN => n12775);
   U1652 : NOR2_X1 port map( A1 => n12548, A2 => DATA2(14), ZN => n12703);
   U1653 : INV_X1 port map( A => n12703, ZN => n12779);
   U1654 : NAND3_X1 port map( A1 => n12551, A2 => n12550, A3 => n12549, ZN => 
                           n12552);
   U1655 : OAI221_X1 port map( B1 => n12641, B2 => n12775, C1 => n12641, C2 => 
                           n12779, A => n12552, ZN => n12563);
   U1656 : AOI22_X1 port map( A1 => n12627, A2 => n12554, B1 => n12585, B2 => 
                           n12553, ZN => n12555);
   U1657 : INV_X1 port map( A => n12555, ZN => n12561);
   U1658 : INV_X1 port map( A => n12556, ZN => n12558);
   U1659 : NOR2_X1 port map( A1 => n12558, A2 => n12557, ZN => n12560);
   U1660 : MUX2_X1 port map( A => n12561, B => n12560, S => n12559, Z => n12562
                           );
   U1661 : NOR4_X1 port map( A1 => n12565, A2 => n12564, A3 => n12563, A4 => 
                           n12562, ZN => n12566);
   U1662 : OAI21_X1 port map( B1 => n12567, B2 => n12603, A => n12566, ZN => 
                           OUTALU(14));
   U1663 : AOI222_X1 port map( A1 => n12593, A2 => n12570, B1 => n12619, B2 => 
                           n12569, C1 => n12568, C2 => n12617, ZN => n12592);
   U1664 : AOI22_X1 port map( A1 => n12573, A2 => n12572, B1 => n12879, B2 => 
                           n12571, ZN => n12577);
   U1665 : AOI22_X1 port map( A1 => n12883, A2 => n12575, B1 => n12877, B2 => 
                           n12574, ZN => n12576);
   U1666 : AOI21_X1 port map( B1 => n12577, B2 => n12576, A => n12603, ZN => 
                           n12584);
   U1667 : AOI22_X1 port map( A1 => DATA1(12), A2 => n12947, B1 => DATA2(12), 
                           B2 => n12772, ZN => n12768);
   U1668 : OAI211_X1 port map( C1 => n12586, C2 => n12579, A => n12627, B => 
                           n12578, ZN => n12582);
   U1669 : NAND3_X1 port map( A1 => DATA2(12), A2 => DATA1(12), A3 => n12580, 
                           ZN => n12581);
   U1670 : OAI211_X1 port map( C1 => n12768, C2 => n12641, A => n12582, B => 
                           n12581, ZN => n12583);
   U1671 : AOI211_X1 port map( C1 => n12649, C2 => dataout_mul_12_port, A => 
                           n12584, B => n12583, ZN => n12591);
   U1672 : INV_X1 port map( A => n12587, ZN => n12589);
   U1673 : OAI221_X1 port map( B1 => n12589, B2 => n12588, C1 => n12587, C2 => 
                           n12586, A => n12585, ZN => n12590);
   U1674 : OAI211_X1 port map( C1 => n12592, C2 => n12610, A => n12591, B => 
                           n12590, ZN => OUTALU(12));
   U1675 : AOI22_X1 port map( A1 => n12594, A2 => n12619, B1 => n12617, B2 => 
                           n12593, ZN => n12611);
   U1676 : NAND2_X1 port map( A1 => n12595, A2 => DATA2(11), ZN => n12767);
   U1677 : NAND2_X1 port map( A1 => DATA1(11), A2 => n12948, ZN => n12700);
   U1678 : AOI21_X1 port map( B1 => n12767, B2 => n12700, A => n12641, ZN => 
                           n12597);
   U1679 : NOR3_X1 port map( A1 => n12616, A2 => n12948, A3 => n12595, ZN => 
                           n12596);
   U1680 : AOI211_X1 port map( C1 => dataout_mul_11_port, C2 => n12615, A => 
                           n12597, B => n12596, ZN => n12609);
   U1681 : INV_X1 port map( A => n12601, ZN => n12599);
   U1682 : XNOR2_X1 port map( A => n12598, B => n12599, ZN => n12607);
   U1683 : INV_X1 port map( A => n12602, ZN => n12600);
   U1684 : AOI221_X1 port map( B1 => n12602, B2 => n12601, C1 => n12600, C2 => 
                           n12599, A => n12612, ZN => n12606);
   U1685 : NOR3_X1 port map( A1 => n12604, A2 => n12624, A3 => n12603, ZN => 
                           n12605);
   U1686 : AOI211_X1 port map( C1 => n12607, C2 => n12627, A => n12606, B => 
                           n12605, ZN => n12608);
   U1687 : OAI211_X1 port map( C1 => n12611, C2 => n12610, A => n12609, B => 
                           n12608, ZN => OUTALU(11));
   U1688 : NOR2_X1 port map( A1 => n12613, A2 => n12612, ZN => n12631);
   U1689 : AOI22_X1 port map( A1 => n12615, A2 => dataout_mul_10_port, B1 => 
                           n12614, B2 => n12631, ZN => n12638);
   U1690 : AOI22_X1 port map( A1 => DATA1(10), A2 => DATA2(10), B1 => n12949, 
                           B2 => n12651, ZN => n12764);
   U1691 : NOR3_X1 port map( A1 => n12616, A2 => n12949, A3 => n12651, ZN => 
                           n12621);
   U1692 : AND3_X1 port map( A1 => n12619, A2 => n12618, A3 => n12617, ZN => 
                           n12620);
   U1693 : AOI211_X1 port map( C1 => n12622, C2 => n12764, A => n12621, B => 
                           n12620, ZN => n12637);
   U1694 : OAI22_X1 port map( A1 => n12626, A2 => n12625, B1 => n12624, B2 => 
                           n12623, ZN => n12630);
   U1695 : AND2_X1 port map( A1 => n12628, A2 => n12627, ZN => n12632);
   U1696 : AOI22_X1 port map( A1 => n12917, A2 => n12630, B1 => n12629, B2 => 
                           n12632, ZN => n12636);
   U1697 : OAI22_X1 port map( A1 => n12634, A2 => n12633, B1 => n12632, B2 => 
                           n12631, ZN => n12635);
   U1698 : NAND4_X1 port map( A1 => n12638, A2 => n12637, A3 => n12636, A4 => 
                           n12635, ZN => OUTALU(10));
   U1699 : OAI21_X1 port map( B1 => DATA1(0), B2 => DATA2_I_0_port, A => n12639
                           , ZN => n12645);
   U1700 : OAI22_X1 port map( A1 => n12961, A2 => n12640, B1 => DATA1(0), B2 =>
                           DATA2(0), ZN => n12661);
   U1701 : OR2_X1 port map( A1 => n12641, A2 => n12661, ZN => n12642);
   U1702 : OAI21_X1 port map( B1 => n12643, B2 => n12645, A => n12642, ZN => 
                           n12644);
   U1703 : AOI21_X1 port map( B1 => n12646, B2 => n12645, A => n12644, ZN => 
                           n12925);
   U1704 : OAI21_X1 port map( B1 => n12961, B2 => n12648, A => n12647, ZN => 
                           n12650);
   U1705 : AOI22_X1 port map( A1 => DATA1(0), A2 => n12650, B1 => n12649, B2 =>
                           dataout_mul_0_port, ZN => n12924);
   U1706 : OAI21_X1 port map( B1 => DATA2(10), B2 => n12651, A => n12700, ZN =>
                           n12769);
   U1707 : AOI22_X1 port map( A1 => DATA2(5), A2 => n12652, B1 => DATA2(6), B2 
                           => n12691, ZN => n12752);
   U1708 : NOR4_X1 port map( A1 => n12656, A2 => n12655, A3 => n12654, A4 => 
                           n12653, ZN => n12657);
   U1709 : NAND3_X1 port map( A1 => n12752, A2 => n12658, A3 => n12657, ZN => 
                           n12681);
   U1710 : INV_X1 port map( A => n12659, ZN => n12709);
   U1711 : INV_X1 port map( A => n12660, ZN => n12717);
   U1712 : NAND2_X1 port map( A1 => n12709, A2 => n12717, ZN => n12794);
   U1713 : NAND4_X1 port map( A1 => FUNC(2), A2 => n12692, A3 => n12779, A4 => 
                           n12815, ZN => n12663);
   U1714 : INV_X1 port map( A => n12727, ZN => n12814);
   U1715 : NAND4_X1 port map( A1 => n12661, A2 => n12792, A3 => n12688, A4 => 
                           n12814, ZN => n12662);
   U1716 : NOR4_X1 port map( A1 => n12794, A2 => n12664, A3 => n12663, A4 => 
                           n12662, ZN => n12677);
   U1717 : NAND2_X1 port map( A1 => n12775, A2 => n12783, ZN => n12707);
   U1718 : AOI21_X1 port map( B1 => DATA1(15), B2 => n12944, A => n12784, ZN =>
                           n12780);
   U1719 : INV_X1 port map( A => n12780, ZN => n12666);
   U1720 : INV_X1 port map( A => n12665, ZN => n12782);
   U1721 : NAND2_X1 port map( A1 => n12782, A2 => n12741, ZN => n12706);
   U1722 : NAND2_X1 port map( A1 => n12785, A2 => n12788, ZN => n12710);
   U1723 : OR4_X1 port map( A1 => n12707, A2 => n12666, A3 => n12706, A4 => 
                           n12710, ZN => n12675);
   U1724 : NAND2_X1 port map( A1 => n12690, A2 => n12685, ZN => n12753);
   U1725 : INV_X1 port map( A => n12768, ZN => n12667);
   U1726 : OAI21_X1 port map( B1 => n12949, B2 => DATA1(10), A => n12767, ZN =>
                           n12701);
   U1727 : OR4_X1 port map( A1 => n12753, A2 => n12742, A3 => n12667, A4 => 
                           n12701, ZN => n12674);
   U1728 : INV_X1 port map( A => n12668, ZN => n12811);
   U1729 : NOR2_X1 port map( A1 => n12811, A2 => n12822, ZN => n12729);
   U1730 : NAND4_X1 port map( A1 => n12670, A2 => n12729, A3 => n12820, A4 => 
                           n12669, ZN => n12673);
   U1731 : NOR2_X1 port map( A1 => n12799, A2 => n12789, ZN => n12714);
   U1732 : INV_X1 port map( A => n12715, ZN => n12797);
   U1733 : INV_X1 port map( A => n12671, ZN => n12756);
   U1734 : NAND4_X1 port map( A1 => n12714, A2 => n12797, A3 => n12803, A4 => 
                           n12756, ZN => n12672);
   U1735 : NOR4_X1 port map( A1 => n12675, A2 => n12674, A3 => n12673, A4 => 
                           n12672, ZN => n12676);
   U1736 : NAND4_X1 port map( A1 => n12679, A2 => n12678, A3 => n12677, A4 => 
                           n12676, ZN => n12680);
   U1737 : NOR4_X1 port map( A1 => n12769, A2 => n12682, A3 => n12681, A4 => 
                           n12680, ZN => n12739);
   U1738 : AOI21_X1 port map( B1 => DATA2(12), B2 => n12772, A => n12773, ZN =>
                           n12705);
   U1739 : NOR2_X1 port map( A1 => DATA1(0), A2 => n12961, ZN => n12683);
   U1740 : AOI21_X1 port map( B1 => n12683, B2 => n12743, A => n12745, ZN => 
                           n12684);
   U1741 : OAI22_X1 port map( A1 => DATA1(2), A2 => n12959, B1 => n12684, B2 =>
                           n12742, ZN => n12686);
   U1742 : OAI211_X1 port map( C1 => n12749, C2 => n12686, A => n12685, B => 
                           n12750, ZN => n12687);
   U1743 : OAI211_X1 port map( C1 => n13261, C2 => n12956, A => n12688, B => 
                           n12687, ZN => n12689);
   U1744 : AOI22_X1 port map( A1 => DATA2(6), A2 => n12691, B1 => n12690, B2 =>
                           n12689, ZN => n12694);
   U1745 : OAI21_X1 port map( B1 => DATA2(7), B2 => n12693, A => n12692, ZN => 
                           n12759);
   U1746 : OAI21_X1 port map( B1 => n12694, B2 => n12759, A => n12757, ZN => 
                           n12695);
   U1747 : AOI22_X1 port map( A1 => DATA2(8), A2 => n12696, B1 => n12762, B2 =>
                           n12695, ZN => n12698);
   U1748 : AOI211_X1 port map( C1 => n12699, C2 => n12698, A => n12697, B => 
                           n12764, ZN => n12702);
   U1749 : OAI211_X1 port map( C1 => n12702, C2 => n12701, A => n12768, B => 
                           n12700, ZN => n12704);
   U1750 : AOI211_X1 port map( C1 => n12705, C2 => n12704, A => n12777, B => 
                           n12703, ZN => n12708);
   U1751 : AOI221_X1 port map( B1 => n12708, B2 => n12780, C1 => n12707, C2 => 
                           n12780, A => n12706, ZN => n12711);
   U1752 : OAI211_X1 port map( C1 => n12711, C2 => n12710, A => n12792, B => 
                           n12709, ZN => n12713);
   U1753 : AOI21_X1 port map( B1 => n12714, B2 => n12713, A => n12712, ZN => 
                           n12718);
   U1754 : AOI211_X1 port map( C1 => n12718, C2 => n12717, A => n12716, B => 
                           n12715, ZN => n12719);
   U1755 : AOI21_X1 port map( B1 => DATA2(22), B2 => n12801, A => n12719, ZN =>
                           n12721);
   U1756 : AOI211_X1 port map( C1 => n12721, C2 => n12802, A => n12805, B => 
                           n12720, ZN => n12722);
   U1757 : AOI211_X1 port map( C1 => DATA2(24), C2 => n12723, A => n12722, B =>
                           n12809, ZN => n12726);
   U1758 : NAND2_X1 port map( A1 => n12806, A2 => n12724, ZN => n12725);
   U1759 : OAI211_X1 port map( C1 => n12726, C2 => n12725, A => n12813, B => 
                           n12815, ZN => n12728);
   U1760 : AOI21_X1 port map( B1 => n12729, B2 => n12728, A => n12727, ZN => 
                           n12732);
   U1761 : AOI211_X1 port map( C1 => n12732, C2 => n12819, A => n12731, B => 
                           n12730, ZN => n12734);
   U1762 : AOI211_X1 port map( C1 => DATA2(30), C2 => n12825, A => n12734, B =>
                           n12733, ZN => n12735);
   U1763 : NOR4_X1 port map( A1 => FUNC(3), A2 => FUNC(2), A3 => n12736, A4 => 
                           n12735, ZN => n12738);
   U1764 : NOR4_X1 port map( A1 => n12739, A2 => FUNC(1), A3 => n12738, A4 => 
                           n12737, ZN => n12919);
   U1765 : NAND2_X1 port map( A1 => n12740, A2 => n12935, ZN => n12808);
   U1766 : INV_X1 port map( A => n12741, ZN => n12787);
   U1767 : INV_X1 port map( A => n12742, ZN => n12747);
   U1768 : NAND2_X1 port map( A1 => DATA1(0), A2 => n12961, ZN => n12744);
   U1769 : OAI21_X1 port map( B1 => n12745, B2 => n12744, A => n12743, ZN => 
                           n12746);
   U1770 : AOI22_X1 port map( A1 => n12747, A2 => n12746, B1 => n13260, B2 => 
                           n12959, ZN => n12751);
   U1771 : AOI211_X1 port map( C1 => n12751, C2 => n12750, A => n12749, B => 
                           n12748, ZN => n12754);
   U1772 : OAI21_X1 port map( B1 => n12754, B2 => n12753, A => n12752, ZN => 
                           n12755);
   U1773 : INV_X1 port map( A => n12755, ZN => n12758);
   U1774 : OAI211_X1 port map( C1 => n12759, C2 => n12758, A => n12757, B => 
                           n12756, ZN => n12761);
   U1775 : AOI21_X1 port map( B1 => n12762, B2 => n12761, A => n12760, ZN => 
                           n12763);
   U1776 : INV_X1 port map( A => n12763, ZN => n12765);
   U1777 : AOI21_X1 port map( B1 => n12766, B2 => n12765, A => n12764, ZN => 
                           n12770);
   U1778 : OAI211_X1 port map( C1 => n12770, C2 => n12769, A => n12768, B => 
                           n12767, ZN => n12771);
   U1779 : OAI21_X1 port map( B1 => DATA2(12), B2 => n12772, A => n12771, ZN =>
                           n12776);
   U1780 : INV_X1 port map( A => n12773, ZN => n12774);
   U1781 : OAI211_X1 port map( C1 => n12777, C2 => n12776, A => n12775, B => 
                           n12774, ZN => n12778);
   U1782 : NAND3_X1 port map( A1 => n12780, A2 => n12779, A3 => n12778, ZN => 
                           n12781);
   U1783 : OAI211_X1 port map( C1 => n12784, C2 => n12783, A => n12782, B => 
                           n12781, ZN => n12786);
   U1784 : OAI21_X1 port map( B1 => n12787, B2 => n12786, A => n12785, ZN => 
                           n12791);
   U1785 : INV_X1 port map( A => n12788, ZN => n12790);
   U1786 : AOI211_X1 port map( C1 => n12792, C2 => n12791, A => n12790, B => 
                           n12789, ZN => n12795);
   U1787 : OAI21_X1 port map( B1 => n12795, B2 => n12794, A => n12793, ZN => 
                           n12798);
   U1788 : OAI211_X1 port map( C1 => n12799, C2 => n12798, A => n12797, B => 
                           n12796, ZN => n12800);
   U1789 : OAI21_X1 port map( B1 => DATA2(22), B2 => n12801, A => n12800, ZN =>
                           n12804);
   U1790 : OAI211_X1 port map( C1 => n12805, C2 => n12804, A => n12803, B => 
                           n12802, ZN => n12807);
   U1791 : OAI221_X1 port map( B1 => n12809, B2 => n12808, C1 => n12809, C2 => 
                           n12807, A => n12806, ZN => n12812);
   U1792 : AOI211_X1 port map( C1 => n12813, C2 => n12812, A => n12811, B => 
                           n12810, ZN => n12818);
   U1793 : NAND2_X1 port map( A1 => n12815, A2 => n12814, ZN => n12817);
   U1794 : OAI21_X1 port map( B1 => n12818, B2 => n12817, A => n12816, ZN => 
                           n12821);
   U1795 : OAI211_X1 port map( C1 => n12822, C2 => n12821, A => n12820, B => 
                           n12819, ZN => n12823);
   U1796 : OAI211_X1 port map( C1 => DATA2(30), C2 => n12825, A => n12824, B =>
                           n12823, ZN => n12826);
   U1797 : OAI221_X1 port map( B1 => FUNC(2), B2 => n12827, C1 => FUNC(2), C2 
                           => n12826, A => FUNC(3), ZN => n12918);
   U1798 : AOI22_X1 port map( A1 => n12831, A2 => n12830, B1 => n12829, B2 => 
                           n12828, ZN => n12893);
   U1799 : INV_X1 port map( A => n12832, ZN => n12887);
   U1800 : INV_X1 port map( A => n12833, ZN => n12868);
   U1801 : AOI22_X1 port map( A1 => n12835, A2 => DATA1(1), B1 => n12834, B2 =>
                           DATA1(0), ZN => n12839);
   U1802 : NAND4_X1 port map( A1 => n12839, A2 => n12838, A3 => n12837, A4 => 
                           n12836, ZN => n12843);
   U1803 : AOI222_X1 port map( A1 => n12845, A2 => n12844, B1 => n12843, B2 => 
                           n12842, C1 => n12841, C2 => n12840, ZN => n12848);
   U1804 : OAI22_X1 port map( A1 => n12849, A2 => n12848, B1 => n12847, B2 => 
                           n12846, ZN => n12855);
   U1805 : OAI22_X1 port map( A1 => n12853, A2 => n12852, B1 => n12851, B2 => 
                           n12850, ZN => n12854);
   U1806 : AOI211_X1 port map( C1 => n12857, C2 => n12856, A => n12855, B => 
                           n12854, ZN => n12859);
   U1807 : OAI22_X1 port map( A1 => n12861, A2 => n12860, B1 => n12859, B2 => 
                           n12858, ZN => n12867);
   U1808 : OAI22_X1 port map( A1 => n12865, A2 => n12864, B1 => n12863, B2 => 
                           n12862, ZN => n12866);
   U1809 : AOI211_X1 port map( C1 => n12869, C2 => n12868, A => n12867, B => 
                           n12866, ZN => n12872);
   U1810 : OAI222_X1 port map( A1 => n12875, A2 => n12874, B1 => n12873, B2 => 
                           n12872, C1 => n12871, C2 => n12870, ZN => n12876);
   U1811 : AOI22_X1 port map( A1 => n12879, A2 => n12878, B1 => n12877, B2 => 
                           n12876, ZN => n12885);
   U1812 : AOI22_X1 port map( A1 => n12883, A2 => n12882, B1 => n12881, B2 => 
                           n12880, ZN => n12884);
   U1813 : OAI211_X1 port map( C1 => n12887, C2 => n12886, A => n12885, B => 
                           n12884, ZN => n12888);
   U1814 : AOI22_X1 port map( A1 => n12891, A2 => n12890, B1 => n12889, B2 => 
                           n12888, ZN => n12892);
   U1815 : OAI211_X1 port map( C1 => n12895, C2 => n12894, A => n12893, B => 
                           n12892, ZN => n12903);
   U1816 : INV_X1 port map( A => n12896, ZN => n12900);
   U1817 : INV_X1 port map( A => n12897, ZN => n12898);
   U1818 : AOI222_X1 port map( A1 => n12903, A2 => n12902, B1 => n12901, B2 => 
                           n12900, C1 => n12899, C2 => n12898, ZN => n12915);
   U1819 : AOI22_X1 port map( A1 => n12907, A2 => n12906, B1 => n12905, B2 => 
                           n12904, ZN => n12913);
   U1820 : AOI22_X1 port map( A1 => n12911, A2 => n12910, B1 => n12909, B2 => 
                           n12908, ZN => n12912);
   U1821 : OAI211_X1 port map( C1 => n12915, C2 => n12914, A => n12913, B => 
                           n12912, ZN => n12916);
   U1822 : AOI22_X1 port map( A1 => n12919, A2 => n12918, B1 => n12917, B2 => 
                           n12916, ZN => n12923);
   U1823 : NAND3_X1 port map( A1 => FUNC(3), A2 => n12921, A3 => n12920, ZN => 
                           n12922);
   U1824 : NAND4_X1 port map( A1 => n12925, A2 => n12924, A3 => n12923, A4 => 
                           n12922, ZN => OUTALU(0));
   U1825 : NAND2_X1 port map( A1 => n12927, A2 => n12926, ZN => n12963);
   U1826 : CLKBUF_X1 port map( A => n12963, Z => n12953);
   U1827 : NAND2_X1 port map( A1 => FUNC(3), A2 => n12927, ZN => n12962);
   U1828 : AOI22_X1 port map( A1 => DATA2(31), A2 => n12953, B1 => n12952, B2 
                           => n12928, ZN => N2548);
   U1829 : AOI22_X1 port map( A1 => DATA2(30), A2 => n12963, B1 => n12962, B2 
                           => n12929, ZN => N2547);
   U1830 : INV_X1 port map( A => DATA2(29), ZN => n12930);
   U1831 : AOI22_X1 port map( A1 => DATA2(29), A2 => n12953, B1 => n12952, B2 
                           => n12930, ZN => N2546);
   U1832 : AOI22_X1 port map( A1 => DATA2(28), A2 => n12963, B1 => n12962, B2 
                           => n12931, ZN => N2545);
   U1833 : AOI22_X1 port map( A1 => DATA2(27), A2 => n12953, B1 => n12952, B2 
                           => n12932, ZN => N2544);
   U1834 : INV_X1 port map( A => DATA2(26), ZN => n12933);
   U1835 : AOI22_X1 port map( A1 => DATA2(26), A2 => n12963, B1 => n12962, B2 
                           => n12933, ZN => N2543);
   U1836 : AOI22_X1 port map( A1 => DATA2(25), A2 => n12953, B1 => n12952, B2 
                           => n12934, ZN => N2542);
   U1837 : AOI22_X1 port map( A1 => DATA2(24), A2 => n12963, B1 => n12962, B2 
                           => n12935, ZN => N2541);
   U1838 : INV_X1 port map( A => DATA2(23), ZN => n12936);
   U1839 : AOI22_X1 port map( A1 => DATA2(23), A2 => n12953, B1 => n12952, B2 
                           => n12936, ZN => N2540);
   U1840 : AOI22_X1 port map( A1 => DATA2(22), A2 => n12963, B1 => n12962, B2 
                           => n12937, ZN => N2539);
   U1841 : AOI22_X1 port map( A1 => DATA2(21), A2 => n12963, B1 => n12962, B2 
                           => n12938, ZN => N2538);
   U1842 : AOI22_X1 port map( A1 => DATA2(20), A2 => n12963, B1 => n12962, B2 
                           => n12939, ZN => N2537);
   U1843 : AOI22_X1 port map( A1 => DATA2(19), A2 => n12953, B1 => n12952, B2 
                           => n12940, ZN => N2536);
   U1844 : AOI22_X1 port map( A1 => DATA2(18), A2 => n12953, B1 => n12952, B2 
                           => n12941, ZN => N2535);
   U1845 : AOI22_X1 port map( A1 => DATA2(17), A2 => n12953, B1 => n12952, B2 
                           => n12942, ZN => N2534);
   U1846 : AOI22_X1 port map( A1 => DATA2(16), A2 => n12953, B1 => n12952, B2 
                           => n12943, ZN => N2533);
   U1847 : AOI22_X1 port map( A1 => DATA2(15), A2 => n12953, B1 => n12952, B2 
                           => n12944, ZN => N2532);
   U1848 : AOI22_X1 port map( A1 => DATA2(14), A2 => n12953, B1 => n12952, B2 
                           => n12945, ZN => N2531);
   U1849 : AOI22_X1 port map( A1 => DATA2(13), A2 => n12953, B1 => n12952, B2 
                           => n12946, ZN => N2530);
   U1850 : AOI22_X1 port map( A1 => DATA2(12), A2 => n12953, B1 => n12952, B2 
                           => n12947, ZN => N2529);
   U1851 : AOI22_X1 port map( A1 => DATA2(11), A2 => n12953, B1 => n12952, B2 
                           => n12948, ZN => N2528);
   U1852 : AOI22_X1 port map( A1 => DATA2(10), A2 => n12953, B1 => n12952, B2 
                           => n12949, ZN => N2527);
   U1853 : AOI22_X1 port map( A1 => DATA2(9), A2 => n12953, B1 => n12952, B2 =>
                           n12950, ZN => N2526);
   U1854 : AOI22_X1 port map( A1 => DATA2(8), A2 => n12953, B1 => n12952, B2 =>
                           n12951, ZN => N2525);
   U1855 : INV_X1 port map( A => DATA2(7), ZN => n12954);
   U1856 : AOI22_X1 port map( A1 => DATA2(7), A2 => n12963, B1 => n12962, B2 =>
                           n12954, ZN => N2524);
   U1857 : AOI22_X1 port map( A1 => DATA2(6), A2 => n12963, B1 => n12962, B2 =>
                           n12955, ZN => N2523);
   U1858 : AOI22_X1 port map( A1 => DATA2(5), A2 => n12963, B1 => n12962, B2 =>
                           n12956, ZN => N2522);
   U1859 : AOI22_X1 port map( A1 => DATA2(4), A2 => n12963, B1 => n12962, B2 =>
                           n12957, ZN => N2521);
   U1860 : AOI22_X1 port map( A1 => DATA2(3), A2 => n12963, B1 => n12962, B2 =>
                           n12958, ZN => N2520);
   U1861 : AOI22_X1 port map( A1 => DATA2(2), A2 => n12963, B1 => n12962, B2 =>
                           n12959, ZN => N2519);
   U1862 : AOI22_X1 port map( A1 => DATA2(1), A2 => n12963, B1 => n12962, B2 =>
                           n12960, ZN => N2518);
   U1863 : AOI22_X1 port map( A1 => DATA2(0), A2 => n12963, B1 => n12962, B2 =>
                           n12961, ZN => N2517);
   U1864 : NOR2_X1 port map( A1 => n12964, A2 => n2008, ZN => 
                           boothmul_pipelined_i_sum_out_1_0_port);
   U1865 : NAND2_X1 port map( A1 => n13005, A2 => data2_mul_3_port, ZN => 
                           n12968);
   U1866 : INV_X1 port map( A => data2_mul_3_port, ZN => n13001);
   U1867 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n13001, ZN => n13000);
   U1868 : INV_X1 port map( A => n12965, ZN => n12966);
   U1869 : NOR2_X1 port map( A1 => n12966, A2 => n13001, ZN => n13003);
   U1870 : NOR2_X1 port map( A1 => data2_mul_3_port, A2 => n12966, ZN => n12993
                           );
   U1871 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n13003, B1 => data1_mul_1_port, B2 => n12993, 
                           ZN => n12967);
   U1872 : OAI221_X1 port map( B1 => n2008, B2 => n12968, C1 => n2008, C2 => 
                           n13000, A => n12967, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1873 : INV_X1 port map( A => n12968, ZN => n13002);
   U1874 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n12993, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n13002, ZN => n12970);
   U1875 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n13003, ZN => n12969);
   U1876 : OAI211_X1 port map( C1 => n2007, C2 => n13000, A => n12970, B => 
                           n12969, ZN => boothmul_pipelined_i_mux_out_1_4_port)
                           ;
   U1877 : CLKBUF_X1 port map( A => n12993, Z => n12997);
   U1878 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n13002, B1 => n12997, B2 => data1_mul_3_port, 
                           ZN => n12972);
   U1879 : CLKBUF_X1 port map( A => n13003, Z => n12994);
   U1880 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n12971);
   U1881 : OAI211_X1 port map( C1 => n13000, C2 => n2005, A => n12972, B => 
                           n12971, ZN => boothmul_pipelined_i_mux_out_1_5_port)
                           ;
   U1882 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B1 => 
                           n12997, B2 => data1_mul_4_port, ZN => n12974);
   U1883 : NAND2_X1 port map( A1 => n13003, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n12973);
   U1884 : OAI211_X1 port map( C1 => n2004, C2 => n13000, A => n12974, B => 
                           n12973, ZN => boothmul_pipelined_i_mux_out_1_6_port)
                           ;
   U1885 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n12997, B2 => data1_mul_5_port, ZN => n12976);
   U1886 : NAND2_X1 port map( A1 => n13003, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n12975);
   U1887 : OAI211_X1 port map( C1 => n2002, C2 => n13000, A => n12976, B => 
                           n12975, ZN => boothmul_pipelined_i_mux_out_1_7_port)
                           ;
   U1888 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n12997, B2 => data1_mul_6_port, ZN => n12978);
   U1889 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n12977);
   U1890 : OAI211_X1 port map( C1 => n2000, C2 => n13000, A => n12978, B => 
                           n12977, ZN => boothmul_pipelined_i_mux_out_1_8_port)
                           ;
   U1891 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n12993, B2 => data1_mul_7_port, ZN => n12980);
   U1892 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n12979);
   U1893 : OAI211_X1 port map( C1 => n1998, C2 => n13000, A => n12980, B => 
                           n12979, ZN => boothmul_pipelined_i_mux_out_1_9_port)
                           ;
   U1894 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n12993, B2 => data1_mul_8_port, ZN => n12982);
   U1895 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n12981);
   U1896 : OAI211_X1 port map( C1 => n1993, C2 => n13000, A => n12982, B => 
                           n12981, ZN => boothmul_pipelined_i_mux_out_1_10_port
                           );
   U1897 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n12997, B2 => data1_mul_9_port, ZN => n12984);
   U1898 : NAND2_X1 port map( A1 => n13003, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n12983);
   U1899 : OAI211_X1 port map( C1 => n1990, C2 => n13000, A => n12984, B => 
                           n12983, ZN => boothmul_pipelined_i_mux_out_1_11_port
                           );
   U1900 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n12993, B2 => data1_mul_10_port, ZN => n12986);
   U1901 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n12985);
   U1902 : OAI211_X1 port map( C1 => n1988, C2 => n13000, A => n12986, B => 
                           n12985, ZN => boothmul_pipelined_i_mux_out_1_12_port
                           );
   U1903 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n12997, B2 => data1_mul_11_port, ZN => n12988);
   U1904 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n12987);
   U1905 : OAI211_X1 port map( C1 => n1986, C2 => n13000, A => n12988, B => 
                           n12987, ZN => boothmul_pipelined_i_mux_out_1_13_port
                           );
   U1906 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n12997, B2 => data1_mul_12_port, ZN => n12990);
   U1907 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n12989);
   U1908 : OAI211_X1 port map( C1 => n1984, C2 => n13000, A => n12990, B => 
                           n12989, ZN => boothmul_pipelined_i_mux_out_1_14_port
                           );
   U1909 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n12993, B2 => data1_mul_13_port, ZN => n12992);
   U1910 : NAND2_X1 port map( A1 => n13003, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n12991);
   U1911 : OAI211_X1 port map( C1 => n1982, C2 => n13000, A => n12992, B => 
                           n12991, ZN => boothmul_pipelined_i_mux_out_1_15_port
                           );
   U1912 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n12993, B2 => data1_mul_14_port, ZN => n12996);
   U1913 : NAND2_X1 port map( A1 => n12994, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n12995);
   U1914 : OAI211_X1 port map( C1 => n1980, C2 => n13000, A => n12996, B => 
                           n12995, ZN => boothmul_pipelined_i_mux_out_1_16_port
                           );
   U1915 : AOI22_X1 port map( A1 => n13002, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n12997, B2 => data1_mul_15_port, ZN => n12999);
   U1916 : NAND2_X1 port map( A1 => n13003, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n12998);
   U1917 : OAI211_X1 port map( C1 => n1978, C2 => n13000, A => n12999, B => 
                           n12998, ZN => boothmul_pipelined_i_mux_out_1_17_port
                           );
   U1918 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n13001, ZN => 
                           n13006);
   U1919 : AOI22_X1 port map( A1 => n13003, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n13002, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n13004);
   U1920 : OAI21_X1 port map( B1 => n13006, B2 => n13005, A => n13004, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1921 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n13045);
   U1922 : NAND2_X1 port map( A1 => n13045, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n13009);
   U1923 : NAND3_X1 port map( A1 => n3076, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n13041);
   U1924 : NOR2_X1 port map( A1 => n3076, A2 => n13007, ZN => n13022);
   U1925 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n13007, ZN => n13035);
   U1926 : CLKBUF_X1 port map( A => n13035, Z => n13038);
   U1927 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n13022, B1 => data1_mul_1_port, B2 => n13038, 
                           ZN => n13008);
   U1928 : OAI221_X1 port map( B1 => n2008, B2 => n13009, C1 => n2008, C2 => 
                           n13041, A => n13008, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1929 : INV_X1 port map( A => n13009, ZN => n13043);
   U1930 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n13035, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n13043, ZN => n13011);
   U1931 : CLKBUF_X1 port map( A => n13022, Z => n13042);
   U1932 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n13042, ZN => n13010);
   U1933 : OAI211_X1 port map( C1 => n13041, C2 => n2007, A => n13011, B => 
                           n13010, ZN => boothmul_pipelined_i_mux_out_2_6_port)
                           ;
   U1934 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n13043, B1 => data1_mul_3_port, B2 => n13038, 
                           ZN => n13013);
   U1935 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n13022, ZN => n13012);
   U1936 : OAI211_X1 port map( C1 => n13041, C2 => n2005, A => n13013, B => 
                           n13012, ZN => boothmul_pipelined_i_mux_out_2_7_port)
                           ;
   U1937 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n13043, B1 => data1_mul_4_port, B2 => n13038, 
                           ZN => n13015);
   U1938 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n13022, ZN => n13014);
   U1939 : OAI211_X1 port map( C1 => n13041, C2 => n2004, A => n13015, B => 
                           n13014, ZN => boothmul_pipelined_i_mux_out_2_8_port)
                           ;
   U1940 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n13043, B1 => data1_mul_5_port, B2 => n13035, 
                           ZN => n13017);
   U1941 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n13022, ZN => n13016);
   U1942 : OAI211_X1 port map( C1 => n13041, C2 => n2002, A => n13017, B => 
                           n13016, ZN => boothmul_pipelined_i_mux_out_2_9_port)
                           ;
   U1943 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n13043, B1 => data1_mul_6_port, B2 => n13038, 
                           ZN => n13019);
   U1944 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n13022, ZN => n13018);
   U1945 : OAI211_X1 port map( C1 => n13041, C2 => n2000, A => n13019, B => 
                           n13018, ZN => boothmul_pipelined_i_mux_out_2_10_port
                           );
   U1946 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n13043, B1 => data1_mul_7_port, B2 => n13035, 
                           ZN => n13021);
   U1947 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n13022, ZN => n13020);
   U1948 : OAI211_X1 port map( C1 => n13041, C2 => n1998, A => n13021, B => 
                           n13020, ZN => boothmul_pipelined_i_mux_out_2_11_port
                           );
   U1949 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n13043, B1 => data1_mul_8_port, B2 => n13038, 
                           ZN => n13024);
   U1950 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n13022, ZN => n13023);
   U1951 : OAI211_X1 port map( C1 => n13041, C2 => n1993, A => n13024, B => 
                           n13023, ZN => boothmul_pipelined_i_mux_out_2_12_port
                           );
   U1952 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n13043, B1 => data1_mul_9_port, B2 => n13038, 
                           ZN => n13026);
   U1953 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n13042, ZN => n13025);
   U1954 : OAI211_X1 port map( C1 => n13041, C2 => n1990, A => n13026, B => 
                           n13025, ZN => boothmul_pipelined_i_mux_out_2_13_port
                           );
   U1955 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n13043, B1 => data1_mul_10_port, B2 => n13035,
                           ZN => n13028);
   U1956 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n13042, ZN => n13027);
   U1957 : OAI211_X1 port map( C1 => n13041, C2 => n1988, A => n13028, B => 
                           n13027, ZN => boothmul_pipelined_i_mux_out_2_14_port
                           );
   U1958 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n13043, B1 => data1_mul_11_port, B2 => n13035,
                           ZN => n13030);
   U1959 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n13042, ZN => n13029);
   U1960 : OAI211_X1 port map( C1 => n13041, C2 => n1986, A => n13030, B => 
                           n13029, ZN => boothmul_pipelined_i_mux_out_2_15_port
                           );
   U1961 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n13043, B1 => data1_mul_12_port, B2 => n13038,
                           ZN => n13032);
   U1962 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n13042, ZN => n13031);
   U1963 : OAI211_X1 port map( C1 => n13041, C2 => n1984, A => n13032, B => 
                           n13031, ZN => boothmul_pipelined_i_mux_out_2_16_port
                           );
   U1964 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n13043, B1 => data1_mul_13_port, B2 => n13035,
                           ZN => n13034);
   U1965 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n13042, ZN => n13033);
   U1966 : OAI211_X1 port map( C1 => n13041, C2 => n1982, A => n13034, B => 
                           n13033, ZN => boothmul_pipelined_i_mux_out_2_17_port
                           );
   U1967 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n13043, B1 => data1_mul_14_port, B2 => n13035,
                           ZN => n13037);
   U1968 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n13042, ZN => n13036);
   U1969 : OAI211_X1 port map( C1 => n13041, C2 => n1980, A => n13037, B => 
                           n13036, ZN => boothmul_pipelined_i_mux_out_2_18_port
                           );
   U1970 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n13043, B1 => data1_mul_15_port, B2 => n13038,
                           ZN => n13040);
   U1971 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n13042, ZN => n13039);
   U1972 : OAI211_X1 port map( C1 => n13041, C2 => n1978, A => n13040, B => 
                           n13039, ZN => boothmul_pipelined_i_mux_out_2_19_port
                           );
   U1973 : NAND2_X1 port map( A1 => n3076, A2 => data1_mul_15_port, ZN => 
                           n13046);
   U1974 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n13043, B1 => n13042, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n13044);
   U1975 : OAI21_X1 port map( B1 => n13046, B2 => n13045, A => n13044, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U1976 : NAND3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n13256);
   U1977 : NOR3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_6_port, 
                           ZN => n13254);
   U1978 : INV_X1 port map( A => n13254, ZN => n13050);
   U1979 : INV_X1 port map( A => n13048, ZN => n13047);
   U1980 : NAND2_X1 port map( A1 => n3082, A2 => n13047, ZN => n13257);
   U1981 : INV_X1 port map( A => n13257, ZN => n13076);
   U1982 : NOR2_X1 port map( A1 => n3082, A2 => n13048, ZN => n13080);
   U1983 : CLKBUF_X1 port map( A => n13080, Z => n13253);
   U1984 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_60_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n13049);
   U1985 : OAI221_X1 port map( B1 => n3077, B2 => n13256, C1 => n3077, C2 => 
                           n13050, A => n13049, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1986 : INV_X1 port map( A => n13256, ZN => n13079);
   U1987 : CLKBUF_X1 port map( A => n13254, Z => n13075);
   U1988 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_3_60_port, A2
                           => n13079, B1 => n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n13052);
   U1989 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => 
                           n13080, B2 => 
                           boothmul_pipelined_i_muxes_in_3_175_port, ZN => 
                           n13051);
   U1990 : NAND2_X1 port map( A1 => n13052, A2 => n13051, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1991 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => 
                           n13254, B2 => 
                           boothmul_pipelined_i_muxes_in_3_175_port, ZN => 
                           n13054);
   U1992 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => 
                           n13080, B2 => 
                           boothmul_pipelined_i_muxes_in_3_174_port, ZN => 
                           n13053);
   U1993 : NAND2_X1 port map( A1 => n13054, A2 => n13053, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1994 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => 
                           n13254, B2 => 
                           boothmul_pipelined_i_muxes_in_3_174_port, ZN => 
                           n13056);
   U1995 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => 
                           n13080, B2 => 
                           boothmul_pipelined_i_muxes_in_3_173_port, ZN => 
                           n13055);
   U1996 : NAND2_X1 port map( A1 => n13056, A2 => n13055, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1997 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_173_port, ZN => 
                           n13058);
   U1998 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_172_port, ZN => 
                           n13057);
   U1999 : NAND2_X1 port map( A1 => n13058, A2 => n13057, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U2000 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_172_port, ZN => 
                           n13060);
   U2001 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => 
                           n13080, B2 => 
                           boothmul_pipelined_i_muxes_in_3_171_port, ZN => 
                           n13059);
   U2002 : NAND2_X1 port map( A1 => n13060, A2 => n13059, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U2003 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_171_port, ZN => 
                           n13062);
   U2004 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_170_port, ZN => 
                           n13061);
   U2005 : NAND2_X1 port map( A1 => n13062, A2 => n13061, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U2006 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_170_port, ZN => 
                           n13064);
   U2007 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_169_port, ZN => 
                           n13063);
   U2008 : NAND2_X1 port map( A1 => n13064, A2 => n13063, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U2009 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_169_port, ZN => 
                           n13066);
   U2010 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_168_port, ZN => 
                           n13065);
   U2011 : NAND2_X1 port map( A1 => n13066, A2 => n13065, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U2012 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_168_port, ZN => 
                           n13068);
   U2013 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => 
                           n13080, B2 => 
                           boothmul_pipelined_i_muxes_in_3_167_port, ZN => 
                           n13067);
   U2014 : NAND2_X1 port map( A1 => n13068, A2 => n13067, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U2015 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_167_port, ZN => 
                           n13070);
   U2016 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_166_port, ZN => 
                           n13069);
   U2017 : NAND2_X1 port map( A1 => n13070, A2 => n13069, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U2018 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_166_port, ZN => 
                           n13072);
   U2019 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_165_port, ZN => 
                           n13071);
   U2020 : NAND2_X1 port map( A1 => n13072, A2 => n13071, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U2021 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => 
                           n13254, B2 => 
                           boothmul_pipelined_i_muxes_in_3_165_port, ZN => 
                           n13074);
   U2022 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_164_port, ZN => 
                           n13073);
   U2023 : NAND2_X1 port map( A1 => n13074, A2 => n13073, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U2024 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => 
                           n13075, B2 => 
                           boothmul_pipelined_i_muxes_in_3_164_port, ZN => 
                           n13078);
   U2025 : AOI22_X1 port map( A1 => n13076, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => 
                           n13080, B2 => 
                           boothmul_pipelined_i_muxes_in_3_163_port, ZN => 
                           n13077);
   U2026 : NAND2_X1 port map( A1 => n13078, A2 => n13077, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U2027 : AOI22_X1 port map( A1 => n13079, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => 
                           n13254, B2 => 
                           boothmul_pipelined_i_muxes_in_3_163_port, ZN => 
                           n13082);
   U2028 : NAND2_X1 port map( A1 => n13080, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, ZN => 
                           n13081);
   U2029 : OAI211_X1 port map( C1 => n7164, C2 => n13257, A => n13082, B => 
                           n13081, ZN => boothmul_pipelined_i_mux_out_3_21_port
                           );
   U2030 : NAND3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n13241);
   U2031 : NOR3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_8_port, 
                           ZN => n13239);
   U2032 : INV_X1 port map( A => n13239, ZN => n13086);
   U2033 : INV_X1 port map( A => n13084, ZN => n13083);
   U2034 : NAND2_X1 port map( A1 => n3078, A2 => n13083, ZN => n13242);
   U2035 : INV_X1 port map( A => n13242, ZN => n13112);
   U2036 : NOR2_X1 port map( A1 => n3078, A2 => n13084, ZN => n13116);
   U2037 : CLKBUF_X1 port map( A => n13116, Z => n13238);
   U2038 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, ZN => 
                           n13085);
   U2039 : OAI221_X1 port map( B1 => n5121, B2 => n13241, C1 => n5121, C2 => 
                           n13086, A => n13085, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U2040 : INV_X1 port map( A => n13241, ZN => n13115);
   U2041 : CLKBUF_X1 port map( A => n13239, Z => n13111);
   U2042 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_64_port, A2
                           => n13115, B1 => n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, ZN => 
                           n13088);
   U2043 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => 
                           n13116, B2 => 
                           boothmul_pipelined_i_muxes_in_4_189_port, ZN => 
                           n13087);
   U2044 : NAND2_X1 port map( A1 => n13088, A2 => n13087, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U2045 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => 
                           n13239, B2 => 
                           boothmul_pipelined_i_muxes_in_4_189_port, ZN => 
                           n13090);
   U2046 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => 
                           n13116, B2 => 
                           boothmul_pipelined_i_muxes_in_4_188_port, ZN => 
                           n13089);
   U2047 : NAND2_X1 port map( A1 => n13090, A2 => n13089, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U2048 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => 
                           n13239, B2 => 
                           boothmul_pipelined_i_muxes_in_4_188_port, ZN => 
                           n13092);
   U2049 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => 
                           n13116, B2 => 
                           boothmul_pipelined_i_muxes_in_4_187_port, ZN => 
                           n13091);
   U2050 : NAND2_X1 port map( A1 => n13092, A2 => n13091, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U2051 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_187_port, ZN => 
                           n13094);
   U2052 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_186_port, ZN => 
                           n13093);
   U2053 : NAND2_X1 port map( A1 => n13094, A2 => n13093, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U2054 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_186_port, ZN => 
                           n13096);
   U2055 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => 
                           n13116, B2 => 
                           boothmul_pipelined_i_muxes_in_4_185_port, ZN => 
                           n13095);
   U2056 : NAND2_X1 port map( A1 => n13096, A2 => n13095, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U2057 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_185_port, ZN => 
                           n13098);
   U2058 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_184_port, ZN => 
                           n13097);
   U2059 : NAND2_X1 port map( A1 => n13098, A2 => n13097, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U2060 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_184_port, ZN => 
                           n13100);
   U2061 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_183_port, ZN => 
                           n13099);
   U2062 : NAND2_X1 port map( A1 => n13100, A2 => n13099, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U2063 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_183_port, ZN => 
                           n13102);
   U2064 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_182_port, ZN => 
                           n13101);
   U2065 : NAND2_X1 port map( A1 => n13102, A2 => n13101, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U2066 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_182_port, ZN => 
                           n13104);
   U2067 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => 
                           n13116, B2 => 
                           boothmul_pipelined_i_muxes_in_4_181_port, ZN => 
                           n13103);
   U2068 : NAND2_X1 port map( A1 => n13104, A2 => n13103, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U2069 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_181_port, ZN => 
                           n13106);
   U2070 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_180_port, ZN => 
                           n13105);
   U2071 : NAND2_X1 port map( A1 => n13106, A2 => n13105, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U2072 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_180_port, ZN => 
                           n13108);
   U2073 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_179_port, ZN => 
                           n13107);
   U2074 : NAND2_X1 port map( A1 => n13108, A2 => n13107, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U2075 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => 
                           n13239, B2 => 
                           boothmul_pipelined_i_muxes_in_4_179_port, ZN => 
                           n13110);
   U2076 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_178_port, ZN => 
                           n13109);
   U2077 : NAND2_X1 port map( A1 => n13110, A2 => n13109, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U2078 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => 
                           n13111, B2 => 
                           boothmul_pipelined_i_muxes_in_4_178_port, ZN => 
                           n13114);
   U2079 : AOI22_X1 port map( A1 => n13112, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => 
                           n13116, B2 => 
                           boothmul_pipelined_i_muxes_in_4_177_port, ZN => 
                           n13113);
   U2080 : NAND2_X1 port map( A1 => n13114, A2 => n13113, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U2081 : AOI22_X1 port map( A1 => n13115, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => 
                           n13239, B2 => 
                           boothmul_pipelined_i_muxes_in_4_177_port, ZN => 
                           n13118);
   U2082 : NAND2_X1 port map( A1 => n13116, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, ZN => 
                           n13117);
   U2083 : OAI211_X1 port map( C1 => n5127, C2 => n13242, A => n13118, B => 
                           n13117, ZN => boothmul_pipelined_i_mux_out_4_23_port
                           );
   U2084 : NAND3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n13246);
   U2085 : NOR3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_10_port, 
                           ZN => n13244);
   U2086 : INV_X1 port map( A => n13244, ZN => n13122);
   U2087 : INV_X1 port map( A => n13120, ZN => n13119);
   U2088 : NAND2_X1 port map( A1 => n3079, A2 => n13119, ZN => n13247);
   U2089 : INV_X1 port map( A => n13247, ZN => n13148);
   U2090 : NOR2_X1 port map( A1 => n3079, A2 => n13120, ZN => n13152);
   U2091 : CLKBUF_X1 port map( A => n13152, Z => n13243);
   U2092 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_68_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, ZN => 
                           n13121);
   U2093 : OAI221_X1 port map( B1 => n5122, B2 => n13246, C1 => n5122, C2 => 
                           n13122, A => n13121, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2094 : INV_X1 port map( A => n13246, ZN => n13151);
   U2095 : CLKBUF_X1 port map( A => n13244, Z => n13147);
   U2096 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_5_68_port, A2
                           => n13151, B1 => n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, ZN => 
                           n13124);
   U2097 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => 
                           n13152, B2 => 
                           boothmul_pipelined_i_muxes_in_5_203_port, ZN => 
                           n13123);
   U2098 : NAND2_X1 port map( A1 => n13124, A2 => n13123, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2099 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => 
                           n13244, B2 => 
                           boothmul_pipelined_i_muxes_in_5_203_port, ZN => 
                           n13126);
   U2100 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => 
                           n13152, B2 => 
                           boothmul_pipelined_i_muxes_in_5_202_port, ZN => 
                           n13125);
   U2101 : NAND2_X1 port map( A1 => n13126, A2 => n13125, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2102 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => 
                           n13244, B2 => 
                           boothmul_pipelined_i_muxes_in_5_202_port, ZN => 
                           n13128);
   U2103 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => 
                           n13152, B2 => 
                           boothmul_pipelined_i_muxes_in_5_201_port, ZN => 
                           n13127);
   U2104 : NAND2_X1 port map( A1 => n13128, A2 => n13127, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2105 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_201_port, ZN => 
                           n13130);
   U2106 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_200_port, ZN => 
                           n13129);
   U2107 : NAND2_X1 port map( A1 => n13130, A2 => n13129, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2108 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_200_port, ZN => 
                           n13132);
   U2109 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => 
                           n13152, B2 => 
                           boothmul_pipelined_i_muxes_in_5_199_port, ZN => 
                           n13131);
   U2110 : NAND2_X1 port map( A1 => n13132, A2 => n13131, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2111 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_199_port, ZN => 
                           n13134);
   U2112 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_198_port, ZN => 
                           n13133);
   U2113 : NAND2_X1 port map( A1 => n13134, A2 => n13133, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2114 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_198_port, ZN => 
                           n13136);
   U2115 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_197_port, ZN => 
                           n13135);
   U2116 : NAND2_X1 port map( A1 => n13136, A2 => n13135, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2117 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_197_port, ZN => 
                           n13138);
   U2118 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_196_port, ZN => 
                           n13137);
   U2119 : NAND2_X1 port map( A1 => n13138, A2 => n13137, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2120 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_196_port, ZN => 
                           n13140);
   U2121 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => 
                           n13152, B2 => 
                           boothmul_pipelined_i_muxes_in_5_195_port, ZN => 
                           n13139);
   U2122 : NAND2_X1 port map( A1 => n13140, A2 => n13139, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2123 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_195_port, ZN => 
                           n13142);
   U2124 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_194_port, ZN => 
                           n13141);
   U2125 : NAND2_X1 port map( A1 => n13142, A2 => n13141, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2126 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_194_port, ZN => 
                           n13144);
   U2127 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_193_port, ZN => 
                           n13143);
   U2128 : NAND2_X1 port map( A1 => n13144, A2 => n13143, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2129 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => 
                           n13244, B2 => 
                           boothmul_pipelined_i_muxes_in_5_193_port, ZN => 
                           n13146);
   U2130 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_192_port, ZN => 
                           n13145);
   U2131 : NAND2_X1 port map( A1 => n13146, A2 => n13145, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2132 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => 
                           n13147, B2 => 
                           boothmul_pipelined_i_muxes_in_5_192_port, ZN => 
                           n13150);
   U2133 : AOI22_X1 port map( A1 => n13148, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => 
                           n13152, B2 => 
                           boothmul_pipelined_i_muxes_in_5_191_port, ZN => 
                           n13149);
   U2134 : NAND2_X1 port map( A1 => n13150, A2 => n13149, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2135 : AOI22_X1 port map( A1 => n13151, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => 
                           n13244, B2 => 
                           boothmul_pipelined_i_muxes_in_5_191_port, ZN => 
                           n13154);
   U2136 : NAND2_X1 port map( A1 => n13152, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, ZN => 
                           n13153);
   U2137 : OAI211_X1 port map( C1 => n5128, C2 => n13247, A => n13154, B => 
                           n13153, ZN => boothmul_pipelined_i_mux_out_5_25_port
                           );
   U2138 : NAND3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n13251);
   U2139 : NOR3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_12_port, 
                           ZN => n13249);
   U2140 : INV_X1 port map( A => n13249, ZN => n13158);
   U2141 : INV_X1 port map( A => n13156, ZN => n13155);
   U2142 : NAND2_X1 port map( A1 => n3080, A2 => n13155, ZN => n13252);
   U2143 : INV_X1 port map( A => n13252, ZN => n13184);
   U2144 : NOR2_X1 port map( A1 => n3080, A2 => n13156, ZN => n13188);
   U2145 : CLKBUF_X1 port map( A => n13188, Z => n13248);
   U2146 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_72_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, ZN => 
                           n13157);
   U2147 : OAI221_X1 port map( B1 => n5123, B2 => n13251, C1 => n5123, C2 => 
                           n13158, A => n13157, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2148 : INV_X1 port map( A => n13251, ZN => n13187);
   U2149 : CLKBUF_X1 port map( A => n13249, Z => n13183);
   U2150 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_6_72_port, A2
                           => n13187, B1 => n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, ZN => 
                           n13160);
   U2151 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => 
                           n13188, B2 => 
                           boothmul_pipelined_i_muxes_in_6_217_port, ZN => 
                           n13159);
   U2152 : NAND2_X1 port map( A1 => n13160, A2 => n13159, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2153 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => 
                           n13249, B2 => 
                           boothmul_pipelined_i_muxes_in_6_217_port, ZN => 
                           n13162);
   U2154 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => 
                           n13188, B2 => 
                           boothmul_pipelined_i_muxes_in_6_216_port, ZN => 
                           n13161);
   U2155 : NAND2_X1 port map( A1 => n13162, A2 => n13161, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2156 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => 
                           n13249, B2 => 
                           boothmul_pipelined_i_muxes_in_6_216_port, ZN => 
                           n13164);
   U2157 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => 
                           n13188, B2 => 
                           boothmul_pipelined_i_muxes_in_6_215_port, ZN => 
                           n13163);
   U2158 : NAND2_X1 port map( A1 => n13164, A2 => n13163, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2159 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_215_port, ZN => 
                           n13166);
   U2160 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_214_port, ZN => 
                           n13165);
   U2161 : NAND2_X1 port map( A1 => n13166, A2 => n13165, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2162 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_214_port, ZN => 
                           n13168);
   U2163 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => 
                           n13188, B2 => 
                           boothmul_pipelined_i_muxes_in_6_213_port, ZN => 
                           n13167);
   U2164 : NAND2_X1 port map( A1 => n13168, A2 => n13167, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2165 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_213_port, ZN => 
                           n13170);
   U2166 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_212_port, ZN => 
                           n13169);
   U2167 : NAND2_X1 port map( A1 => n13170, A2 => n13169, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2168 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_212_port, ZN => 
                           n13172);
   U2169 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_211_port, ZN => 
                           n13171);
   U2170 : NAND2_X1 port map( A1 => n13172, A2 => n13171, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2171 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_211_port, ZN => 
                           n13174);
   U2172 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_210_port, ZN => 
                           n13173);
   U2173 : NAND2_X1 port map( A1 => n13174, A2 => n13173, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2174 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_210_port, ZN => 
                           n13176);
   U2175 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => 
                           n13188, B2 => 
                           boothmul_pipelined_i_muxes_in_6_209_port, ZN => 
                           n13175);
   U2176 : NAND2_X1 port map( A1 => n13176, A2 => n13175, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2177 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_209_port, ZN => 
                           n13178);
   U2178 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_208_port, ZN => 
                           n13177);
   U2179 : NAND2_X1 port map( A1 => n13178, A2 => n13177, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2180 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_208_port, ZN => 
                           n13180);
   U2181 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_207_port, ZN => 
                           n13179);
   U2182 : NAND2_X1 port map( A1 => n13180, A2 => n13179, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2183 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => 
                           n13249, B2 => 
                           boothmul_pipelined_i_muxes_in_6_207_port, ZN => 
                           n13182);
   U2184 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_206_port, ZN => 
                           n13181);
   U2185 : NAND2_X1 port map( A1 => n13182, A2 => n13181, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2186 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => 
                           n13183, B2 => 
                           boothmul_pipelined_i_muxes_in_6_206_port, ZN => 
                           n13186);
   U2187 : AOI22_X1 port map( A1 => n13184, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => 
                           n13188, B2 => 
                           boothmul_pipelined_i_muxes_in_6_205_port, ZN => 
                           n13185);
   U2188 : NAND2_X1 port map( A1 => n13186, A2 => n13185, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2189 : AOI22_X1 port map( A1 => n13187, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => 
                           n13249, B2 => 
                           boothmul_pipelined_i_muxes_in_6_205_port, ZN => 
                           n13190);
   U2190 : NAND2_X1 port map( A1 => n13188, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, ZN => 
                           n13189);
   U2191 : OAI211_X1 port map( C1 => n5129, C2 => n13252, A => n13190, B => 
                           n13189, ZN => boothmul_pipelined_i_mux_out_6_27_port
                           );
   U2192 : NOR2_X1 port map( A1 => n13191, A2 => n13258, ZN => n13208);
   U2193 : INV_X1 port map( A => n13208, ZN => n13195);
   U2194 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A3 => n7165, ZN => n13231);
   U2195 : INV_X1 port map( A => n13231, ZN => n13194);
   U2196 : NOR2_X1 port map( A1 => n13192, A2 => n13258, ZN => n13225);
   U2197 : CLKBUF_X1 port map( A => n13225, Z => n13229);
   U2198 : NOR2_X1 port map( A1 => n7165, A2 => n13192, ZN => n13209);
   U2199 : CLKBUF_X1 port map( A => n13209, Z => n13230);
   U2200 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_76_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, ZN => 
                           n13193);
   U2201 : OAI221_X1 port map( B1 => n5134, B2 => n13195, C1 => n5134, C2 => 
                           n13194, A => n13193, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2202 : CLKBUF_X1 port map( A => n13231, Z => n13224);
   U2203 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_7_76_port, A2
                           => n13208, B1 => n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, ZN => 
                           n13197);
   U2204 : AOI22_X1 port map( A1 => n13225, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => 
                           n13209, B2 => 
                           boothmul_pipelined_i_muxes_in_7_231_port, ZN => 
                           n13196);
   U2205 : NAND2_X1 port map( A1 => n13197, A2 => n13196, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2206 : CLKBUF_X1 port map( A => n13208, Z => n13228);
   U2207 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => 
                           n13231, B2 => 
                           boothmul_pipelined_i_muxes_in_7_231_port, ZN => 
                           n13199);
   U2208 : AOI22_X1 port map( A1 => n13225, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => 
                           n13209, B2 => 
                           boothmul_pipelined_i_muxes_in_7_230_port, ZN => 
                           n13198);
   U2209 : NAND2_X1 port map( A1 => n13199, A2 => n13198, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2210 : AOI22_X1 port map( A1 => n13208, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => 
                           n13231, B2 => 
                           boothmul_pipelined_i_muxes_in_7_230_port, ZN => 
                           n13201);
   U2211 : AOI22_X1 port map( A1 => n13225, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => 
                           n13209, B2 => 
                           boothmul_pipelined_i_muxes_in_7_229_port, ZN => 
                           n13200);
   U2212 : NAND2_X1 port map( A1 => n13201, A2 => n13200, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2213 : AOI22_X1 port map( A1 => n13208, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_229_port, ZN => 
                           n13203);
   U2214 : AOI22_X1 port map( A1 => n13225, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => 
                           n13209, B2 => 
                           boothmul_pipelined_i_muxes_in_7_228_port, ZN => 
                           n13202);
   U2215 : NAND2_X1 port map( A1 => n13203, A2 => n13202, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2216 : AOI22_X1 port map( A1 => n13208, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_228_port, ZN => 
                           n13205);
   U2217 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => 
                           n13209, B2 => 
                           boothmul_pipelined_i_muxes_in_7_227_port, ZN => 
                           n13204);
   U2218 : NAND2_X1 port map( A1 => n13205, A2 => n13204, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2219 : AOI22_X1 port map( A1 => n13208, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_227_port, ZN => 
                           n13207);
   U2220 : AOI22_X1 port map( A1 => n13225, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => 
                           n13209, B2 => 
                           boothmul_pipelined_i_muxes_in_7_226_port, ZN => 
                           n13206);
   U2221 : NAND2_X1 port map( A1 => n13207, A2 => n13206, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2222 : AOI22_X1 port map( A1 => n13208, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_226_port, ZN => 
                           n13211);
   U2223 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => 
                           n13209, B2 => 
                           boothmul_pipelined_i_muxes_in_7_225_port, ZN => 
                           n13210);
   U2224 : NAND2_X1 port map( A1 => n13211, A2 => n13210, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2225 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_225_port, ZN => 
                           n13213);
   U2226 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_224_port, ZN => 
                           n13212);
   U2227 : NAND2_X1 port map( A1 => n13213, A2 => n13212, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2228 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => 
                           n13231, B2 => 
                           boothmul_pipelined_i_muxes_in_7_224_port, ZN => 
                           n13215);
   U2229 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_223_port, ZN => 
                           n13214);
   U2230 : NAND2_X1 port map( A1 => n13215, A2 => n13214, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2231 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_223_port, ZN => 
                           n13217);
   U2232 : AOI22_X1 port map( A1 => n13225, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_222_port, ZN => 
                           n13216);
   U2233 : NAND2_X1 port map( A1 => n13217, A2 => n13216, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2234 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_222_port, ZN => 
                           n13219);
   U2235 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_221_port, ZN => 
                           n13218);
   U2236 : NAND2_X1 port map( A1 => n13219, A2 => n13218, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2237 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_221_port, ZN => 
                           n13221);
   U2238 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_220_port, ZN => 
                           n13220);
   U2239 : NAND2_X1 port map( A1 => n13221, A2 => n13220, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2240 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => 
                           n13231, B2 => 
                           boothmul_pipelined_i_muxes_in_7_220_port, ZN => 
                           n13223);
   U2241 : AOI22_X1 port map( A1 => n13229, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_219_port, ZN => 
                           n13222);
   U2242 : NAND2_X1 port map( A1 => n13223, A2 => n13222, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2243 : AOI22_X1 port map( A1 => n13228, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => 
                           n13224, B2 => 
                           boothmul_pipelined_i_muxes_in_7_219_port, ZN => 
                           n13227);
   U2244 : AOI22_X1 port map( A1 => n13225, A2 => 
                           boothmul_pipelined_i_muxes_in_7_62_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, ZN => 
                           n13226);
   U2245 : NAND2_X1 port map( A1 => n13227, A2 => n13226, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2246 : OAI21_X1 port map( B1 => n13229, B2 => n13228, A => 
                           boothmul_pipelined_i_muxes_in_7_62_port, ZN => 
                           n13233);
   U2247 : AOI22_X1 port map( A1 => n13231, A2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, B1 => 
                           n13230, B2 => 
                           boothmul_pipelined_i_muxes_in_7_217_port, ZN => 
                           n13232);
   U2248 : NAND2_X1 port map( A1 => n13233, A2 => n13232, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2249 : AOI22_X1 port map( A1 => n13235, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n13234, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n13236);
   U2250 : OAI21_X1 port map( B1 => n13237, B2 => n1976, A => n13236, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2251 : AOI22_X1 port map( A1 => n13239, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, B1 => 
                           n13238, B2 => 
                           boothmul_pipelined_i_muxes_in_4_175_port, ZN => 
                           n13240);
   U2252 : OAI221_X1 port map( B1 => n5127, B2 => n13242, C1 => n5127, C2 => 
                           n13241, A => n13240, ZN => n1997);
   U2253 : AOI22_X1 port map( A1 => n13244, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, B1 => 
                           n13243, B2 => 
                           boothmul_pipelined_i_muxes_in_5_189_port, ZN => 
                           n13245);
   U2254 : OAI221_X1 port map( B1 => n5128, B2 => n13247, C1 => n5128, C2 => 
                           n13246, A => n13245, ZN => n1996);
   U2255 : AOI22_X1 port map( A1 => n13249, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, B1 => 
                           n13248, B2 => 
                           boothmul_pipelined_i_muxes_in_6_203_port, ZN => 
                           n13250);
   U2256 : OAI221_X1 port map( B1 => n5129, B2 => n13252, C1 => n5129, C2 => 
                           n13251, A => n13250, ZN => n1995);
   U2257 : AOI22_X1 port map( A1 => n13254, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, B1 => 
                           n13253, B2 => 
                           boothmul_pipelined_i_muxes_in_3_161_port, ZN => 
                           n13255);
   U2258 : OAI221_X1 port map( B1 => n7164, B2 => n13257, C1 => n7164, C2 => 
                           n13256, A => n13255, ZN => n1991);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N385, N386, N387, N388, N389, N390, N391, N392, N393
      , N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, 
      n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, 
      n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, 
      n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, 
      n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, 
      n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, 
      n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, 
      n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, 
      n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, 
      n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, 
      n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, 
      n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, 
      n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, 
      n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, 
      n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, 
      n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, 
      n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, 
      n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, 
      n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, 
      n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, 
      n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, 
      n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, 
      n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, 
      n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, 
      n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, 
      n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, 
      n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, 
      n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, 
      n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, 
      n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, 
      n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, 
      n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, 
      n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, 
      n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, 
      n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, 
      n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, 
      n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, 
      n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, 
      n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, 
      n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, 
      n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, 
      n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, 
      n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, 
      n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, 
      n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, 
      n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, 
      n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, 
      n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, 
      n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, 
      n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, 
      n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, 
      n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, 
      n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, 
      n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, 
      n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, 
      n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, 
      n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, 
      n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, 
      n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, 
      n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, 
      n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, 
      n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, 
      n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, 
      n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, 
      n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, 
      n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, 
      n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, 
      n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, 
      n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, 
      n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, 
      n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, 
      n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, 
      n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, 
      n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, 
      n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, 
      n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, 
      n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, 
      n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, 
      n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, 
      n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, 
      n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, 
      n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, 
      n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, 
      n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, 
      n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, 
      n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, 
      n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, 
      n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, 
      n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, 
      n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, 
      n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, 
      n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, 
      n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, 
      n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, 
      n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, 
      n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, 
      n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, 
      n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, 
      n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, 
      n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, 
      n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, 
      n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, 
      n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, 
      n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, 
      n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, 
      n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, 
      n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, 
      n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, 
      n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, 
      n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, 
      n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, 
      n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, 
      n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, 
      n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, 
      n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, 
      n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, 
      n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, 
      n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, 
      n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, 
      n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, 
      n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, 
      n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, 
      n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, 
      n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, 
      n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, 
      n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, 
      n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, 
      n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, 
      n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, 
      n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, 
      n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, 
      n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, 
      n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, 
      n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, 
      n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, 
      n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, 
      n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, 
      n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, 
      n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, 
      n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, 
      n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, 
      n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, 
      n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, 
      n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, 
      n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, 
      n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, 
      n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, 
      n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, 
      n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, 
      n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, 
      n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, 
      n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, 
      n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, 
      n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, 
      n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, 
      n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, 
      n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, 
      n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, 
      n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, 
      n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, 
      n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, 
      n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, 
      n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, 
      n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, 
      n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, 
      n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, 
      n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, 
      n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, 
      n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, 
      n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, 
      n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, 
      n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, 
      n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, 
      n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, 
      n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, 
      n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, 
      n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, 
      n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, 
      n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, 
      n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, 
      n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, 
      n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, 
      n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, 
      n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, 
      n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, 
      n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, 
      n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, 
      n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, 
      n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, 
      n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, 
      n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, 
      n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, 
      n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, 
      n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, 
      n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, 
      n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, 
      n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, 
      n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, 
      n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, 
      n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, 
      n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, 
      n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, 
      n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, 
      n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, 
      n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, 
      n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, 
      n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, 
      n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, 
      n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, 
      n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, 
      n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, 
      n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, 
      n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, 
      n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, 
      n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, 
      n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, 
      n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, 
      n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, 
      n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, 
      n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, 
      n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, 
      n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, 
      n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, 
      n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, 
      n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, 
      n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, 
      n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, 
      n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, 
      n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, 
      n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, 
      n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, 
      n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, 
      n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, 
      n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, 
      n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, 
      n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, 
      n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, 
      n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, 
      n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, 
      n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, 
      n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, 
      n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, 
      n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, 
      n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, 
      n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, 
      n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, 
      n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, 
      n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, 
      n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, 
      n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, 
      n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, 
      n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, 
      n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, 
      n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, 
      n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, 
      n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, 
      n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, 
      n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, 
      n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, 
      n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, 
      n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, 
      n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, 
      n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, 
      n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, 
      n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, 
      n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, 
      n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, 
      n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, 
      n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, 
      n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, 
      n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, 
      n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, 
      n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, 
      n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, 
      n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, 
      n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, 
      n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, 
      n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, 
      n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, 
      n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, 
      n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, 
      n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, 
      n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, 
      n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, 
      n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, 
      n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, 
      n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, 
      n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, 
      n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, 
      n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, 
      n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, 
      n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, 
      n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, 
      n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, 
      n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, 
      n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, 
      n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, 
      n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, 
      n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, 
      n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, 
      n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, 
      n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, 
      n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, 
      n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, 
      n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, 
      n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, 
      n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, 
      n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, 
      n19552, n19553, n19554, n19555, n_1349, n_1350, n_1351, n_1352, n_1353, 
      n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, 
      n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, 
      n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, 
      n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, 
      n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, 
      n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, 
      n_1408, n_1409, n_1410, n_1411, n_1412 : std_logic;

begin
   
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n18539);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n18795);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n19053);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n18540);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n18796);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n18541);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n18797);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n18798);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n18799);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n18800);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n19306);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n18542);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n18543);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n18801);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n18544);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n19307);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n18545);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n18802);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n18546);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n18803);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n18804);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n18547);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n19308);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n18805);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n19054);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n19055);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n18548);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n19309);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n19056);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n18806);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           REGISTERS_1_28_port, QN => n19310);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n18549);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n19057);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n18550);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n18807);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n18808);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n18551);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n19058);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n19311);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n19059);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n19312);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n19060);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n18809);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n18552);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n19061);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n19313);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n18553);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n19062);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n18554);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n19314);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n19315);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n19063);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n19316);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n18810);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n18811);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n18555);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n18812);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n19317);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n19064);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n18813);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n18814);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n18556);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n18557);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n18558);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n18559);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n19318);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n18815);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n19319);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n18560);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n18816);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n18561);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n18817);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n18562);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n19065);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n18563);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n19320);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n18818);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n18819);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n18820);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n18821);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n18564);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n18565);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n18566);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n18822);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n18567);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n18823);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n18824);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n18825);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n18568);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n18569);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n18826);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n19321);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n18570);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n19322);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n18827);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n18828);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n19066);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n18571);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n19323);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n18572);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n19067);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n18573);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n19068);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n18574);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n18575);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n18576);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n18577);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n19069);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n19324);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n18578);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n19325);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n18579);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n19326);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n18829);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n18830);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n18831);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n19070);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n19071);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n19327);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n19072);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n18580);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n18581);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n18582);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n19073);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n19328);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n19329);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n19074);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n19330);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n18832);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n19075);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n19331);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n19076);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n19332);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n19077);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n19078);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n19333);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n19079);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n18833);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n19080);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n19334);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n19081);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n19082);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n19335);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n19083);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n19336);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n19084);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n19337);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n19338);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n19085);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n19086);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n18583);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n19087);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n19088);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n18834);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n19339);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n18835);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n18584);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n19340);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n19341);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n19342);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n19343);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n19089);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n18585);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n19344);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n19090);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n19345);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n18836);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n19346);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n19091);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n19347);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           REGISTERS_5_16_port, QN => n19348);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n18837);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n18586);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n19092);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n19093);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n18838);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n19349);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n19094);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n19095);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n19096);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n18587);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n19350);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n19097);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n19098);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n19351);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n19099);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n19352);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n19100);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n19101);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n19102);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n19103);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n19104);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n19353);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n19354);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n19105);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n19106);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n19355);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n19356);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n19357);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n19107);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n19358);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n19359);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n19360);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n19361);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n19362);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n19108);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n19109);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n19363);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n19110);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n19111);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n19112);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n19113);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n19364);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n19365);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n19114);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n19366);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n19367);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n19368);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n19115);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n18588);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n18839);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n18589);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n18590);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n18840);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n18841);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n18842);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n18591);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n18843);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n18844);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n18845);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n18592);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n18593);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n18846);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n18594);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n18595);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n18596);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n18847);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n18848);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n18849);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n18597);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n18850);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n18851);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n18852);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n18598);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n18853);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n18599);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n18600);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n18854);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n18855);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n18856);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n18857);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n18858);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n19116);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n18601);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n18602);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n19117);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n18859);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n18603);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n18604);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n18605);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n18606);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n18860);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n19369);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n18607);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n18608);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n19118);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n18609);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n19119);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n18610);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n19120);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n19121);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n18611);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n18861);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n18612);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n19122);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n19370);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n18613);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n19371);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n18614);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n19123);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n18615);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n18616);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n18617);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n19372);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n19373);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n19374);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n18862);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n19124);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n19125);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n19126);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n19375);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n19127);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n19376);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n18618);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n18863);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n18619);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n18864);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n19377);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n19128);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n19378);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n19379);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n18865);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n19129);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n19130);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n18620);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n19380);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n18621);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n19131);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n18866);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n18867);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n19381);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n19382);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n19383);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n18622);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n18623);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n19132);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n18624);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n18625);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n18868);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n18626);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n18869);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n18870);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n18627);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n18871);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n18628);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n18629);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n18872);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n19133);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n18873);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n18630);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n18874);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n18631);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n18632);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           REGISTERS_10_13_port, QN => n18875);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n18876);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n18633);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n18634);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n18635);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           REGISTERS_10_8_port, QN => n18636);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n18877);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n18878);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n18637);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n18638);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n18639);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n18879);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n18880);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n18881);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n18882);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n18883);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n19384);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n19134);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n18884);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n18640);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n18885);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n18886);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n19135);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n19136);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n19385);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n18641);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n19386);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n19137);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n18887);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n18888);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n18889);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n19387);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n19138);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n18642);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n19388);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n19139);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n18890);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n18891);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n18892);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n19140);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n18893);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n19389);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n18894);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n18643);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n19141);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n19142);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n18644);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n19390);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n18895);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n19143);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n19391);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n19144);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n19392);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n19393);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n19394);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n18896);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n19395);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n19145);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n19146);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n19396);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n18897);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n19397);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n18645);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n18898);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n18646);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           REGISTERS_12_12_port, QN => n18899);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n18900);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n19147);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n19148);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n19398);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n19149);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n19399);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n19150);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n18647);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n18648);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n19151);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n19152);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n19400);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n19153);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n18649);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n19154);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n19155);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n18901);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n19401);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n19156);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n19157);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n18902);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n19402);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n19403);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n19404);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n18903);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n19405);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n19158);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n19159);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n19406);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n19160);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n19407);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n19161);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n19162);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n19408);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n19409);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n19163);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n18650);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n19410);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n19411);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n19412);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n19164);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n19413);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n19414);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n19415);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n19416);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n19165);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n19166);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n19417);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n19418);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n19167);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n19168);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n19419);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n19169);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n19420);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n19170);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n19171);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n19421);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n19172);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n19173);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n19174);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n19175);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n19176);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n19177);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n19422);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n19423);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n19424);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n19425);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n19426);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n19178);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n19179);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n19180);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n19181);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n19427);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n19182);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n19428);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n19183);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n18651);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n18904);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n18905);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n18906);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n18652);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n18907);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n18908);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n18653);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n18909);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n18654);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n18655);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n18656);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n18910);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n18657);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n18911);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n18912);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n18913);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n18914);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n18915);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n18916);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n18917);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n18918);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n18658);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n18919);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n18920);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n18659);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n18660);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n18921);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n18922);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n18923);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n18924);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n18925);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n18788);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n19429);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n19184);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n18926);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n19185);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n19430);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n19431);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n19432);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n18927);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n18661);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n19186);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n19433);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n18662);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n19187);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n18928);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n18929);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n19188);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n19189);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n19434);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n19190);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n18663);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n19435);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n18930);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n19191);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n19436);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n18664);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n19437);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n18665);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n19192);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n18931);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n18932);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n18933);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n18532);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n18934);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n18666);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n18935);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n19438);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           REGISTERS_17_26_port, QN => n18667);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n18936);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n19193);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n19194);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n18937);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n19439);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n19195);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n19196);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n19440);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n19197);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n18668);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n18669);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n19198);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n19199);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n19200);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n18670);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n18938);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n18939);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n19441);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n19442);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n19443);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n18940);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n19201);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n19444);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n18941);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n19445);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n18942);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n18533);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n18671);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n18672);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n18673);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n18674);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n19202);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n19446);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n18943);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n18675);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n19447);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n18944);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n18676);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n19448);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n18677);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n18945);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n19449);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n19450);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n19451);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n18678);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n18679);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n19452);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n19453);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n18680);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n18681);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n18946);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n18682);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n18683);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n19203);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n18947);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n19454);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           REGISTERS_18_1_port, QN => n18948);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n18684);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n18534);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n19204);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n18685);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n19205);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n18686);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n18687);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n18688);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n19206);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n18689);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n18690);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n18691);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n19455);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n18692);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n18693);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n18694);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n19207);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n18949);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n18695);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n18696);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n19208);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n19456);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n18950);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n19457);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n18951);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n19458);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n19459);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n19209);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n18952);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n19460);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n18697);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n19210);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n18698);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n18789);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n19461);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n18699);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n19462);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n19463);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n18700);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n18953);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n18701);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n18954);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n18702);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n19464);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n18955);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n19211);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n19212);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           REGISTERS_20_17_port, QN => n19213);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n19465);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n19214);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n19215);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n19216);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n19466);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n19217);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n19467);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n18956);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n18703);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n19218);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n19219);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n19468);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n19220);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n18704);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n19469);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n19221);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n19222);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n18790);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n19223);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n19470);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n19471);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n19224);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n19225);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n19226);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n19227);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n19472);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n19473);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n19474);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n19475);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n18957);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n19476);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n19477);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n19478);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n19479);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n19480);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n19228);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n19481);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n19229);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n19230);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n19231);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n19482);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n19232);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n18705);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n19483);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n19233);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n19234);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n19484);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n18706);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n19485);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n19047);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n19486);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n19487);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n19235);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n19236);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n19488);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n19237);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n19489);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n19490);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n19491);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n19492);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n19493);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n19494);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n19238);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n19239);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n19240);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n19495);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n19496);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n19497);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n19241);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n19242);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n19243);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n19244);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n19245);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n19498);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n19499);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n19246);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n19500);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n19501);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n19502);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n19247);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n19503);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n19048);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n19248);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n18958);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n18707);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n18959);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n18960);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n18961);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n18962);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n19504);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n18963);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n18708);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n18964);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n18965);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           REGISTERS_23_18_port, QN => n19505);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n19249);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n19506);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n18966);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n18709);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n19507);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n18710);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n18967);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n18711);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n18968);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n18969);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n18712);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n18970);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n18971);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n18713);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n19508);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n18972);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n18973);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n18714);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n18791);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n18974);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n18715);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n18975);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n18976);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n18977);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n18716);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n18717);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n18718);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n18978);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n18979);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n18980);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n18981);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n18982);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n18719);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n18983);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n18984);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n18985);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n18720);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n18986);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n18987);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n19250);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n18721);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n18722);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n18723);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n19509);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n18724);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n18725);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n18726);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n18727);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n18728);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n18988);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n18792);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n18729);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n19251);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n19252);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n19253);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n19510);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n19254);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n19511);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n19255);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n19256);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n18989);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n19257);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n19512);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n18730);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n19258);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n18731);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n19259);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n19260);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n19513);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n18990);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n18991);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n18992);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n19261);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n19514);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n19262);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n19263);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n19515);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n19516);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n19264);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n19265);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n19517);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n19518);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n18793);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n18993);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n19519);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n19520);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n18994);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n19521);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n19522);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n19523);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n19266);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n19267);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n18732);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n18733);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n19268);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n19269);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n18995);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n18734);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n19270);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n18735);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n18996);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n19271);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n19524);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n19272);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n19525);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n19273);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n18736);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n18737);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n18997);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n19526);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n18738);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n19274);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n18998);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n19527);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n19049);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n19528);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n19529);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n19275);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n19530);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n19531);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n19276);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n18739);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n19532);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n19533);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n19277);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n19534);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n19278);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n18999);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n19535);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n19536);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n18740);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n19537);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           REGISTERS_27_13_port, QN => n18741);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n19000);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n19279);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n18742);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n19280);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n19538);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n19281);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n19282);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n19283);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n19539);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n18743);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n19284);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n19285);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n19286);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n19050);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n19540);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n19541);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n18744);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n19287);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n19288);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n19289);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n19290);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n19291);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n19292);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n19293);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n19294);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n19295);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n19296);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n19542);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n19297);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n18745);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n19001);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n19002);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n19543);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n19544);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n19545);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n19298);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n19546);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n19003);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n19299);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n18746);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n19004);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n19547);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n19300);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n19301);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n19548);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n18535);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n18747);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n19005);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n18748);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n19006);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n19007);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n19008);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n19009);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           REGISTERS_29_23_port, QN => n19010);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n18749);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n19011);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n18750);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n18751);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n19012);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n19013);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n19014);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n18752);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n19015);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n19016);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n19017);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n19018);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n18753);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n18754);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n18755);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n19019);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n19020);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n18756);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n19021);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n19022);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n18757);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n19023);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n18758);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n19051);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n18759);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n19549);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n19550);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n18760);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n18761);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n18762);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n19024);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n18763);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n19302);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n19303);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           REGISTERS_30_20_port, QN => n18764);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n19025);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n19026);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n19027);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n18765);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n19551);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n19028);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n19552);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n18766);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n18767);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n18768);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n19553);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n19029);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n19030);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n19031);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n18769);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n19032);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n18770);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n19033);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n19554);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n18771);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n18536);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n18772);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n18773);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n19034);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n19035);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n18774);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n19036);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n18775);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n19037);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n19038);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n18776);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n18777);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n19039);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n19040);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n18778);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n18779);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n19041);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n18780);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n18781);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n19042);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n18782);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n19043);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n19044);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n18783);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n18784);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n19045);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n19555);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n18785);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n19046);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n18786);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n18787);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n19304);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT1(31), QN 
                           => n_1349);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT1(30), QN 
                           => n_1350);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT1(29), QN 
                           => n_1351);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT1(28), QN 
                           => n_1352);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT1(27), QN 
                           => n_1353);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT1(26), QN 
                           => n_1354);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT1(25), QN 
                           => n_1355);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT1(24), QN 
                           => n_1356);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT1(23), QN 
                           => n_1357);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => CLK, Q => OUT1(22), QN 
                           => n_1358);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => CLK, Q => OUT1(21), QN 
                           => n_1359);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => CLK, Q => OUT1(20), QN 
                           => n_1360);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => CLK, Q => OUT1(19), QN 
                           => n_1361);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => CLK, Q => OUT1(18), QN 
                           => n_1362);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => CLK, Q => OUT1(17), QN 
                           => n_1363);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => CLK, Q => OUT1(16), QN 
                           => n_1364);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => CLK, Q => OUT1(15), QN 
                           => n_1365);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => CLK, Q => OUT1(14), QN 
                           => n_1366);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => CLK, Q => OUT1(13), QN 
                           => n_1367);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => CLK, Q => OUT1(12), QN 
                           => n_1368);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => CLK, Q => OUT1(11), QN 
                           => n_1369);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => CLK, Q => OUT1(10), QN 
                           => n_1370);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => CLK, Q => OUT1(9), QN =>
                           n_1371);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => CLK, Q => OUT1(8), QN =>
                           n_1372);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => CLK, Q => OUT1(7), QN =>
                           n_1373);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => CLK, Q => OUT1(6), QN =>
                           n_1374);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => CLK, Q => OUT1(5), QN =>
                           n_1375);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => CLK, Q => OUT1(4), QN =>
                           n_1376);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => CLK, Q => OUT1(3), QN =>
                           n_1377);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => CLK, Q => OUT1(2), QN =>
                           n_1378);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => CLK, Q => OUT1(1), QN =>
                           n_1379);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT2(31), QN 
                           => n_1380);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT2(30), QN 
                           => n_1381);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT2(29), QN 
                           => n_1382);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT2(28), QN 
                           => n_1383);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT2(27), QN 
                           => n_1384);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT2(26), QN 
                           => n_1385);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT2(25), QN 
                           => n_1386);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT2(24), QN 
                           => n_1387);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT2(23), QN 
                           => n_1388);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(22), QN 
                           => n_1389);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(21), QN 
                           => n_1390);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(20), QN 
                           => n_1391);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(19), QN 
                           => n_1392);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(18), QN 
                           => n_1393);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(17), QN 
                           => n_1394);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(16), QN 
                           => n_1395);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(15), QN 
                           => n_1396);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(14), QN 
                           => n_1397);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(13), QN 
                           => n_1398);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(12), QN 
                           => n_1399);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(11), QN 
                           => n_1400);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(10), QN 
                           => n_1401);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(9), QN =>
                           n_1402);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(8), QN =>
                           n_1403);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(7), QN =>
                           n_1404);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(6), QN =>
                           n_1405);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(5), QN =>
                           n_1406);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(4), QN =>
                           n_1407);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(3), QN =>
                           n_1408);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(2), QN =>
                           n_1409);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(1), QN =>
                           n_1410);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(0), QN =>
                           n_1411);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => CLK, Q => OUT1(0), QN =>
                           n_1412);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n18537);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n19305);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n18538);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n18794);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n19052);
   U3 : CLKBUF_X1 port map( A => RESET_BAR, Z => n16780);
   U4 : CLKBUF_X1 port map( A => RESET_BAR, Z => n16781);
   U5 : CLKBUF_X1 port map( A => RESET_BAR, Z => n16782);
   U6 : CLKBUF_X1 port map( A => RESET_BAR, Z => n16783);
   U7 : NAND2_X2 port map( A1 => n16780, A2 => n16956, ZN => n16968);
   U8 : NAND2_X2 port map( A1 => n16783, A2 => n16929, ZN => n16931);
   U9 : NAND2_X2 port map( A1 => n16780, A2 => n16920, ZN => n16922);
   U10 : NAND2_X2 port map( A1 => n16780, A2 => n16916, ZN => n16918);
   U11 : NAND2_X2 port map( A1 => n16781, A2 => n16912, ZN => n16914);
   U12 : NAND2_X2 port map( A1 => n16780, A2 => n16903, ZN => n16905);
   U13 : NAND2_X2 port map( A1 => n16780, A2 => n16839, ZN => n16841);
   U14 : NAND2_X2 port map( A1 => n16781, A2 => n16831, ZN => n16833);
   U15 : NAND2_X2 port map( A1 => n16780, A2 => n16828, ZN => n16830);
   U16 : NAND2_X2 port map( A1 => n16780, A2 => n16825, ZN => n16827);
   U17 : NAND2_X2 port map( A1 => n16780, A2 => n16822, ZN => n16824);
   U18 : NAND2_X2 port map( A1 => n16783, A2 => n16819, ZN => n16821);
   U19 : NAND2_X2 port map( A1 => n16780, A2 => n16816, ZN => n16818);
   U20 : NAND2_X2 port map( A1 => n16783, A2 => n16897, ZN => n16899);
   U21 : NAND2_X2 port map( A1 => n16783, A2 => n16892, ZN => n16894);
   U22 : NAND2_X2 port map( A1 => n16783, A2 => n16889, ZN => n16891);
   U23 : NAND2_X2 port map( A1 => n16783, A2 => n16886, ZN => n16888);
   U24 : NAND2_X2 port map( A1 => n16781, A2 => n16883, ZN => n16885);
   U25 : NAND2_X2 port map( A1 => n16783, A2 => n16870, ZN => n16882);
   U26 : NAND2_X2 port map( A1 => n16780, A2 => n16846, ZN => n16848);
   U27 : NAND2_X2 port map( A1 => n16780, A2 => n16843, ZN => n16845);
   U28 : NAND2_X2 port map( A1 => n16781, A2 => n16813, ZN => n16815);
   U29 : NAND2_X2 port map( A1 => n16780, A2 => n16807, ZN => n16809);
   U30 : NAND2_X2 port map( A1 => n16782, A2 => n16803, ZN => n16805);
   U31 : NAND2_X2 port map( A1 => n16783, A2 => n16799, ZN => n16801);
   U32 : INV_X1 port map( A => ADD_WR(4), ZN => n16901);
   U33 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n16810);
   U34 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n16806, ZN => n16911);
   U35 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n16842, ZN => n16812);
   U36 : CLKBUF_X1 port map( A => n17749, Z => n17694);
   U37 : CLKBUF_X1 port map( A => n18531, Z => n18476);
   U38 : NAND2_X1 port map( A1 => n16781, A2 => n16924, ZN => n16927);
   U39 : NAND2_X1 port map( A1 => n16782, A2 => n16907, ZN => n16910);
   U40 : CLKBUF_X1 port map( A => n16870, Z => n16880);
   U41 : NAND2_X1 port map( A1 => n16781, A2 => n16834, ZN => n16837);
   U42 : CLKBUF_X1 port map( A => n16876, Z => n16962);
   U43 : CLKBUF_X1 port map( A => n16860, Z => n16946);
   U44 : CLKBUF_X1 port map( A => n16813, Z => n16814);
   U45 : NAND2_X1 port map( A1 => n16782, A2 => n16795, ZN => n16798);
   U46 : CLKBUF_X1 port map( A => n16789, Z => n16790);
   U47 : CLKBUF_X1 port map( A => n16788, Z => n16785);
   U48 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1), 
                           ZN => n16902);
   U49 : INV_X1 port map( A => ADD_WR(3), ZN => n16784);
   U50 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n16784, ZN => n16842)
                           ;
   U51 : NAND2_X1 port map( A1 => n16902, A2 => n16812, ZN => n16786);
   U52 : CLKBUF_X1 port map( A => n16786, Z => n16787);
   U53 : NAND2_X1 port map( A1 => n16782, A2 => n16787, ZN => n16788);
   U54 : NAND2_X1 port map( A1 => n16783, A2 => DATAIN(31), ZN => n16934);
   U55 : CLKBUF_X1 port map( A => n16934, Z => n16896);
   U56 : OAI22_X1 port map( A1 => n18537, A2 => n16785, B1 => n16896, B2 => 
                           n16787, ZN => n2166);
   U57 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(30), ZN => n16849);
   U58 : OAI22_X1 port map( A1 => n19305, A2 => n16788, B1 => n16787, B2 => 
                           n16849, ZN => n2165);
   U59 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(29), ZN => n16850);
   U60 : OAI22_X1 port map( A1 => n18538, A2 => n16785, B1 => n16787, B2 => 
                           n16850, ZN => n2164);
   U61 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(28), ZN => n16851);
   U62 : OAI22_X1 port map( A1 => n18794, A2 => n16788, B1 => n16787, B2 => 
                           n16851, ZN => n2163);
   U63 : NAND2_X1 port map( A1 => n16783, A2 => DATAIN(27), ZN => n16852);
   U64 : OAI22_X1 port map( A1 => n19052, A2 => n16785, B1 => n16787, B2 => 
                           n16852, ZN => n2162);
   U65 : NAND2_X1 port map( A1 => n16783, A2 => DATAIN(26), ZN => n16853);
   U66 : OAI22_X1 port map( A1 => n18539, A2 => n16788, B1 => n16787, B2 => 
                           n16853, ZN => n2161);
   U67 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(25), ZN => n16854);
   U68 : OAI22_X1 port map( A1 => n18795, A2 => n16785, B1 => n16787, B2 => 
                           n16854, ZN => n2160);
   U69 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(24), ZN => n16855);
   U70 : OAI22_X1 port map( A1 => n19053, A2 => n16788, B1 => n16787, B2 => 
                           n16855, ZN => n2159);
   U71 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(23), ZN => n16856);
   U72 : OAI22_X1 port map( A1 => n18540, A2 => n16785, B1 => n16786, B2 => 
                           n16856, ZN => n2158);
   U73 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(22), ZN => n16857);
   U74 : OAI22_X1 port map( A1 => n18796, A2 => n16788, B1 => n16786, B2 => 
                           n16857, ZN => n2157);
   U75 : NAND2_X1 port map( A1 => n16783, A2 => DATAIN(21), ZN => n16858);
   U76 : OAI22_X1 port map( A1 => n18541, A2 => n16788, B1 => n16786, B2 => 
                           n16858, ZN => n2156);
   U77 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(20), ZN => n16859);
   U78 : OAI22_X1 port map( A1 => n18797, A2 => n16788, B1 => n16786, B2 => 
                           n16859, ZN => n2155);
   U79 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(19), ZN => n16860);
   U80 : OAI22_X1 port map( A1 => n18798, A2 => n16785, B1 => n16786, B2 => 
                           n16860, ZN => n2154);
   U81 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(18), ZN => n16861);
   U82 : OAI22_X1 port map( A1 => n18799, A2 => n16785, B1 => n16786, B2 => 
                           n16861, ZN => n2153);
   U83 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(17), ZN => n16862);
   U84 : OAI22_X1 port map( A1 => n18800, A2 => n16785, B1 => n16786, B2 => 
                           n16862, ZN => n2152);
   U85 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(16), ZN => n16863);
   U86 : OAI22_X1 port map( A1 => n19306, A2 => n16785, B1 => n16786, B2 => 
                           n16863, ZN => n2151);
   U87 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(15), ZN => n16864);
   U88 : OAI22_X1 port map( A1 => n18542, A2 => n16785, B1 => n16787, B2 => 
                           n16864, ZN => n2150);
   U89 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(14), ZN => n16865);
   U90 : OAI22_X1 port map( A1 => n18543, A2 => n16785, B1 => n16786, B2 => 
                           n16865, ZN => n2149);
   U91 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(13), ZN => n16866);
   U92 : OAI22_X1 port map( A1 => n18801, A2 => n16785, B1 => n16787, B2 => 
                           n16866, ZN => n2148);
   U93 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(12), ZN => n16867);
   U94 : OAI22_X1 port map( A1 => n18544, A2 => n16785, B1 => n16786, B2 => 
                           n16867, ZN => n2147);
   U95 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(11), ZN => n16868);
   U96 : OAI22_X1 port map( A1 => n19307, A2 => n16785, B1 => n16786, B2 => 
                           n16868, ZN => n2146);
   U97 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(10), ZN => n16869);
   U98 : OAI22_X1 port map( A1 => n18545, A2 => n16785, B1 => n16786, B2 => 
                           n16869, ZN => n2145);
   U99 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(9), ZN => n16871);
   U100 : OAI22_X1 port map( A1 => n18802, A2 => n16785, B1 => n16787, B2 => 
                           n16871, ZN => n2144);
   U101 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(8), ZN => n16872);
   U102 : OAI22_X1 port map( A1 => n18546, A2 => n16785, B1 => n16786, B2 => 
                           n16872, ZN => n2143);
   U103 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(7), ZN => n16873);
   U104 : OAI22_X1 port map( A1 => n18803, A2 => n16788, B1 => n16787, B2 => 
                           n16873, ZN => n2142);
   U105 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(6), ZN => n16874);
   U106 : OAI22_X1 port map( A1 => n18804, A2 => n16788, B1 => n16786, B2 => 
                           n16874, ZN => n2141);
   U107 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(5), ZN => n16875);
   U108 : OAI22_X1 port map( A1 => n18547, A2 => n16788, B1 => n16787, B2 => 
                           n16875, ZN => n2140);
   U109 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(4), ZN => n16876);
   U110 : OAI22_X1 port map( A1 => n19308, A2 => n16788, B1 => n16786, B2 => 
                           n16876, ZN => n2139);
   U111 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(3), ZN => n16877);
   U112 : OAI22_X1 port map( A1 => n18805, A2 => n16788, B1 => n16787, B2 => 
                           n16877, ZN => n2138);
   U113 : NAND2_X1 port map( A1 => n16782, A2 => DATAIN(2), ZN => n16878);
   U114 : OAI22_X1 port map( A1 => n19054, A2 => n16788, B1 => n16786, B2 => 
                           n16878, ZN => n2137);
   U115 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(1), ZN => n16879);
   U116 : OAI22_X1 port map( A1 => n19055, A2 => n16788, B1 => n16787, B2 => 
                           n16879, ZN => n2136);
   U117 : NAND2_X1 port map( A1 => n16781, A2 => DATAIN(0), ZN => n16881);
   U118 : OAI22_X1 port map( A1 => n18548, A2 => n16788, B1 => n16787, B2 => 
                           n16881, ZN => n2135);
   U119 : INV_X1 port map( A => ADD_WR(0), ZN => n16802);
   U120 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n16802, ZN 
                           => n16906);
   U121 : NAND2_X1 port map( A1 => n16812, A2 => n16906, ZN => n16789);
   U122 : NAND2_X2 port map( A1 => n16783, A2 => n16789, ZN => n16791);
   U123 : OAI22_X1 port map( A1 => n19309, A2 => n16791, B1 => n16934, B2 => 
                           n16790, ZN => n2134);
   U124 : OAI22_X1 port map( A1 => n19056, A2 => n16791, B1 => n16849, B2 => 
                           n16789, ZN => n2133);
   U125 : OAI22_X1 port map( A1 => n18806, A2 => n16791, B1 => n16850, B2 => 
                           n16790, ZN => n2132);
   U126 : OAI22_X1 port map( A1 => n19310, A2 => n16791, B1 => n16851, B2 => 
                           n16789, ZN => n2131);
   U127 : OAI22_X1 port map( A1 => n18549, A2 => n16791, B1 => n16852, B2 => 
                           n16790, ZN => n2130);
   U128 : OAI22_X1 port map( A1 => n19057, A2 => n16791, B1 => n16853, B2 => 
                           n16789, ZN => n2129);
   U129 : OAI22_X1 port map( A1 => n18550, A2 => n16791, B1 => n16854, B2 => 
                           n16790, ZN => n2128);
   U130 : OAI22_X1 port map( A1 => n18807, A2 => n16791, B1 => n16855, B2 => 
                           n16789, ZN => n2127);
   U131 : OAI22_X1 port map( A1 => n18808, A2 => n16791, B1 => n16856, B2 => 
                           n16790, ZN => n2126);
   U132 : OAI22_X1 port map( A1 => n18551, A2 => n16791, B1 => n16857, B2 => 
                           n16789, ZN => n2125);
   U133 : OAI22_X1 port map( A1 => n19058, A2 => n16791, B1 => n16858, B2 => 
                           n16789, ZN => n2124);
   U134 : OAI22_X1 port map( A1 => n19311, A2 => n16791, B1 => n16859, B2 => 
                           n16790, ZN => n2123);
   U135 : OAI22_X1 port map( A1 => n19059, A2 => n16791, B1 => n16860, B2 => 
                           n16789, ZN => n2122);
   U136 : OAI22_X1 port map( A1 => n19312, A2 => n16791, B1 => n16861, B2 => 
                           n16790, ZN => n2121);
   U137 : OAI22_X1 port map( A1 => n19060, A2 => n16791, B1 => n16862, B2 => 
                           n16789, ZN => n2120);
   U138 : OAI22_X1 port map( A1 => n18809, A2 => n16791, B1 => n16863, B2 => 
                           n16790, ZN => n2119);
   U139 : OAI22_X1 port map( A1 => n18552, A2 => n16791, B1 => n16864, B2 => 
                           n16789, ZN => n2118);
   U140 : OAI22_X1 port map( A1 => n19061, A2 => n16791, B1 => n16865, B2 => 
                           n16789, ZN => n2117);
   U141 : OAI22_X1 port map( A1 => n19313, A2 => n16791, B1 => n16866, B2 => 
                           n16789, ZN => n2116);
   U142 : OAI22_X1 port map( A1 => n18553, A2 => n16791, B1 => n16867, B2 => 
                           n16789, ZN => n2115);
   U143 : OAI22_X1 port map( A1 => n19062, A2 => n16791, B1 => n16868, B2 => 
                           n16789, ZN => n2114);
   U144 : OAI22_X1 port map( A1 => n18554, A2 => n16791, B1 => n16869, B2 => 
                           n16789, ZN => n2113);
   U145 : OAI22_X1 port map( A1 => n19314, A2 => n16791, B1 => n16871, B2 => 
                           n16789, ZN => n2112);
   U146 : OAI22_X1 port map( A1 => n19315, A2 => n16791, B1 => n16872, B2 => 
                           n16790, ZN => n2111);
   U147 : OAI22_X1 port map( A1 => n19063, A2 => n16791, B1 => n16873, B2 => 
                           n16790, ZN => n2110);
   U148 : OAI22_X1 port map( A1 => n19316, A2 => n16791, B1 => n16874, B2 => 
                           n16790, ZN => n2109);
   U149 : OAI22_X1 port map( A1 => n18810, A2 => n16791, B1 => n16875, B2 => 
                           n16790, ZN => n2108);
   U150 : OAI22_X1 port map( A1 => n18811, A2 => n16791, B1 => n16876, B2 => 
                           n16790, ZN => n2107);
   U151 : OAI22_X1 port map( A1 => n18555, A2 => n16791, B1 => n16877, B2 => 
                           n16790, ZN => n2106);
   U152 : OAI22_X1 port map( A1 => n18812, A2 => n16791, B1 => n16878, B2 => 
                           n16790, ZN => n2105);
   U153 : OAI22_X1 port map( A1 => n19317, A2 => n16791, B1 => n16879, B2 => 
                           n16790, ZN => n2104);
   U154 : OAI22_X1 port map( A1 => n19064, A2 => n16791, B1 => n16881, B2 => 
                           n16790, ZN => n2103);
   U155 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n16802, ZN => n16806);
   U156 : NAND2_X1 port map( A1 => n16812, A2 => n16911, ZN => n16792);
   U157 : NAND2_X2 port map( A1 => n16780, A2 => n16792, ZN => n16794);
   U158 : CLKBUF_X1 port map( A => n16792, Z => n16793);
   U159 : OAI22_X1 port map( A1 => n18813, A2 => n16794, B1 => n16896, B2 => 
                           n16793, ZN => n2102);
   U160 : OAI22_X1 port map( A1 => n18814, A2 => n16794, B1 => n16849, B2 => 
                           n16792, ZN => n2101);
   U161 : OAI22_X1 port map( A1 => n18556, A2 => n16794, B1 => n16850, B2 => 
                           n16793, ZN => n2100);
   U162 : OAI22_X1 port map( A1 => n18557, A2 => n16794, B1 => n16851, B2 => 
                           n16792, ZN => n2099);
   U163 : OAI22_X1 port map( A1 => n18558, A2 => n16794, B1 => n16852, B2 => 
                           n16793, ZN => n2098);
   U164 : OAI22_X1 port map( A1 => n18559, A2 => n16794, B1 => n16853, B2 => 
                           n16792, ZN => n2097);
   U165 : OAI22_X1 port map( A1 => n19318, A2 => n16794, B1 => n16854, B2 => 
                           n16793, ZN => n2096);
   U166 : OAI22_X1 port map( A1 => n18815, A2 => n16794, B1 => n16855, B2 => 
                           n16792, ZN => n2095);
   U167 : OAI22_X1 port map( A1 => n19319, A2 => n16794, B1 => n16856, B2 => 
                           n16793, ZN => n2094);
   U168 : OAI22_X1 port map( A1 => n18560, A2 => n16794, B1 => n16857, B2 => 
                           n16792, ZN => n2093);
   U169 : OAI22_X1 port map( A1 => n18816, A2 => n16794, B1 => n16858, B2 => 
                           n16792, ZN => n2092);
   U170 : OAI22_X1 port map( A1 => n18561, A2 => n16794, B1 => n16859, B2 => 
                           n16793, ZN => n2091);
   U171 : OAI22_X1 port map( A1 => n18817, A2 => n16794, B1 => n16860, B2 => 
                           n16792, ZN => n2090);
   U172 : OAI22_X1 port map( A1 => n18562, A2 => n16794, B1 => n16861, B2 => 
                           n16793, ZN => n2089);
   U173 : OAI22_X1 port map( A1 => n19065, A2 => n16794, B1 => n16862, B2 => 
                           n16792, ZN => n2088);
   U174 : OAI22_X1 port map( A1 => n18563, A2 => n16794, B1 => n16863, B2 => 
                           n16793, ZN => n2087);
   U175 : OAI22_X1 port map( A1 => n19320, A2 => n16794, B1 => n16864, B2 => 
                           n16792, ZN => n2086);
   U176 : OAI22_X1 port map( A1 => n18818, A2 => n16794, B1 => n16865, B2 => 
                           n16792, ZN => n2085);
   U177 : OAI22_X1 port map( A1 => n18819, A2 => n16794, B1 => n16866, B2 => 
                           n16792, ZN => n2084);
   U178 : OAI22_X1 port map( A1 => n18820, A2 => n16794, B1 => n16867, B2 => 
                           n16792, ZN => n2083);
   U179 : OAI22_X1 port map( A1 => n18821, A2 => n16794, B1 => n16868, B2 => 
                           n16792, ZN => n2082);
   U180 : OAI22_X1 port map( A1 => n18564, A2 => n16794, B1 => n16869, B2 => 
                           n16792, ZN => n2081);
   U181 : OAI22_X1 port map( A1 => n18565, A2 => n16794, B1 => n16871, B2 => 
                           n16792, ZN => n2080);
   U182 : OAI22_X1 port map( A1 => n18566, A2 => n16794, B1 => n16872, B2 => 
                           n16793, ZN => n2079);
   U183 : OAI22_X1 port map( A1 => n18822, A2 => n16794, B1 => n16873, B2 => 
                           n16793, ZN => n2078);
   U184 : OAI22_X1 port map( A1 => n18567, A2 => n16794, B1 => n16874, B2 => 
                           n16793, ZN => n2077);
   U185 : OAI22_X1 port map( A1 => n18823, A2 => n16794, B1 => n16875, B2 => 
                           n16793, ZN => n2076);
   U186 : OAI22_X1 port map( A1 => n18824, A2 => n16794, B1 => n16876, B2 => 
                           n16793, ZN => n2075);
   U187 : OAI22_X1 port map( A1 => n18825, A2 => n16794, B1 => n16877, B2 => 
                           n16793, ZN => n2074);
   U188 : OAI22_X1 port map( A1 => n18568, A2 => n16794, B1 => n16878, B2 => 
                           n16793, ZN => n2073);
   U189 : OAI22_X1 port map( A1 => n18569, A2 => n16794, B1 => n16879, B2 => 
                           n16793, ZN => n2072);
   U190 : OAI22_X1 port map( A1 => n18826, A2 => n16794, B1 => n16881, B2 => 
                           n16793, ZN => n2071);
   U191 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n16810, ZN => n16915);
   U192 : NAND2_X1 port map( A1 => n16812, A2 => n16915, ZN => n16795);
   U193 : CLKBUF_X1 port map( A => n16798, Z => n16796);
   U194 : CLKBUF_X1 port map( A => n16795, Z => n16797);
   U195 : OAI22_X1 port map( A1 => n19321, A2 => n16796, B1 => n16934, B2 => 
                           n16797, ZN => n2070);
   U196 : OAI22_X1 port map( A1 => n18570, A2 => n16798, B1 => n16849, B2 => 
                           n16795, ZN => n2069);
   U197 : OAI22_X1 port map( A1 => n19322, A2 => n16796, B1 => n16850, B2 => 
                           n16797, ZN => n2068);
   U198 : OAI22_X1 port map( A1 => n18827, A2 => n16798, B1 => n16851, B2 => 
                           n16795, ZN => n2067);
   U199 : OAI22_X1 port map( A1 => n18828, A2 => n16796, B1 => n16852, B2 => 
                           n16797, ZN => n2066);
   U200 : OAI22_X1 port map( A1 => n19066, A2 => n16798, B1 => n16853, B2 => 
                           n16795, ZN => n2065);
   U201 : OAI22_X1 port map( A1 => n18571, A2 => n16796, B1 => n16854, B2 => 
                           n16797, ZN => n2064);
   U202 : OAI22_X1 port map( A1 => n19323, A2 => n16798, B1 => n16855, B2 => 
                           n16795, ZN => n2063);
   U203 : OAI22_X1 port map( A1 => n18572, A2 => n16796, B1 => n16856, B2 => 
                           n16797, ZN => n2062);
   U204 : OAI22_X1 port map( A1 => n19067, A2 => n16798, B1 => n16857, B2 => 
                           n16795, ZN => n2061);
   U205 : OAI22_X1 port map( A1 => n18573, A2 => n16798, B1 => n16858, B2 => 
                           n16795, ZN => n2060);
   U206 : OAI22_X1 port map( A1 => n19068, A2 => n16798, B1 => n16859, B2 => 
                           n16797, ZN => n2059);
   U207 : OAI22_X1 port map( A1 => n18574, A2 => n16796, B1 => n16860, B2 => 
                           n16795, ZN => n2058);
   U208 : OAI22_X1 port map( A1 => n18575, A2 => n16796, B1 => n16861, B2 => 
                           n16797, ZN => n2057);
   U209 : OAI22_X1 port map( A1 => n18576, A2 => n16796, B1 => n16862, B2 => 
                           n16795, ZN => n2056);
   U210 : OAI22_X1 port map( A1 => n18577, A2 => n16796, B1 => n16863, B2 => 
                           n16797, ZN => n2055);
   U211 : OAI22_X1 port map( A1 => n19069, A2 => n16796, B1 => n16864, B2 => 
                           n16795, ZN => n2054);
   U212 : OAI22_X1 port map( A1 => n19324, A2 => n16796, B1 => n16865, B2 => 
                           n16795, ZN => n2053);
   U213 : OAI22_X1 port map( A1 => n18578, A2 => n16796, B1 => n16866, B2 => 
                           n16795, ZN => n2052);
   U214 : OAI22_X1 port map( A1 => n19325, A2 => n16796, B1 => n16867, B2 => 
                           n16795, ZN => n2051);
   U215 : OAI22_X1 port map( A1 => n18579, A2 => n16796, B1 => n16868, B2 => 
                           n16795, ZN => n2050);
   U216 : OAI22_X1 port map( A1 => n19326, A2 => n16796, B1 => n16869, B2 => 
                           n16795, ZN => n2049);
   U217 : OAI22_X1 port map( A1 => n18829, A2 => n16796, B1 => n16871, B2 => 
                           n16795, ZN => n2048);
   U218 : OAI22_X1 port map( A1 => n18830, A2 => n16796, B1 => n16872, B2 => 
                           n16797, ZN => n2047);
   U219 : OAI22_X1 port map( A1 => n18831, A2 => n16798, B1 => n16873, B2 => 
                           n16797, ZN => n2046);
   U220 : OAI22_X1 port map( A1 => n19070, A2 => n16798, B1 => n16874, B2 => 
                           n16797, ZN => n2045);
   U221 : OAI22_X1 port map( A1 => n19071, A2 => n16798, B1 => n16875, B2 => 
                           n16797, ZN => n2044);
   U222 : OAI22_X1 port map( A1 => n19327, A2 => n16798, B1 => n16876, B2 => 
                           n16797, ZN => n2043);
   U223 : OAI22_X1 port map( A1 => n19072, A2 => n16798, B1 => n16877, B2 => 
                           n16797, ZN => n2042);
   U224 : OAI22_X1 port map( A1 => n18580, A2 => n16798, B1 => n16878, B2 => 
                           n16797, ZN => n2041);
   U225 : OAI22_X1 port map( A1 => n18581, A2 => n16798, B1 => n16879, B2 => 
                           n16797, ZN => n2040);
   U226 : OAI22_X1 port map( A1 => n18582, A2 => n16798, B1 => n16881, B2 => 
                           n16797, ZN => n2039);
   U227 : INV_X1 port map( A => ADD_WR(2), ZN => n16811);
   U228 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n16811, ZN 
                           => n16919);
   U229 : NAND2_X1 port map( A1 => n16812, A2 => n16919, ZN => n16799);
   U230 : CLKBUF_X1 port map( A => n16799, Z => n16800);
   U231 : OAI22_X1 port map( A1 => n19073, A2 => n16801, B1 => n16896, B2 => 
                           n16800, ZN => n2038);
   U232 : OAI22_X1 port map( A1 => n19328, A2 => n16801, B1 => n16849, B2 => 
                           n16799, ZN => n2037);
   U233 : OAI22_X1 port map( A1 => n19329, A2 => n16801, B1 => n16850, B2 => 
                           n16800, ZN => n2036);
   U234 : OAI22_X1 port map( A1 => n19074, A2 => n16801, B1 => n16851, B2 => 
                           n16799, ZN => n2035);
   U235 : OAI22_X1 port map( A1 => n19330, A2 => n16801, B1 => n16852, B2 => 
                           n16800, ZN => n2034);
   U236 : OAI22_X1 port map( A1 => n18832, A2 => n16801, B1 => n16853, B2 => 
                           n16799, ZN => n2033);
   U237 : OAI22_X1 port map( A1 => n19075, A2 => n16801, B1 => n16854, B2 => 
                           n16800, ZN => n2032);
   U238 : OAI22_X1 port map( A1 => n19331, A2 => n16801, B1 => n16855, B2 => 
                           n16799, ZN => n2031);
   U239 : OAI22_X1 port map( A1 => n19076, A2 => n16801, B1 => n16856, B2 => 
                           n16800, ZN => n2030);
   U240 : OAI22_X1 port map( A1 => n19332, A2 => n16801, B1 => n16857, B2 => 
                           n16799, ZN => n2029);
   U241 : OAI22_X1 port map( A1 => n19077, A2 => n16801, B1 => n16858, B2 => 
                           n16799, ZN => n2028);
   U242 : OAI22_X1 port map( A1 => n19078, A2 => n16801, B1 => n16859, B2 => 
                           n16800, ZN => n2027);
   U243 : OAI22_X1 port map( A1 => n19333, A2 => n16801, B1 => n16860, B2 => 
                           n16799, ZN => n2026);
   U244 : OAI22_X1 port map( A1 => n19079, A2 => n16801, B1 => n16861, B2 => 
                           n16800, ZN => n2025);
   U245 : OAI22_X1 port map( A1 => n18833, A2 => n16801, B1 => n16862, B2 => 
                           n16799, ZN => n2024);
   U246 : OAI22_X1 port map( A1 => n19080, A2 => n16801, B1 => n16863, B2 => 
                           n16800, ZN => n2023);
   U247 : OAI22_X1 port map( A1 => n19334, A2 => n16801, B1 => n16864, B2 => 
                           n16799, ZN => n2022);
   U248 : OAI22_X1 port map( A1 => n19081, A2 => n16801, B1 => n16865, B2 => 
                           n16799, ZN => n2021);
   U249 : OAI22_X1 port map( A1 => n19082, A2 => n16801, B1 => n16866, B2 => 
                           n16799, ZN => n2020);
   U250 : OAI22_X1 port map( A1 => n19335, A2 => n16801, B1 => n16867, B2 => 
                           n16799, ZN => n2019);
   U251 : OAI22_X1 port map( A1 => n19083, A2 => n16801, B1 => n16868, B2 => 
                           n16799, ZN => n2018);
   U252 : OAI22_X1 port map( A1 => n19336, A2 => n16801, B1 => n16869, B2 => 
                           n16799, ZN => n2017);
   U253 : OAI22_X1 port map( A1 => n19084, A2 => n16801, B1 => n16871, B2 => 
                           n16799, ZN => n2016);
   U254 : OAI22_X1 port map( A1 => n19337, A2 => n16801, B1 => n16872, B2 => 
                           n16800, ZN => n2015);
   U255 : OAI22_X1 port map( A1 => n19338, A2 => n16801, B1 => n16873, B2 => 
                           n16800, ZN => n2014);
   U256 : OAI22_X1 port map( A1 => n19085, A2 => n16801, B1 => n16874, B2 => 
                           n16800, ZN => n2013);
   U257 : OAI22_X1 port map( A1 => n19086, A2 => n16801, B1 => n16875, B2 => 
                           n16800, ZN => n2012);
   U258 : OAI22_X1 port map( A1 => n18583, A2 => n16801, B1 => n16876, B2 => 
                           n16800, ZN => n2011);
   U259 : OAI22_X1 port map( A1 => n19087, A2 => n16801, B1 => n16877, B2 => 
                           n16800, ZN => n2010);
   U260 : OAI22_X1 port map( A1 => n19088, A2 => n16801, B1 => n16878, B2 => 
                           n16800, ZN => n2009);
   U261 : OAI22_X1 port map( A1 => n18834, A2 => n16801, B1 => n16879, B2 => 
                           n16800, ZN => n2008);
   U262 : OAI22_X1 port map( A1 => n19339, A2 => n16801, B1 => n16881, B2 => 
                           n16800, ZN => n2007);
   U263 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n16802, A3 => n16811, ZN => 
                           n16923);
   U264 : NAND2_X1 port map( A1 => n16812, A2 => n16923, ZN => n16803);
   U265 : CLKBUF_X1 port map( A => n16803, Z => n16804);
   U266 : OAI22_X1 port map( A1 => n18835, A2 => n16805, B1 => n16934, B2 => 
                           n16804, ZN => n2006);
   U267 : OAI22_X1 port map( A1 => n18584, A2 => n16805, B1 => n16849, B2 => 
                           n16803, ZN => n2005);
   U268 : OAI22_X1 port map( A1 => n19340, A2 => n16805, B1 => n16850, B2 => 
                           n16804, ZN => n2004);
   U269 : OAI22_X1 port map( A1 => n19341, A2 => n16805, B1 => n16851, B2 => 
                           n16803, ZN => n2003);
   U270 : OAI22_X1 port map( A1 => n19342, A2 => n16805, B1 => n16852, B2 => 
                           n16804, ZN => n2002);
   U271 : OAI22_X1 port map( A1 => n19343, A2 => n16805, B1 => n16853, B2 => 
                           n16803, ZN => n2001);
   U272 : OAI22_X1 port map( A1 => n19089, A2 => n16805, B1 => n16854, B2 => 
                           n16804, ZN => n2000);
   U273 : OAI22_X1 port map( A1 => n18585, A2 => n16805, B1 => n16855, B2 => 
                           n16803, ZN => n1999);
   U274 : OAI22_X1 port map( A1 => n19344, A2 => n16805, B1 => n16856, B2 => 
                           n16804, ZN => n1998);
   U275 : OAI22_X1 port map( A1 => n19090, A2 => n16805, B1 => n16857, B2 => 
                           n16803, ZN => n1997);
   U276 : OAI22_X1 port map( A1 => n19345, A2 => n16805, B1 => n16858, B2 => 
                           n16803, ZN => n1996);
   U277 : OAI22_X1 port map( A1 => n18836, A2 => n16805, B1 => n16859, B2 => 
                           n16804, ZN => n1995);
   U278 : OAI22_X1 port map( A1 => n19346, A2 => n16805, B1 => n16860, B2 => 
                           n16803, ZN => n1994);
   U279 : OAI22_X1 port map( A1 => n19091, A2 => n16805, B1 => n16861, B2 => 
                           n16804, ZN => n1993);
   U280 : OAI22_X1 port map( A1 => n19347, A2 => n16805, B1 => n16862, B2 => 
                           n16803, ZN => n1992);
   U281 : OAI22_X1 port map( A1 => n19348, A2 => n16805, B1 => n16863, B2 => 
                           n16804, ZN => n1991);
   U282 : OAI22_X1 port map( A1 => n18837, A2 => n16805, B1 => n16864, B2 => 
                           n16803, ZN => n1990);
   U283 : OAI22_X1 port map( A1 => n18586, A2 => n16805, B1 => n16865, B2 => 
                           n16803, ZN => n1989);
   U284 : OAI22_X1 port map( A1 => n19092, A2 => n16805, B1 => n16866, B2 => 
                           n16803, ZN => n1988);
   U285 : OAI22_X1 port map( A1 => n19093, A2 => n16805, B1 => n16867, B2 => 
                           n16803, ZN => n1987);
   U286 : OAI22_X1 port map( A1 => n18838, A2 => n16805, B1 => n16868, B2 => 
                           n16803, ZN => n1986);
   U287 : OAI22_X1 port map( A1 => n19349, A2 => n16805, B1 => n16869, B2 => 
                           n16803, ZN => n1985);
   U288 : OAI22_X1 port map( A1 => n19094, A2 => n16805, B1 => n16871, B2 => 
                           n16803, ZN => n1984);
   U289 : OAI22_X1 port map( A1 => n19095, A2 => n16805, B1 => n16872, B2 => 
                           n16804, ZN => n1983);
   U290 : OAI22_X1 port map( A1 => n19096, A2 => n16805, B1 => n16873, B2 => 
                           n16804, ZN => n1982);
   U291 : OAI22_X1 port map( A1 => n18587, A2 => n16805, B1 => n16874, B2 => 
                           n16804, ZN => n1981);
   U292 : OAI22_X1 port map( A1 => n19350, A2 => n16805, B1 => n16875, B2 => 
                           n16804, ZN => n1980);
   U293 : OAI22_X1 port map( A1 => n19097, A2 => n16805, B1 => n16876, B2 => 
                           n16804, ZN => n1979);
   U294 : OAI22_X1 port map( A1 => n19098, A2 => n16805, B1 => n16877, B2 => 
                           n16804, ZN => n1978);
   U295 : OAI22_X1 port map( A1 => n19351, A2 => n16805, B1 => n16878, B2 => 
                           n16804, ZN => n1977);
   U296 : OAI22_X1 port map( A1 => n19099, A2 => n16805, B1 => n16879, B2 => 
                           n16804, ZN => n1976);
   U297 : OAI22_X1 port map( A1 => n19352, A2 => n16805, B1 => n16881, B2 => 
                           n16804, ZN => n1975);
   U298 : NOR2_X1 port map( A1 => n16811, A2 => n16806, ZN => n16928);
   U299 : NAND2_X1 port map( A1 => n16812, A2 => n16928, ZN => n16807);
   U300 : CLKBUF_X1 port map( A => n16807, Z => n16808);
   U301 : OAI22_X1 port map( A1 => n19100, A2 => n16809, B1 => n16896, B2 => 
                           n16808, ZN => n1974);
   U302 : OAI22_X1 port map( A1 => n19101, A2 => n16809, B1 => n16849, B2 => 
                           n16807, ZN => n1973);
   U303 : OAI22_X1 port map( A1 => n19102, A2 => n16809, B1 => n16850, B2 => 
                           n16808, ZN => n1972);
   U304 : OAI22_X1 port map( A1 => n19103, A2 => n16809, B1 => n16851, B2 => 
                           n16807, ZN => n1971);
   U305 : OAI22_X1 port map( A1 => n19104, A2 => n16809, B1 => n16852, B2 => 
                           n16808, ZN => n1970);
   U306 : OAI22_X1 port map( A1 => n19353, A2 => n16809, B1 => n16853, B2 => 
                           n16807, ZN => n1969);
   U307 : OAI22_X1 port map( A1 => n19354, A2 => n16809, B1 => n16854, B2 => 
                           n16808, ZN => n1968);
   U308 : OAI22_X1 port map( A1 => n19105, A2 => n16809, B1 => n16855, B2 => 
                           n16807, ZN => n1967);
   U309 : OAI22_X1 port map( A1 => n19106, A2 => n16809, B1 => n16856, B2 => 
                           n16808, ZN => n1966);
   U310 : OAI22_X1 port map( A1 => n19355, A2 => n16809, B1 => n16857, B2 => 
                           n16807, ZN => n1965);
   U311 : OAI22_X1 port map( A1 => n19356, A2 => n16809, B1 => n16858, B2 => 
                           n16807, ZN => n1964);
   U312 : OAI22_X1 port map( A1 => n19357, A2 => n16809, B1 => n16859, B2 => 
                           n16808, ZN => n1963);
   U313 : OAI22_X1 port map( A1 => n19107, A2 => n16809, B1 => n16860, B2 => 
                           n16807, ZN => n1962);
   U314 : OAI22_X1 port map( A1 => n19358, A2 => n16809, B1 => n16861, B2 => 
                           n16808, ZN => n1961);
   U315 : OAI22_X1 port map( A1 => n19359, A2 => n16809, B1 => n16862, B2 => 
                           n16807, ZN => n1960);
   U316 : OAI22_X1 port map( A1 => n19360, A2 => n16809, B1 => n16863, B2 => 
                           n16808, ZN => n1959);
   U317 : OAI22_X1 port map( A1 => n19361, A2 => n16809, B1 => n16864, B2 => 
                           n16807, ZN => n1958);
   U318 : OAI22_X1 port map( A1 => n19362, A2 => n16809, B1 => n16865, B2 => 
                           n16807, ZN => n1957);
   U319 : OAI22_X1 port map( A1 => n19108, A2 => n16809, B1 => n16866, B2 => 
                           n16807, ZN => n1956);
   U320 : OAI22_X1 port map( A1 => n19109, A2 => n16809, B1 => n16867, B2 => 
                           n16807, ZN => n1955);
   U321 : OAI22_X1 port map( A1 => n19363, A2 => n16809, B1 => n16868, B2 => 
                           n16807, ZN => n1954);
   U322 : OAI22_X1 port map( A1 => n19110, A2 => n16809, B1 => n16869, B2 => 
                           n16807, ZN => n1953);
   U323 : OAI22_X1 port map( A1 => n19111, A2 => n16809, B1 => n16871, B2 => 
                           n16807, ZN => n1952);
   U324 : OAI22_X1 port map( A1 => n19112, A2 => n16809, B1 => n16872, B2 => 
                           n16808, ZN => n1951);
   U325 : OAI22_X1 port map( A1 => n19113, A2 => n16809, B1 => n16873, B2 => 
                           n16808, ZN => n1950);
   U326 : OAI22_X1 port map( A1 => n19364, A2 => n16809, B1 => n16874, B2 => 
                           n16808, ZN => n1949);
   U327 : OAI22_X1 port map( A1 => n19365, A2 => n16809, B1 => n16875, B2 => 
                           n16808, ZN => n1948);
   U328 : OAI22_X1 port map( A1 => n19114, A2 => n16809, B1 => n16876, B2 => 
                           n16808, ZN => n1947);
   U329 : OAI22_X1 port map( A1 => n19366, A2 => n16809, B1 => n16877, B2 => 
                           n16808, ZN => n1946);
   U330 : OAI22_X1 port map( A1 => n19367, A2 => n16809, B1 => n16878, B2 => 
                           n16808, ZN => n1945);
   U331 : OAI22_X1 port map( A1 => n19368, A2 => n16809, B1 => n16879, B2 => 
                           n16808, ZN => n1944);
   U332 : OAI22_X1 port map( A1 => n19115, A2 => n16809, B1 => n16881, B2 => 
                           n16808, ZN => n1943);
   U333 : NOR2_X1 port map( A1 => n16811, A2 => n16810, ZN => n16933);
   U334 : NAND2_X1 port map( A1 => n16812, A2 => n16933, ZN => n16813);
   U335 : OAI22_X1 port map( A1 => n18588, A2 => n16815, B1 => n16934, B2 => 
                           n16814, ZN => n1942);
   U336 : OAI22_X1 port map( A1 => n18839, A2 => n16815, B1 => n16849, B2 => 
                           n16813, ZN => n1941);
   U337 : OAI22_X1 port map( A1 => n18589, A2 => n16815, B1 => n16850, B2 => 
                           n16814, ZN => n1940);
   U338 : OAI22_X1 port map( A1 => n18590, A2 => n16815, B1 => n16851, B2 => 
                           n16813, ZN => n1939);
   U339 : OAI22_X1 port map( A1 => n18840, A2 => n16815, B1 => n16852, B2 => 
                           n16814, ZN => n1938);
   U340 : OAI22_X1 port map( A1 => n18841, A2 => n16815, B1 => n16853, B2 => 
                           n16813, ZN => n1937);
   U341 : OAI22_X1 port map( A1 => n18842, A2 => n16815, B1 => n16854, B2 => 
                           n16814, ZN => n1936);
   U342 : OAI22_X1 port map( A1 => n18591, A2 => n16815, B1 => n16855, B2 => 
                           n16813, ZN => n1935);
   U343 : OAI22_X1 port map( A1 => n18843, A2 => n16815, B1 => n16856, B2 => 
                           n16814, ZN => n1934);
   U344 : OAI22_X1 port map( A1 => n18844, A2 => n16815, B1 => n16857, B2 => 
                           n16813, ZN => n1933);
   U345 : OAI22_X1 port map( A1 => n18845, A2 => n16815, B1 => n16858, B2 => 
                           n16813, ZN => n1932);
   U346 : OAI22_X1 port map( A1 => n18592, A2 => n16815, B1 => n16859, B2 => 
                           n16814, ZN => n1931);
   U347 : OAI22_X1 port map( A1 => n18593, A2 => n16815, B1 => n16860, B2 => 
                           n16813, ZN => n1930);
   U348 : OAI22_X1 port map( A1 => n18846, A2 => n16815, B1 => n16861, B2 => 
                           n16814, ZN => n1929);
   U349 : OAI22_X1 port map( A1 => n18594, A2 => n16815, B1 => n16862, B2 => 
                           n16813, ZN => n1928);
   U350 : OAI22_X1 port map( A1 => n18595, A2 => n16815, B1 => n16863, B2 => 
                           n16814, ZN => n1927);
   U351 : OAI22_X1 port map( A1 => n18596, A2 => n16815, B1 => n16864, B2 => 
                           n16813, ZN => n1926);
   U352 : OAI22_X1 port map( A1 => n18847, A2 => n16815, B1 => n16865, B2 => 
                           n16813, ZN => n1925);
   U353 : OAI22_X1 port map( A1 => n18848, A2 => n16815, B1 => n16866, B2 => 
                           n16813, ZN => n1924);
   U354 : OAI22_X1 port map( A1 => n18849, A2 => n16815, B1 => n16867, B2 => 
                           n16813, ZN => n1923);
   U355 : OAI22_X1 port map( A1 => n18597, A2 => n16815, B1 => n16868, B2 => 
                           n16813, ZN => n1922);
   U356 : OAI22_X1 port map( A1 => n18850, A2 => n16815, B1 => n16869, B2 => 
                           n16813, ZN => n1921);
   U357 : OAI22_X1 port map( A1 => n18851, A2 => n16815, B1 => n16871, B2 => 
                           n16813, ZN => n1920);
   U358 : OAI22_X1 port map( A1 => n18852, A2 => n16815, B1 => n16872, B2 => 
                           n16814, ZN => n1919);
   U359 : OAI22_X1 port map( A1 => n18598, A2 => n16815, B1 => n16873, B2 => 
                           n16814, ZN => n1918);
   U360 : OAI22_X1 port map( A1 => n18853, A2 => n16815, B1 => n16874, B2 => 
                           n16814, ZN => n1917);
   U361 : OAI22_X1 port map( A1 => n18599, A2 => n16815, B1 => n16875, B2 => 
                           n16814, ZN => n1916);
   U362 : OAI22_X1 port map( A1 => n18600, A2 => n16815, B1 => n16876, B2 => 
                           n16814, ZN => n1915);
   U363 : OAI22_X1 port map( A1 => n18854, A2 => n16815, B1 => n16877, B2 => 
                           n16814, ZN => n1914);
   U364 : OAI22_X1 port map( A1 => n18855, A2 => n16815, B1 => n16878, B2 => 
                           n16814, ZN => n1913);
   U365 : OAI22_X1 port map( A1 => n18856, A2 => n16815, B1 => n16879, B2 => 
                           n16814, ZN => n1912);
   U366 : OAI22_X1 port map( A1 => n18857, A2 => n16815, B1 => n16881, B2 => 
                           n16814, ZN => n1911);
   U367 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => ADD_WR(3), ZN => 
                           n16900);
   U368 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n16900, ZN => n16838);
   U369 : NAND2_X1 port map( A1 => n16902, A2 => n16838, ZN => n16816);
   U370 : CLKBUF_X1 port map( A => n16816, Z => n16817);
   U371 : OAI22_X1 port map( A1 => n18858, A2 => n16818, B1 => n16896, B2 => 
                           n16817, ZN => n1910);
   U372 : OAI22_X1 port map( A1 => n19116, A2 => n16818, B1 => n16849, B2 => 
                           n16816, ZN => n1909);
   U373 : OAI22_X1 port map( A1 => n18601, A2 => n16818, B1 => n16850, B2 => 
                           n16817, ZN => n1908);
   U374 : OAI22_X1 port map( A1 => n18602, A2 => n16818, B1 => n16851, B2 => 
                           n16816, ZN => n1907);
   U375 : OAI22_X1 port map( A1 => n19117, A2 => n16818, B1 => n16852, B2 => 
                           n16817, ZN => n1906);
   U376 : OAI22_X1 port map( A1 => n18859, A2 => n16818, B1 => n16853, B2 => 
                           n16816, ZN => n1905);
   U377 : OAI22_X1 port map( A1 => n18603, A2 => n16818, B1 => n16854, B2 => 
                           n16817, ZN => n1904);
   U378 : OAI22_X1 port map( A1 => n18604, A2 => n16818, B1 => n16855, B2 => 
                           n16816, ZN => n1903);
   U379 : OAI22_X1 port map( A1 => n18605, A2 => n16818, B1 => n16856, B2 => 
                           n16817, ZN => n1902);
   U380 : OAI22_X1 port map( A1 => n18606, A2 => n16818, B1 => n16857, B2 => 
                           n16816, ZN => n1901);
   U381 : OAI22_X1 port map( A1 => n18860, A2 => n16818, B1 => n16858, B2 => 
                           n16816, ZN => n1900);
   U382 : OAI22_X1 port map( A1 => n19369, A2 => n16818, B1 => n16859, B2 => 
                           n16817, ZN => n1899);
   U383 : OAI22_X1 port map( A1 => n18607, A2 => n16818, B1 => n16860, B2 => 
                           n16816, ZN => n1898);
   U384 : OAI22_X1 port map( A1 => n18608, A2 => n16818, B1 => n16861, B2 => 
                           n16817, ZN => n1897);
   U385 : OAI22_X1 port map( A1 => n19118, A2 => n16818, B1 => n16862, B2 => 
                           n16816, ZN => n1896);
   U386 : OAI22_X1 port map( A1 => n18609, A2 => n16818, B1 => n16863, B2 => 
                           n16817, ZN => n1895);
   U387 : OAI22_X1 port map( A1 => n19119, A2 => n16818, B1 => n16864, B2 => 
                           n16816, ZN => n1894);
   U388 : OAI22_X1 port map( A1 => n18610, A2 => n16818, B1 => n16865, B2 => 
                           n16816, ZN => n1893);
   U389 : OAI22_X1 port map( A1 => n19120, A2 => n16818, B1 => n16866, B2 => 
                           n16816, ZN => n1892);
   U390 : OAI22_X1 port map( A1 => n19121, A2 => n16818, B1 => n16867, B2 => 
                           n16816, ZN => n1891);
   U391 : OAI22_X1 port map( A1 => n18611, A2 => n16818, B1 => n16868, B2 => 
                           n16816, ZN => n1890);
   U392 : OAI22_X1 port map( A1 => n18861, A2 => n16818, B1 => n16869, B2 => 
                           n16816, ZN => n1889);
   U393 : OAI22_X1 port map( A1 => n18612, A2 => n16818, B1 => n16871, B2 => 
                           n16816, ZN => n1888);
   U394 : OAI22_X1 port map( A1 => n19122, A2 => n16818, B1 => n16872, B2 => 
                           n16817, ZN => n1887);
   U395 : OAI22_X1 port map( A1 => n19370, A2 => n16818, B1 => n16873, B2 => 
                           n16817, ZN => n1886);
   U396 : OAI22_X1 port map( A1 => n18613, A2 => n16818, B1 => n16874, B2 => 
                           n16817, ZN => n1885);
   U397 : OAI22_X1 port map( A1 => n19371, A2 => n16818, B1 => n16875, B2 => 
                           n16817, ZN => n1884);
   U398 : OAI22_X1 port map( A1 => n18614, A2 => n16818, B1 => n16876, B2 => 
                           n16817, ZN => n1883);
   U399 : OAI22_X1 port map( A1 => n19123, A2 => n16818, B1 => n16877, B2 => 
                           n16817, ZN => n1882);
   U400 : OAI22_X1 port map( A1 => n18615, A2 => n16818, B1 => n16878, B2 => 
                           n16817, ZN => n1881);
   U401 : OAI22_X1 port map( A1 => n18616, A2 => n16818, B1 => n16879, B2 => 
                           n16817, ZN => n1880);
   U402 : OAI22_X1 port map( A1 => n18617, A2 => n16818, B1 => n16881, B2 => 
                           n16817, ZN => n1879);
   U403 : NAND2_X1 port map( A1 => n16906, A2 => n16838, ZN => n16819);
   U404 : CLKBUF_X1 port map( A => n16819, Z => n16820);
   U405 : OAI22_X1 port map( A1 => n19372, A2 => n16821, B1 => n16934, B2 => 
                           n16820, ZN => n1878);
   U406 : OAI22_X1 port map( A1 => n19373, A2 => n16821, B1 => n16849, B2 => 
                           n16819, ZN => n1877);
   U407 : OAI22_X1 port map( A1 => n19374, A2 => n16821, B1 => n16850, B2 => 
                           n16820, ZN => n1876);
   U408 : OAI22_X1 port map( A1 => n18862, A2 => n16821, B1 => n16851, B2 => 
                           n16819, ZN => n1875);
   U409 : OAI22_X1 port map( A1 => n19124, A2 => n16821, B1 => n16852, B2 => 
                           n16820, ZN => n1874);
   U410 : OAI22_X1 port map( A1 => n19125, A2 => n16821, B1 => n16853, B2 => 
                           n16819, ZN => n1873);
   U411 : OAI22_X1 port map( A1 => n19126, A2 => n16821, B1 => n16854, B2 => 
                           n16820, ZN => n1872);
   U412 : OAI22_X1 port map( A1 => n19375, A2 => n16821, B1 => n16855, B2 => 
                           n16819, ZN => n1871);
   U413 : OAI22_X1 port map( A1 => n19127, A2 => n16821, B1 => n16856, B2 => 
                           n16820, ZN => n1870);
   U414 : OAI22_X1 port map( A1 => n19376, A2 => n16821, B1 => n16857, B2 => 
                           n16819, ZN => n1869);
   U415 : OAI22_X1 port map( A1 => n18618, A2 => n16821, B1 => n16858, B2 => 
                           n16819, ZN => n1868);
   U416 : OAI22_X1 port map( A1 => n18863, A2 => n16821, B1 => n16859, B2 => 
                           n16820, ZN => n1867);
   U417 : OAI22_X1 port map( A1 => n18619, A2 => n16821, B1 => n16860, B2 => 
                           n16819, ZN => n1866);
   U418 : OAI22_X1 port map( A1 => n18864, A2 => n16821, B1 => n16861, B2 => 
                           n16820, ZN => n1865);
   U419 : OAI22_X1 port map( A1 => n19377, A2 => n16821, B1 => n16862, B2 => 
                           n16819, ZN => n1864);
   U420 : OAI22_X1 port map( A1 => n19128, A2 => n16821, B1 => n16863, B2 => 
                           n16820, ZN => n1863);
   U421 : OAI22_X1 port map( A1 => n19378, A2 => n16821, B1 => n16864, B2 => 
                           n16819, ZN => n1862);
   U422 : OAI22_X1 port map( A1 => n19379, A2 => n16821, B1 => n16865, B2 => 
                           n16819, ZN => n1861);
   U423 : OAI22_X1 port map( A1 => n18865, A2 => n16821, B1 => n16866, B2 => 
                           n16819, ZN => n1860);
   U424 : OAI22_X1 port map( A1 => n19129, A2 => n16821, B1 => n16867, B2 => 
                           n16819, ZN => n1859);
   U425 : OAI22_X1 port map( A1 => n19130, A2 => n16821, B1 => n16868, B2 => 
                           n16819, ZN => n1858);
   U426 : OAI22_X1 port map( A1 => n18620, A2 => n16821, B1 => n16869, B2 => 
                           n16819, ZN => n1857);
   U427 : OAI22_X1 port map( A1 => n19380, A2 => n16821, B1 => n16871, B2 => 
                           n16819, ZN => n1856);
   U428 : OAI22_X1 port map( A1 => n18621, A2 => n16821, B1 => n16872, B2 => 
                           n16820, ZN => n1855);
   U429 : OAI22_X1 port map( A1 => n19131, A2 => n16821, B1 => n16873, B2 => 
                           n16820, ZN => n1854);
   U430 : OAI22_X1 port map( A1 => n18866, A2 => n16821, B1 => n16874, B2 => 
                           n16820, ZN => n1853);
   U431 : OAI22_X1 port map( A1 => n18867, A2 => n16821, B1 => n16875, B2 => 
                           n16820, ZN => n1852);
   U432 : OAI22_X1 port map( A1 => n19381, A2 => n16821, B1 => n16876, B2 => 
                           n16820, ZN => n1851);
   U433 : OAI22_X1 port map( A1 => n19382, A2 => n16821, B1 => n16877, B2 => 
                           n16820, ZN => n1850);
   U434 : OAI22_X1 port map( A1 => n19383, A2 => n16821, B1 => n16878, B2 => 
                           n16820, ZN => n1849);
   U435 : OAI22_X1 port map( A1 => n18622, A2 => n16821, B1 => n16879, B2 => 
                           n16820, ZN => n1848);
   U436 : OAI22_X1 port map( A1 => n18623, A2 => n16821, B1 => n16881, B2 => 
                           n16820, ZN => n1847);
   U437 : NAND2_X1 port map( A1 => n16911, A2 => n16838, ZN => n16822);
   U438 : CLKBUF_X1 port map( A => n16822, Z => n16823);
   U439 : OAI22_X1 port map( A1 => n19132, A2 => n16824, B1 => n16934, B2 => 
                           n16823, ZN => n1846);
   U440 : OAI22_X1 port map( A1 => n18624, A2 => n16824, B1 => n16849, B2 => 
                           n16822, ZN => n1845);
   U441 : OAI22_X1 port map( A1 => n18625, A2 => n16824, B1 => n16850, B2 => 
                           n16823, ZN => n1844);
   U442 : OAI22_X1 port map( A1 => n18868, A2 => n16824, B1 => n16851, B2 => 
                           n16822, ZN => n1843);
   U443 : OAI22_X1 port map( A1 => n18626, A2 => n16824, B1 => n16852, B2 => 
                           n16823, ZN => n1842);
   U444 : OAI22_X1 port map( A1 => n18869, A2 => n16824, B1 => n16853, B2 => 
                           n16822, ZN => n1841);
   U445 : OAI22_X1 port map( A1 => n18870, A2 => n16824, B1 => n16854, B2 => 
                           n16823, ZN => n1840);
   U446 : OAI22_X1 port map( A1 => n18627, A2 => n16824, B1 => n16855, B2 => 
                           n16822, ZN => n1839);
   U447 : OAI22_X1 port map( A1 => n18871, A2 => n16824, B1 => n16856, B2 => 
                           n16823, ZN => n1838);
   U448 : OAI22_X1 port map( A1 => n18628, A2 => n16824, B1 => n16857, B2 => 
                           n16822, ZN => n1837);
   U449 : OAI22_X1 port map( A1 => n18629, A2 => n16824, B1 => n16858, B2 => 
                           n16822, ZN => n1836);
   U450 : OAI22_X1 port map( A1 => n18872, A2 => n16824, B1 => n16859, B2 => 
                           n16823, ZN => n1835);
   U451 : OAI22_X1 port map( A1 => n19133, A2 => n16824, B1 => n16860, B2 => 
                           n16822, ZN => n1834);
   U452 : OAI22_X1 port map( A1 => n18873, A2 => n16824, B1 => n16861, B2 => 
                           n16823, ZN => n1833);
   U453 : OAI22_X1 port map( A1 => n18630, A2 => n16824, B1 => n16862, B2 => 
                           n16822, ZN => n1832);
   U454 : OAI22_X1 port map( A1 => n18874, A2 => n16824, B1 => n16863, B2 => 
                           n16823, ZN => n1831);
   U455 : OAI22_X1 port map( A1 => n18631, A2 => n16824, B1 => n16864, B2 => 
                           n16822, ZN => n1830);
   U456 : OAI22_X1 port map( A1 => n18632, A2 => n16824, B1 => n16865, B2 => 
                           n16822, ZN => n1829);
   U457 : OAI22_X1 port map( A1 => n18875, A2 => n16824, B1 => n16866, B2 => 
                           n16822, ZN => n1828);
   U458 : OAI22_X1 port map( A1 => n18876, A2 => n16824, B1 => n16867, B2 => 
                           n16822, ZN => n1827);
   U459 : OAI22_X1 port map( A1 => n18633, A2 => n16824, B1 => n16868, B2 => 
                           n16822, ZN => n1826);
   U460 : OAI22_X1 port map( A1 => n18634, A2 => n16824, B1 => n16869, B2 => 
                           n16822, ZN => n1825);
   U461 : OAI22_X1 port map( A1 => n18635, A2 => n16824, B1 => n16871, B2 => 
                           n16822, ZN => n1824);
   U462 : OAI22_X1 port map( A1 => n18636, A2 => n16824, B1 => n16872, B2 => 
                           n16823, ZN => n1823);
   U463 : OAI22_X1 port map( A1 => n18877, A2 => n16824, B1 => n16873, B2 => 
                           n16823, ZN => n1822);
   U464 : OAI22_X1 port map( A1 => n18878, A2 => n16824, B1 => n16874, B2 => 
                           n16823, ZN => n1821);
   U465 : OAI22_X1 port map( A1 => n18637, A2 => n16824, B1 => n16875, B2 => 
                           n16823, ZN => n1820);
   U466 : OAI22_X1 port map( A1 => n18638, A2 => n16824, B1 => n16876, B2 => 
                           n16823, ZN => n1819);
   U467 : OAI22_X1 port map( A1 => n18639, A2 => n16824, B1 => n16877, B2 => 
                           n16823, ZN => n1818);
   U468 : OAI22_X1 port map( A1 => n18879, A2 => n16824, B1 => n16878, B2 => 
                           n16823, ZN => n1817);
   U469 : OAI22_X1 port map( A1 => n18880, A2 => n16824, B1 => n16879, B2 => 
                           n16823, ZN => n1816);
   U470 : OAI22_X1 port map( A1 => n18881, A2 => n16824, B1 => n16881, B2 => 
                           n16823, ZN => n1815);
   U471 : NAND2_X1 port map( A1 => n16915, A2 => n16838, ZN => n16825);
   U472 : CLKBUF_X1 port map( A => n16825, Z => n16826);
   U473 : OAI22_X1 port map( A1 => n18882, A2 => n16827, B1 => n16934, B2 => 
                           n16826, ZN => n1814);
   U474 : CLKBUF_X1 port map( A => n16849, Z => n16935);
   U475 : OAI22_X1 port map( A1 => n18883, A2 => n16827, B1 => n16935, B2 => 
                           n16825, ZN => n1813);
   U476 : CLKBUF_X1 port map( A => n16850, Z => n16936);
   U477 : OAI22_X1 port map( A1 => n19384, A2 => n16827, B1 => n16936, B2 => 
                           n16826, ZN => n1812);
   U478 : CLKBUF_X1 port map( A => n16851, Z => n16937);
   U479 : OAI22_X1 port map( A1 => n19134, A2 => n16827, B1 => n16937, B2 => 
                           n16825, ZN => n1811);
   U480 : CLKBUF_X1 port map( A => n16852, Z => n16938);
   U481 : OAI22_X1 port map( A1 => n18884, A2 => n16827, B1 => n16938, B2 => 
                           n16826, ZN => n1810);
   U482 : CLKBUF_X1 port map( A => n16853, Z => n16939);
   U483 : OAI22_X1 port map( A1 => n18640, A2 => n16827, B1 => n16939, B2 => 
                           n16825, ZN => n1809);
   U484 : CLKBUF_X1 port map( A => n16854, Z => n16940);
   U485 : OAI22_X1 port map( A1 => n18885, A2 => n16827, B1 => n16940, B2 => 
                           n16826, ZN => n1808);
   U486 : CLKBUF_X1 port map( A => n16855, Z => n16941);
   U487 : OAI22_X1 port map( A1 => n18886, A2 => n16827, B1 => n16941, B2 => 
                           n16825, ZN => n1807);
   U488 : CLKBUF_X1 port map( A => n16856, Z => n16942);
   U489 : OAI22_X1 port map( A1 => n19135, A2 => n16827, B1 => n16942, B2 => 
                           n16826, ZN => n1806);
   U490 : CLKBUF_X1 port map( A => n16857, Z => n16943);
   U491 : OAI22_X1 port map( A1 => n19136, A2 => n16827, B1 => n16943, B2 => 
                           n16825, ZN => n1805);
   U492 : CLKBUF_X1 port map( A => n16858, Z => n16944);
   U493 : OAI22_X1 port map( A1 => n19385, A2 => n16827, B1 => n16944, B2 => 
                           n16825, ZN => n1804);
   U494 : CLKBUF_X1 port map( A => n16859, Z => n16945);
   U495 : OAI22_X1 port map( A1 => n18641, A2 => n16827, B1 => n16945, B2 => 
                           n16826, ZN => n1803);
   U496 : OAI22_X1 port map( A1 => n19386, A2 => n16827, B1 => n16946, B2 => 
                           n16825, ZN => n1802);
   U497 : CLKBUF_X1 port map( A => n16861, Z => n16947);
   U498 : OAI22_X1 port map( A1 => n19137, A2 => n16827, B1 => n16947, B2 => 
                           n16826, ZN => n1801);
   U499 : CLKBUF_X1 port map( A => n16862, Z => n16948);
   U500 : OAI22_X1 port map( A1 => n18887, A2 => n16827, B1 => n16948, B2 => 
                           n16825, ZN => n1800);
   U501 : CLKBUF_X1 port map( A => n16863, Z => n16949);
   U502 : OAI22_X1 port map( A1 => n18888, A2 => n16827, B1 => n16949, B2 => 
                           n16826, ZN => n1799);
   U503 : CLKBUF_X1 port map( A => n16864, Z => n16950);
   U504 : OAI22_X1 port map( A1 => n18889, A2 => n16827, B1 => n16950, B2 => 
                           n16825, ZN => n1798);
   U505 : CLKBUF_X1 port map( A => n16865, Z => n16951);
   U506 : OAI22_X1 port map( A1 => n19387, A2 => n16827, B1 => n16951, B2 => 
                           n16825, ZN => n1797);
   U507 : CLKBUF_X1 port map( A => n16866, Z => n16952);
   U508 : OAI22_X1 port map( A1 => n19138, A2 => n16827, B1 => n16952, B2 => 
                           n16825, ZN => n1796);
   U509 : CLKBUF_X1 port map( A => n16867, Z => n16953);
   U510 : OAI22_X1 port map( A1 => n18642, A2 => n16827, B1 => n16953, B2 => 
                           n16825, ZN => n1795);
   U511 : CLKBUF_X1 port map( A => n16868, Z => n16954);
   U512 : OAI22_X1 port map( A1 => n19388, A2 => n16827, B1 => n16954, B2 => 
                           n16825, ZN => n1794);
   U513 : CLKBUF_X1 port map( A => n16869, Z => n16955);
   U514 : OAI22_X1 port map( A1 => n19139, A2 => n16827, B1 => n16955, B2 => 
                           n16825, ZN => n1793);
   U515 : CLKBUF_X1 port map( A => n16871, Z => n16957);
   U516 : OAI22_X1 port map( A1 => n18890, A2 => n16827, B1 => n16957, B2 => 
                           n16825, ZN => n1792);
   U517 : CLKBUF_X1 port map( A => n16872, Z => n16958);
   U518 : OAI22_X1 port map( A1 => n18891, A2 => n16827, B1 => n16958, B2 => 
                           n16826, ZN => n1791);
   U519 : CLKBUF_X1 port map( A => n16873, Z => n16959);
   U520 : OAI22_X1 port map( A1 => n18892, A2 => n16827, B1 => n16959, B2 => 
                           n16826, ZN => n1790);
   U521 : CLKBUF_X1 port map( A => n16874, Z => n16960);
   U522 : OAI22_X1 port map( A1 => n19140, A2 => n16827, B1 => n16960, B2 => 
                           n16826, ZN => n1789);
   U523 : CLKBUF_X1 port map( A => n16875, Z => n16961);
   U524 : OAI22_X1 port map( A1 => n18893, A2 => n16827, B1 => n16961, B2 => 
                           n16826, ZN => n1788);
   U525 : OAI22_X1 port map( A1 => n19389, A2 => n16827, B1 => n16962, B2 => 
                           n16826, ZN => n1787);
   U526 : CLKBUF_X1 port map( A => n16877, Z => n16963);
   U527 : OAI22_X1 port map( A1 => n18894, A2 => n16827, B1 => n16963, B2 => 
                           n16826, ZN => n1786);
   U528 : CLKBUF_X1 port map( A => n16878, Z => n16964);
   U529 : OAI22_X1 port map( A1 => n18643, A2 => n16827, B1 => n16964, B2 => 
                           n16826, ZN => n1785);
   U530 : CLKBUF_X1 port map( A => n16879, Z => n16965);
   U531 : OAI22_X1 port map( A1 => n19141, A2 => n16827, B1 => n16965, B2 => 
                           n16826, ZN => n1784);
   U532 : CLKBUF_X1 port map( A => n16881, Z => n16967);
   U533 : OAI22_X1 port map( A1 => n19142, A2 => n16827, B1 => n16967, B2 => 
                           n16826, ZN => n1783);
   U534 : NAND2_X1 port map( A1 => n16919, A2 => n16838, ZN => n16828);
   U535 : CLKBUF_X1 port map( A => n16828, Z => n16829);
   U536 : OAI22_X1 port map( A1 => n18644, A2 => n16830, B1 => n16896, B2 => 
                           n16829, ZN => n1782);
   U537 : OAI22_X1 port map( A1 => n19390, A2 => n16830, B1 => n16849, B2 => 
                           n16828, ZN => n1781);
   U538 : OAI22_X1 port map( A1 => n18895, A2 => n16830, B1 => n16850, B2 => 
                           n16829, ZN => n1780);
   U539 : OAI22_X1 port map( A1 => n19143, A2 => n16830, B1 => n16851, B2 => 
                           n16828, ZN => n1779);
   U540 : OAI22_X1 port map( A1 => n19391, A2 => n16830, B1 => n16852, B2 => 
                           n16829, ZN => n1778);
   U541 : OAI22_X1 port map( A1 => n19144, A2 => n16830, B1 => n16853, B2 => 
                           n16828, ZN => n1777);
   U542 : OAI22_X1 port map( A1 => n19392, A2 => n16830, B1 => n16854, B2 => 
                           n16829, ZN => n1776);
   U543 : OAI22_X1 port map( A1 => n19393, A2 => n16830, B1 => n16855, B2 => 
                           n16828, ZN => n1775);
   U544 : OAI22_X1 port map( A1 => n19394, A2 => n16830, B1 => n16856, B2 => 
                           n16829, ZN => n1774);
   U545 : OAI22_X1 port map( A1 => n18896, A2 => n16830, B1 => n16857, B2 => 
                           n16828, ZN => n1773);
   U546 : OAI22_X1 port map( A1 => n19395, A2 => n16830, B1 => n16858, B2 => 
                           n16828, ZN => n1772);
   U547 : OAI22_X1 port map( A1 => n19145, A2 => n16830, B1 => n16859, B2 => 
                           n16829, ZN => n1771);
   U548 : OAI22_X1 port map( A1 => n19146, A2 => n16830, B1 => n16860, B2 => 
                           n16828, ZN => n1770);
   U549 : OAI22_X1 port map( A1 => n19396, A2 => n16830, B1 => n16861, B2 => 
                           n16829, ZN => n1769);
   U550 : OAI22_X1 port map( A1 => n18897, A2 => n16830, B1 => n16862, B2 => 
                           n16828, ZN => n1768);
   U551 : OAI22_X1 port map( A1 => n19397, A2 => n16830, B1 => n16863, B2 => 
                           n16829, ZN => n1767);
   U552 : OAI22_X1 port map( A1 => n18645, A2 => n16830, B1 => n16864, B2 => 
                           n16828, ZN => n1766);
   U553 : OAI22_X1 port map( A1 => n18898, A2 => n16830, B1 => n16865, B2 => 
                           n16828, ZN => n1765);
   U554 : OAI22_X1 port map( A1 => n18646, A2 => n16830, B1 => n16866, B2 => 
                           n16828, ZN => n1764);
   U555 : OAI22_X1 port map( A1 => n18899, A2 => n16830, B1 => n16867, B2 => 
                           n16828, ZN => n1763);
   U556 : OAI22_X1 port map( A1 => n18900, A2 => n16830, B1 => n16868, B2 => 
                           n16828, ZN => n1762);
   U557 : OAI22_X1 port map( A1 => n19147, A2 => n16830, B1 => n16869, B2 => 
                           n16828, ZN => n1761);
   U558 : OAI22_X1 port map( A1 => n19148, A2 => n16830, B1 => n16871, B2 => 
                           n16828, ZN => n1760);
   U559 : OAI22_X1 port map( A1 => n19398, A2 => n16830, B1 => n16872, B2 => 
                           n16829, ZN => n1759);
   U560 : OAI22_X1 port map( A1 => n19149, A2 => n16830, B1 => n16873, B2 => 
                           n16829, ZN => n1758);
   U561 : OAI22_X1 port map( A1 => n19399, A2 => n16830, B1 => n16874, B2 => 
                           n16829, ZN => n1757);
   U562 : OAI22_X1 port map( A1 => n19150, A2 => n16830, B1 => n16875, B2 => 
                           n16829, ZN => n1756);
   U563 : OAI22_X1 port map( A1 => n18647, A2 => n16830, B1 => n16876, B2 => 
                           n16829, ZN => n1755);
   U564 : OAI22_X1 port map( A1 => n18648, A2 => n16830, B1 => n16877, B2 => 
                           n16829, ZN => n1754);
   U565 : OAI22_X1 port map( A1 => n19151, A2 => n16830, B1 => n16878, B2 => 
                           n16829, ZN => n1753);
   U566 : OAI22_X1 port map( A1 => n19152, A2 => n16830, B1 => n16879, B2 => 
                           n16829, ZN => n1752);
   U567 : OAI22_X1 port map( A1 => n19400, A2 => n16830, B1 => n16881, B2 => 
                           n16829, ZN => n1751);
   U568 : NAND2_X1 port map( A1 => n16923, A2 => n16838, ZN => n16831);
   U569 : CLKBUF_X1 port map( A => n16831, Z => n16832);
   U570 : OAI22_X1 port map( A1 => n19153, A2 => n16833, B1 => n16896, B2 => 
                           n16832, ZN => n1750);
   U571 : OAI22_X1 port map( A1 => n18649, A2 => n16833, B1 => n16935, B2 => 
                           n16831, ZN => n1749);
   U572 : OAI22_X1 port map( A1 => n19154, A2 => n16833, B1 => n16936, B2 => 
                           n16832, ZN => n1748);
   U573 : OAI22_X1 port map( A1 => n19155, A2 => n16833, B1 => n16937, B2 => 
                           n16831, ZN => n1747);
   U574 : OAI22_X1 port map( A1 => n18901, A2 => n16833, B1 => n16938, B2 => 
                           n16832, ZN => n1746);
   U575 : OAI22_X1 port map( A1 => n19401, A2 => n16833, B1 => n16939, B2 => 
                           n16831, ZN => n1745);
   U576 : OAI22_X1 port map( A1 => n19156, A2 => n16833, B1 => n16940, B2 => 
                           n16832, ZN => n1744);
   U577 : OAI22_X1 port map( A1 => n19157, A2 => n16833, B1 => n16941, B2 => 
                           n16831, ZN => n1743);
   U578 : OAI22_X1 port map( A1 => n18902, A2 => n16833, B1 => n16942, B2 => 
                           n16832, ZN => n1742);
   U579 : OAI22_X1 port map( A1 => n19402, A2 => n16833, B1 => n16943, B2 => 
                           n16831, ZN => n1741);
   U580 : OAI22_X1 port map( A1 => n19403, A2 => n16833, B1 => n16944, B2 => 
                           n16831, ZN => n1740);
   U581 : OAI22_X1 port map( A1 => n19404, A2 => n16833, B1 => n16945, B2 => 
                           n16832, ZN => n1739);
   U582 : OAI22_X1 port map( A1 => n18903, A2 => n16833, B1 => n16946, B2 => 
                           n16831, ZN => n1738);
   U583 : OAI22_X1 port map( A1 => n19405, A2 => n16833, B1 => n16947, B2 => 
                           n16832, ZN => n1737);
   U584 : OAI22_X1 port map( A1 => n19158, A2 => n16833, B1 => n16948, B2 => 
                           n16831, ZN => n1736);
   U585 : OAI22_X1 port map( A1 => n19159, A2 => n16833, B1 => n16949, B2 => 
                           n16832, ZN => n1735);
   U586 : OAI22_X1 port map( A1 => n19406, A2 => n16833, B1 => n16950, B2 => 
                           n16831, ZN => n1734);
   U587 : OAI22_X1 port map( A1 => n19160, A2 => n16833, B1 => n16951, B2 => 
                           n16831, ZN => n1733);
   U588 : OAI22_X1 port map( A1 => n19407, A2 => n16833, B1 => n16952, B2 => 
                           n16831, ZN => n1732);
   U589 : OAI22_X1 port map( A1 => n19161, A2 => n16833, B1 => n16953, B2 => 
                           n16831, ZN => n1731);
   U590 : OAI22_X1 port map( A1 => n19162, A2 => n16833, B1 => n16954, B2 => 
                           n16831, ZN => n1730);
   U591 : OAI22_X1 port map( A1 => n19408, A2 => n16833, B1 => n16955, B2 => 
                           n16831, ZN => n1729);
   U592 : OAI22_X1 port map( A1 => n19409, A2 => n16833, B1 => n16957, B2 => 
                           n16831, ZN => n1728);
   U593 : OAI22_X1 port map( A1 => n19163, A2 => n16833, B1 => n16958, B2 => 
                           n16832, ZN => n1727);
   U594 : OAI22_X1 port map( A1 => n18650, A2 => n16833, B1 => n16959, B2 => 
                           n16832, ZN => n1726);
   U595 : OAI22_X1 port map( A1 => n19410, A2 => n16833, B1 => n16960, B2 => 
                           n16832, ZN => n1725);
   U596 : OAI22_X1 port map( A1 => n19411, A2 => n16833, B1 => n16961, B2 => 
                           n16832, ZN => n1724);
   U597 : OAI22_X1 port map( A1 => n19412, A2 => n16833, B1 => n16962, B2 => 
                           n16832, ZN => n1723);
   U598 : OAI22_X1 port map( A1 => n19164, A2 => n16833, B1 => n16963, B2 => 
                           n16832, ZN => n1722);
   U599 : OAI22_X1 port map( A1 => n19413, A2 => n16833, B1 => n16964, B2 => 
                           n16832, ZN => n1721);
   U600 : OAI22_X1 port map( A1 => n19414, A2 => n16833, B1 => n16965, B2 => 
                           n16832, ZN => n1720);
   U601 : OAI22_X1 port map( A1 => n19415, A2 => n16833, B1 => n16967, B2 => 
                           n16832, ZN => n1719);
   U602 : NAND2_X1 port map( A1 => n16928, A2 => n16838, ZN => n16834);
   U603 : CLKBUF_X1 port map( A => n16837, Z => n16835);
   U604 : CLKBUF_X1 port map( A => n16834, Z => n16836);
   U605 : OAI22_X1 port map( A1 => n19416, A2 => n16835, B1 => n16896, B2 => 
                           n16836, ZN => n1718);
   U606 : OAI22_X1 port map( A1 => n19165, A2 => n16837, B1 => n16849, B2 => 
                           n16834, ZN => n1717);
   U607 : OAI22_X1 port map( A1 => n19166, A2 => n16835, B1 => n16850, B2 => 
                           n16836, ZN => n1716);
   U608 : OAI22_X1 port map( A1 => n19417, A2 => n16837, B1 => n16851, B2 => 
                           n16834, ZN => n1715);
   U609 : OAI22_X1 port map( A1 => n19418, A2 => n16835, B1 => n16852, B2 => 
                           n16836, ZN => n1714);
   U610 : OAI22_X1 port map( A1 => n19167, A2 => n16837, B1 => n16853, B2 => 
                           n16834, ZN => n1713);
   U611 : OAI22_X1 port map( A1 => n19168, A2 => n16835, B1 => n16854, B2 => 
                           n16836, ZN => n1712);
   U612 : OAI22_X1 port map( A1 => n19419, A2 => n16837, B1 => n16855, B2 => 
                           n16834, ZN => n1711);
   U613 : OAI22_X1 port map( A1 => n19169, A2 => n16835, B1 => n16856, B2 => 
                           n16836, ZN => n1710);
   U614 : OAI22_X1 port map( A1 => n19420, A2 => n16837, B1 => n16857, B2 => 
                           n16834, ZN => n1709);
   U615 : OAI22_X1 port map( A1 => n19170, A2 => n16837, B1 => n16858, B2 => 
                           n16834, ZN => n1708);
   U616 : OAI22_X1 port map( A1 => n19171, A2 => n16837, B1 => n16859, B2 => 
                           n16836, ZN => n1707);
   U617 : OAI22_X1 port map( A1 => n19421, A2 => n16835, B1 => n16860, B2 => 
                           n16834, ZN => n1706);
   U618 : OAI22_X1 port map( A1 => n19172, A2 => n16835, B1 => n16861, B2 => 
                           n16836, ZN => n1705);
   U619 : OAI22_X1 port map( A1 => n19173, A2 => n16835, B1 => n16862, B2 => 
                           n16834, ZN => n1704);
   U620 : OAI22_X1 port map( A1 => n19174, A2 => n16835, B1 => n16863, B2 => 
                           n16836, ZN => n1703);
   U621 : OAI22_X1 port map( A1 => n19175, A2 => n16835, B1 => n16864, B2 => 
                           n16834, ZN => n1702);
   U622 : OAI22_X1 port map( A1 => n19176, A2 => n16835, B1 => n16865, B2 => 
                           n16834, ZN => n1701);
   U623 : OAI22_X1 port map( A1 => n19177, A2 => n16835, B1 => n16866, B2 => 
                           n16834, ZN => n1700);
   U624 : OAI22_X1 port map( A1 => n19422, A2 => n16835, B1 => n16867, B2 => 
                           n16834, ZN => n1699);
   U625 : OAI22_X1 port map( A1 => n19423, A2 => n16835, B1 => n16868, B2 => 
                           n16834, ZN => n1698);
   U626 : OAI22_X1 port map( A1 => n19424, A2 => n16835, B1 => n16869, B2 => 
                           n16834, ZN => n1697);
   U627 : OAI22_X1 port map( A1 => n19425, A2 => n16835, B1 => n16871, B2 => 
                           n16834, ZN => n1696);
   U628 : OAI22_X1 port map( A1 => n19426, A2 => n16835, B1 => n16872, B2 => 
                           n16836, ZN => n1695);
   U629 : OAI22_X1 port map( A1 => n19178, A2 => n16837, B1 => n16873, B2 => 
                           n16836, ZN => n1694);
   U630 : OAI22_X1 port map( A1 => n19179, A2 => n16837, B1 => n16874, B2 => 
                           n16836, ZN => n1693);
   U631 : OAI22_X1 port map( A1 => n19180, A2 => n16837, B1 => n16875, B2 => 
                           n16836, ZN => n1692);
   U632 : OAI22_X1 port map( A1 => n19181, A2 => n16837, B1 => n16876, B2 => 
                           n16836, ZN => n1691);
   U633 : OAI22_X1 port map( A1 => n19427, A2 => n16837, B1 => n16877, B2 => 
                           n16836, ZN => n1690);
   U634 : OAI22_X1 port map( A1 => n19182, A2 => n16837, B1 => n16878, B2 => 
                           n16836, ZN => n1689);
   U635 : OAI22_X1 port map( A1 => n19428, A2 => n16837, B1 => n16879, B2 => 
                           n16836, ZN => n1688);
   U636 : OAI22_X1 port map( A1 => n19183, A2 => n16837, B1 => n16881, B2 => 
                           n16836, ZN => n1687);
   U637 : NAND2_X1 port map( A1 => n16933, A2 => n16838, ZN => n16839);
   U638 : CLKBUF_X1 port map( A => n16839, Z => n16840);
   U639 : OAI22_X1 port map( A1 => n18651, A2 => n16841, B1 => n16896, B2 => 
                           n16840, ZN => n1686);
   U640 : OAI22_X1 port map( A1 => n18904, A2 => n16841, B1 => n16935, B2 => 
                           n16839, ZN => n1685);
   U641 : OAI22_X1 port map( A1 => n18905, A2 => n16841, B1 => n16936, B2 => 
                           n16840, ZN => n1684);
   U642 : OAI22_X1 port map( A1 => n18906, A2 => n16841, B1 => n16937, B2 => 
                           n16839, ZN => n1683);
   U643 : OAI22_X1 port map( A1 => n18652, A2 => n16841, B1 => n16938, B2 => 
                           n16840, ZN => n1682);
   U644 : OAI22_X1 port map( A1 => n18907, A2 => n16841, B1 => n16939, B2 => 
                           n16839, ZN => n1681);
   U645 : OAI22_X1 port map( A1 => n18908, A2 => n16841, B1 => n16940, B2 => 
                           n16840, ZN => n1680);
   U646 : OAI22_X1 port map( A1 => n18653, A2 => n16841, B1 => n16941, B2 => 
                           n16839, ZN => n1679);
   U647 : OAI22_X1 port map( A1 => n18909, A2 => n16841, B1 => n16942, B2 => 
                           n16840, ZN => n1678);
   U648 : OAI22_X1 port map( A1 => n18654, A2 => n16841, B1 => n16943, B2 => 
                           n16839, ZN => n1677);
   U649 : OAI22_X1 port map( A1 => n18655, A2 => n16841, B1 => n16944, B2 => 
                           n16839, ZN => n1676);
   U650 : OAI22_X1 port map( A1 => n18656, A2 => n16841, B1 => n16945, B2 => 
                           n16840, ZN => n1675);
   U651 : OAI22_X1 port map( A1 => n18910, A2 => n16841, B1 => n16946, B2 => 
                           n16839, ZN => n1674);
   U652 : OAI22_X1 port map( A1 => n18657, A2 => n16841, B1 => n16947, B2 => 
                           n16840, ZN => n1673);
   U653 : OAI22_X1 port map( A1 => n18911, A2 => n16841, B1 => n16948, B2 => 
                           n16839, ZN => n1672);
   U654 : OAI22_X1 port map( A1 => n18912, A2 => n16841, B1 => n16949, B2 => 
                           n16840, ZN => n1671);
   U655 : OAI22_X1 port map( A1 => n18913, A2 => n16841, B1 => n16950, B2 => 
                           n16839, ZN => n1670);
   U656 : OAI22_X1 port map( A1 => n18914, A2 => n16841, B1 => n16951, B2 => 
                           n16839, ZN => n1669);
   U657 : OAI22_X1 port map( A1 => n18915, A2 => n16841, B1 => n16952, B2 => 
                           n16839, ZN => n1668);
   U658 : OAI22_X1 port map( A1 => n18916, A2 => n16841, B1 => n16953, B2 => 
                           n16839, ZN => n1667);
   U659 : OAI22_X1 port map( A1 => n18917, A2 => n16841, B1 => n16954, B2 => 
                           n16839, ZN => n1666);
   U660 : OAI22_X1 port map( A1 => n18918, A2 => n16841, B1 => n16955, B2 => 
                           n16839, ZN => n1665);
   U661 : OAI22_X1 port map( A1 => n18658, A2 => n16841, B1 => n16957, B2 => 
                           n16839, ZN => n1664);
   U662 : OAI22_X1 port map( A1 => n18919, A2 => n16841, B1 => n16958, B2 => 
                           n16840, ZN => n1663);
   U663 : OAI22_X1 port map( A1 => n18920, A2 => n16841, B1 => n16959, B2 => 
                           n16840, ZN => n1662);
   U664 : OAI22_X1 port map( A1 => n18659, A2 => n16841, B1 => n16960, B2 => 
                           n16840, ZN => n1661);
   U665 : OAI22_X1 port map( A1 => n18660, A2 => n16841, B1 => n16961, B2 => 
                           n16840, ZN => n1660);
   U666 : OAI22_X1 port map( A1 => n18921, A2 => n16841, B1 => n16962, B2 => 
                           n16840, ZN => n1659);
   U667 : OAI22_X1 port map( A1 => n18922, A2 => n16841, B1 => n16963, B2 => 
                           n16840, ZN => n1658);
   U668 : OAI22_X1 port map( A1 => n18923, A2 => n16841, B1 => n16964, B2 => 
                           n16840, ZN => n1657);
   U669 : OAI22_X1 port map( A1 => n18924, A2 => n16841, B1 => n16965, B2 => 
                           n16840, ZN => n1656);
   U670 : OAI22_X1 port map( A1 => n18925, A2 => n16841, B1 => n16967, B2 => 
                           n16840, ZN => n1655);
   U671 : NOR2_X1 port map( A1 => n16901, A2 => n16842, ZN => n16895);
   U672 : NAND2_X1 port map( A1 => n16902, A2 => n16895, ZN => n16843);
   U673 : CLKBUF_X1 port map( A => n16843, Z => n16844);
   U674 : OAI22_X1 port map( A1 => n18788, A2 => n16845, B1 => n16896, B2 => 
                           n16844, ZN => n1654);
   U675 : OAI22_X1 port map( A1 => n19429, A2 => n16845, B1 => n16849, B2 => 
                           n16843, ZN => n1653);
   U676 : OAI22_X1 port map( A1 => n19184, A2 => n16845, B1 => n16850, B2 => 
                           n16844, ZN => n1652);
   U677 : OAI22_X1 port map( A1 => n18926, A2 => n16845, B1 => n16851, B2 => 
                           n16843, ZN => n1651);
   U678 : OAI22_X1 port map( A1 => n19185, A2 => n16845, B1 => n16852, B2 => 
                           n16844, ZN => n1650);
   U679 : OAI22_X1 port map( A1 => n19430, A2 => n16845, B1 => n16853, B2 => 
                           n16843, ZN => n1649);
   U680 : OAI22_X1 port map( A1 => n19431, A2 => n16845, B1 => n16854, B2 => 
                           n16844, ZN => n1648);
   U681 : OAI22_X1 port map( A1 => n19432, A2 => n16845, B1 => n16855, B2 => 
                           n16843, ZN => n1647);
   U682 : OAI22_X1 port map( A1 => n18927, A2 => n16845, B1 => n16856, B2 => 
                           n16844, ZN => n1646);
   U683 : OAI22_X1 port map( A1 => n18661, A2 => n16845, B1 => n16857, B2 => 
                           n16843, ZN => n1645);
   U684 : OAI22_X1 port map( A1 => n19186, A2 => n16845, B1 => n16858, B2 => 
                           n16843, ZN => n1644);
   U685 : OAI22_X1 port map( A1 => n19433, A2 => n16845, B1 => n16859, B2 => 
                           n16844, ZN => n1643);
   U686 : OAI22_X1 port map( A1 => n18662, A2 => n16845, B1 => n16860, B2 => 
                           n16843, ZN => n1642);
   U687 : OAI22_X1 port map( A1 => n19187, A2 => n16845, B1 => n16861, B2 => 
                           n16844, ZN => n1641);
   U688 : OAI22_X1 port map( A1 => n18928, A2 => n16845, B1 => n16862, B2 => 
                           n16843, ZN => n1640);
   U689 : OAI22_X1 port map( A1 => n18929, A2 => n16845, B1 => n16863, B2 => 
                           n16844, ZN => n1639);
   U690 : OAI22_X1 port map( A1 => n19188, A2 => n16845, B1 => n16864, B2 => 
                           n16843, ZN => n1638);
   U691 : OAI22_X1 port map( A1 => n19189, A2 => n16845, B1 => n16865, B2 => 
                           n16843, ZN => n1637);
   U692 : OAI22_X1 port map( A1 => n19434, A2 => n16845, B1 => n16866, B2 => 
                           n16843, ZN => n1636);
   U693 : OAI22_X1 port map( A1 => n19190, A2 => n16845, B1 => n16867, B2 => 
                           n16843, ZN => n1635);
   U694 : OAI22_X1 port map( A1 => n18663, A2 => n16845, B1 => n16868, B2 => 
                           n16843, ZN => n1634);
   U695 : OAI22_X1 port map( A1 => n19435, A2 => n16845, B1 => n16869, B2 => 
                           n16843, ZN => n1633);
   U696 : OAI22_X1 port map( A1 => n18930, A2 => n16845, B1 => n16871, B2 => 
                           n16843, ZN => n1632);
   U697 : OAI22_X1 port map( A1 => n19191, A2 => n16845, B1 => n16872, B2 => 
                           n16844, ZN => n1631);
   U698 : OAI22_X1 port map( A1 => n19436, A2 => n16845, B1 => n16873, B2 => 
                           n16844, ZN => n1630);
   U699 : OAI22_X1 port map( A1 => n18664, A2 => n16845, B1 => n16874, B2 => 
                           n16844, ZN => n1629);
   U700 : OAI22_X1 port map( A1 => n19437, A2 => n16845, B1 => n16875, B2 => 
                           n16844, ZN => n1628);
   U701 : OAI22_X1 port map( A1 => n18665, A2 => n16845, B1 => n16876, B2 => 
                           n16844, ZN => n1627);
   U702 : OAI22_X1 port map( A1 => n19192, A2 => n16845, B1 => n16877, B2 => 
                           n16844, ZN => n1626);
   U703 : OAI22_X1 port map( A1 => n18931, A2 => n16845, B1 => n16878, B2 => 
                           n16844, ZN => n1625);
   U704 : OAI22_X1 port map( A1 => n18932, A2 => n16845, B1 => n16879, B2 => 
                           n16844, ZN => n1624);
   U705 : OAI22_X1 port map( A1 => n18933, A2 => n16845, B1 => n16881, B2 => 
                           n16844, ZN => n1623);
   U706 : NAND2_X1 port map( A1 => n16906, A2 => n16895, ZN => n16846);
   U707 : CLKBUF_X1 port map( A => n16846, Z => n16847);
   U708 : OAI22_X1 port map( A1 => n18532, A2 => n16848, B1 => n16896, B2 => 
                           n16847, ZN => n1622);
   U709 : OAI22_X1 port map( A1 => n18934, A2 => n16848, B1 => n16935, B2 => 
                           n16846, ZN => n1621);
   U710 : OAI22_X1 port map( A1 => n18666, A2 => n16848, B1 => n16936, B2 => 
                           n16847, ZN => n1620);
   U711 : OAI22_X1 port map( A1 => n18935, A2 => n16848, B1 => n16937, B2 => 
                           n16846, ZN => n1619);
   U712 : OAI22_X1 port map( A1 => n19438, A2 => n16848, B1 => n16938, B2 => 
                           n16847, ZN => n1618);
   U713 : OAI22_X1 port map( A1 => n18667, A2 => n16848, B1 => n16939, B2 => 
                           n16846, ZN => n1617);
   U714 : OAI22_X1 port map( A1 => n18936, A2 => n16848, B1 => n16940, B2 => 
                           n16847, ZN => n1616);
   U715 : OAI22_X1 port map( A1 => n19193, A2 => n16848, B1 => n16941, B2 => 
                           n16846, ZN => n1615);
   U716 : OAI22_X1 port map( A1 => n19194, A2 => n16848, B1 => n16942, B2 => 
                           n16847, ZN => n1614);
   U717 : OAI22_X1 port map( A1 => n18937, A2 => n16848, B1 => n16943, B2 => 
                           n16846, ZN => n1613);
   U718 : OAI22_X1 port map( A1 => n19439, A2 => n16848, B1 => n16944, B2 => 
                           n16846, ZN => n1612);
   U719 : OAI22_X1 port map( A1 => n19195, A2 => n16848, B1 => n16945, B2 => 
                           n16847, ZN => n1611);
   U720 : OAI22_X1 port map( A1 => n19196, A2 => n16848, B1 => n16946, B2 => 
                           n16846, ZN => n1610);
   U721 : OAI22_X1 port map( A1 => n19440, A2 => n16848, B1 => n16947, B2 => 
                           n16847, ZN => n1609);
   U722 : OAI22_X1 port map( A1 => n19197, A2 => n16848, B1 => n16948, B2 => 
                           n16846, ZN => n1608);
   U723 : OAI22_X1 port map( A1 => n18668, A2 => n16848, B1 => n16949, B2 => 
                           n16847, ZN => n1607);
   U724 : OAI22_X1 port map( A1 => n18669, A2 => n16848, B1 => n16950, B2 => 
                           n16846, ZN => n1606);
   U725 : OAI22_X1 port map( A1 => n19198, A2 => n16848, B1 => n16951, B2 => 
                           n16846, ZN => n1605);
   U726 : OAI22_X1 port map( A1 => n19199, A2 => n16848, B1 => n16952, B2 => 
                           n16846, ZN => n1604);
   U727 : OAI22_X1 port map( A1 => n19200, A2 => n16848, B1 => n16953, B2 => 
                           n16846, ZN => n1603);
   U728 : OAI22_X1 port map( A1 => n18670, A2 => n16848, B1 => n16954, B2 => 
                           n16846, ZN => n1602);
   U729 : OAI22_X1 port map( A1 => n18938, A2 => n16848, B1 => n16955, B2 => 
                           n16846, ZN => n1601);
   U730 : OAI22_X1 port map( A1 => n18939, A2 => n16848, B1 => n16957, B2 => 
                           n16846, ZN => n1600);
   U731 : OAI22_X1 port map( A1 => n19441, A2 => n16848, B1 => n16958, B2 => 
                           n16847, ZN => n1599);
   U732 : OAI22_X1 port map( A1 => n19442, A2 => n16848, B1 => n16959, B2 => 
                           n16847, ZN => n1598);
   U733 : OAI22_X1 port map( A1 => n19443, A2 => n16848, B1 => n16960, B2 => 
                           n16847, ZN => n1597);
   U734 : OAI22_X1 port map( A1 => n18940, A2 => n16848, B1 => n16961, B2 => 
                           n16847, ZN => n1596);
   U735 : OAI22_X1 port map( A1 => n19201, A2 => n16848, B1 => n16962, B2 => 
                           n16847, ZN => n1595);
   U736 : OAI22_X1 port map( A1 => n19444, A2 => n16848, B1 => n16963, B2 => 
                           n16847, ZN => n1594);
   U737 : OAI22_X1 port map( A1 => n18941, A2 => n16848, B1 => n16964, B2 => 
                           n16847, ZN => n1593);
   U738 : OAI22_X1 port map( A1 => n19445, A2 => n16848, B1 => n16965, B2 => 
                           n16847, ZN => n1592);
   U739 : OAI22_X1 port map( A1 => n18942, A2 => n16848, B1 => n16967, B2 => 
                           n16847, ZN => n1591);
   U740 : NAND2_X1 port map( A1 => n16911, A2 => n16895, ZN => n16870);
   U741 : OAI22_X1 port map( A1 => n18533, A2 => n16882, B1 => n16896, B2 => 
                           n16880, ZN => n1590);
   U742 : OAI22_X1 port map( A1 => n18671, A2 => n16882, B1 => n16849, B2 => 
                           n16870, ZN => n1589);
   U743 : OAI22_X1 port map( A1 => n18672, A2 => n16882, B1 => n16850, B2 => 
                           n16880, ZN => n1588);
   U744 : OAI22_X1 port map( A1 => n18673, A2 => n16882, B1 => n16851, B2 => 
                           n16870, ZN => n1587);
   U745 : OAI22_X1 port map( A1 => n18674, A2 => n16882, B1 => n16852, B2 => 
                           n16880, ZN => n1586);
   U746 : OAI22_X1 port map( A1 => n19202, A2 => n16882, B1 => n16853, B2 => 
                           n16870, ZN => n1585);
   U747 : OAI22_X1 port map( A1 => n19446, A2 => n16882, B1 => n16854, B2 => 
                           n16880, ZN => n1584);
   U748 : OAI22_X1 port map( A1 => n18943, A2 => n16882, B1 => n16855, B2 => 
                           n16870, ZN => n1583);
   U749 : OAI22_X1 port map( A1 => n18675, A2 => n16882, B1 => n16856, B2 => 
                           n16880, ZN => n1582);
   U750 : OAI22_X1 port map( A1 => n19447, A2 => n16882, B1 => n16857, B2 => 
                           n16870, ZN => n1581);
   U751 : OAI22_X1 port map( A1 => n18944, A2 => n16882, B1 => n16858, B2 => 
                           n16870, ZN => n1580);
   U752 : OAI22_X1 port map( A1 => n18676, A2 => n16882, B1 => n16859, B2 => 
                           n16880, ZN => n1579);
   U753 : OAI22_X1 port map( A1 => n19448, A2 => n16882, B1 => n16860, B2 => 
                           n16870, ZN => n1578);
   U754 : OAI22_X1 port map( A1 => n18677, A2 => n16882, B1 => n16861, B2 => 
                           n16880, ZN => n1577);
   U755 : OAI22_X1 port map( A1 => n18945, A2 => n16882, B1 => n16862, B2 => 
                           n16870, ZN => n1576);
   U756 : OAI22_X1 port map( A1 => n19449, A2 => n16882, B1 => n16863, B2 => 
                           n16880, ZN => n1575);
   U757 : OAI22_X1 port map( A1 => n19450, A2 => n16882, B1 => n16864, B2 => 
                           n16870, ZN => n1574);
   U758 : OAI22_X1 port map( A1 => n19451, A2 => n16882, B1 => n16865, B2 => 
                           n16870, ZN => n1573);
   U759 : OAI22_X1 port map( A1 => n18678, A2 => n16882, B1 => n16866, B2 => 
                           n16870, ZN => n1572);
   U760 : OAI22_X1 port map( A1 => n18679, A2 => n16882, B1 => n16867, B2 => 
                           n16870, ZN => n1571);
   U761 : OAI22_X1 port map( A1 => n19452, A2 => n16882, B1 => n16868, B2 => 
                           n16870, ZN => n1570);
   U762 : OAI22_X1 port map( A1 => n19453, A2 => n16882, B1 => n16869, B2 => 
                           n16870, ZN => n1569);
   U763 : OAI22_X1 port map( A1 => n18680, A2 => n16882, B1 => n16871, B2 => 
                           n16870, ZN => n1568);
   U764 : OAI22_X1 port map( A1 => n18681, A2 => n16882, B1 => n16872, B2 => 
                           n16880, ZN => n1567);
   U765 : OAI22_X1 port map( A1 => n18946, A2 => n16882, B1 => n16873, B2 => 
                           n16880, ZN => n1566);
   U766 : OAI22_X1 port map( A1 => n18682, A2 => n16882, B1 => n16874, B2 => 
                           n16880, ZN => n1565);
   U767 : OAI22_X1 port map( A1 => n18683, A2 => n16882, B1 => n16875, B2 => 
                           n16880, ZN => n1564);
   U768 : OAI22_X1 port map( A1 => n19203, A2 => n16882, B1 => n16876, B2 => 
                           n16880, ZN => n1563);
   U769 : OAI22_X1 port map( A1 => n18947, A2 => n16882, B1 => n16877, B2 => 
                           n16880, ZN => n1562);
   U770 : OAI22_X1 port map( A1 => n19454, A2 => n16882, B1 => n16878, B2 => 
                           n16880, ZN => n1561);
   U771 : OAI22_X1 port map( A1 => n18948, A2 => n16882, B1 => n16879, B2 => 
                           n16880, ZN => n1560);
   U772 : OAI22_X1 port map( A1 => n18684, A2 => n16882, B1 => n16881, B2 => 
                           n16880, ZN => n1559);
   U773 : NAND2_X1 port map( A1 => n16915, A2 => n16895, ZN => n16883);
   U774 : CLKBUF_X1 port map( A => n16883, Z => n16884);
   U775 : OAI22_X1 port map( A1 => n18534, A2 => n16885, B1 => n16896, B2 => 
                           n16884, ZN => n1558);
   U776 : OAI22_X1 port map( A1 => n19204, A2 => n16885, B1 => n16935, B2 => 
                           n16883, ZN => n1557);
   U777 : OAI22_X1 port map( A1 => n18685, A2 => n16885, B1 => n16936, B2 => 
                           n16884, ZN => n1556);
   U778 : OAI22_X1 port map( A1 => n19205, A2 => n16885, B1 => n16937, B2 => 
                           n16883, ZN => n1555);
   U779 : OAI22_X1 port map( A1 => n18686, A2 => n16885, B1 => n16938, B2 => 
                           n16884, ZN => n1554);
   U780 : OAI22_X1 port map( A1 => n18687, A2 => n16885, B1 => n16939, B2 => 
                           n16883, ZN => n1553);
   U781 : OAI22_X1 port map( A1 => n18688, A2 => n16885, B1 => n16940, B2 => 
                           n16884, ZN => n1552);
   U782 : OAI22_X1 port map( A1 => n19206, A2 => n16885, B1 => n16941, B2 => 
                           n16883, ZN => n1551);
   U783 : OAI22_X1 port map( A1 => n18689, A2 => n16885, B1 => n16942, B2 => 
                           n16884, ZN => n1550);
   U784 : OAI22_X1 port map( A1 => n18690, A2 => n16885, B1 => n16943, B2 => 
                           n16883, ZN => n1549);
   U785 : OAI22_X1 port map( A1 => n18691, A2 => n16885, B1 => n16944, B2 => 
                           n16883, ZN => n1548);
   U786 : OAI22_X1 port map( A1 => n19455, A2 => n16885, B1 => n16945, B2 => 
                           n16884, ZN => n1547);
   U787 : OAI22_X1 port map( A1 => n18692, A2 => n16885, B1 => n16946, B2 => 
                           n16883, ZN => n1546);
   U788 : OAI22_X1 port map( A1 => n18693, A2 => n16885, B1 => n16947, B2 => 
                           n16884, ZN => n1545);
   U789 : OAI22_X1 port map( A1 => n18694, A2 => n16885, B1 => n16948, B2 => 
                           n16883, ZN => n1544);
   U790 : OAI22_X1 port map( A1 => n19207, A2 => n16885, B1 => n16949, B2 => 
                           n16884, ZN => n1543);
   U791 : OAI22_X1 port map( A1 => n18949, A2 => n16885, B1 => n16950, B2 => 
                           n16883, ZN => n1542);
   U792 : OAI22_X1 port map( A1 => n18695, A2 => n16885, B1 => n16951, B2 => 
                           n16883, ZN => n1541);
   U793 : OAI22_X1 port map( A1 => n18696, A2 => n16885, B1 => n16952, B2 => 
                           n16883, ZN => n1540);
   U794 : OAI22_X1 port map( A1 => n19208, A2 => n16885, B1 => n16953, B2 => 
                           n16883, ZN => n1539);
   U795 : OAI22_X1 port map( A1 => n19456, A2 => n16885, B1 => n16954, B2 => 
                           n16883, ZN => n1538);
   U796 : OAI22_X1 port map( A1 => n18950, A2 => n16885, B1 => n16955, B2 => 
                           n16883, ZN => n1537);
   U797 : OAI22_X1 port map( A1 => n19457, A2 => n16885, B1 => n16957, B2 => 
                           n16883, ZN => n1536);
   U798 : OAI22_X1 port map( A1 => n18951, A2 => n16885, B1 => n16958, B2 => 
                           n16884, ZN => n1535);
   U799 : OAI22_X1 port map( A1 => n19458, A2 => n16885, B1 => n16959, B2 => 
                           n16884, ZN => n1534);
   U800 : OAI22_X1 port map( A1 => n19459, A2 => n16885, B1 => n16960, B2 => 
                           n16884, ZN => n1533);
   U801 : OAI22_X1 port map( A1 => n19209, A2 => n16885, B1 => n16961, B2 => 
                           n16884, ZN => n1532);
   U802 : OAI22_X1 port map( A1 => n18952, A2 => n16885, B1 => n16962, B2 => 
                           n16884, ZN => n1531);
   U803 : OAI22_X1 port map( A1 => n19460, A2 => n16885, B1 => n16963, B2 => 
                           n16884, ZN => n1530);
   U804 : OAI22_X1 port map( A1 => n18697, A2 => n16885, B1 => n16964, B2 => 
                           n16884, ZN => n1529);
   U805 : OAI22_X1 port map( A1 => n19210, A2 => n16885, B1 => n16965, B2 => 
                           n16884, ZN => n1528);
   U806 : OAI22_X1 port map( A1 => n18698, A2 => n16885, B1 => n16967, B2 => 
                           n16884, ZN => n1527);
   U807 : NAND2_X1 port map( A1 => n16919, A2 => n16895, ZN => n16886);
   U808 : CLKBUF_X1 port map( A => n16886, Z => n16887);
   U809 : OAI22_X1 port map( A1 => n18789, A2 => n16888, B1 => n16896, B2 => 
                           n16887, ZN => n1526);
   U810 : OAI22_X1 port map( A1 => n19461, A2 => n16888, B1 => n16935, B2 => 
                           n16886, ZN => n1525);
   U811 : OAI22_X1 port map( A1 => n18699, A2 => n16888, B1 => n16936, B2 => 
                           n16887, ZN => n1524);
   U812 : OAI22_X1 port map( A1 => n19462, A2 => n16888, B1 => n16937, B2 => 
                           n16886, ZN => n1523);
   U813 : OAI22_X1 port map( A1 => n19463, A2 => n16888, B1 => n16938, B2 => 
                           n16887, ZN => n1522);
   U814 : OAI22_X1 port map( A1 => n18700, A2 => n16888, B1 => n16939, B2 => 
                           n16886, ZN => n1521);
   U815 : OAI22_X1 port map( A1 => n18953, A2 => n16888, B1 => n16940, B2 => 
                           n16887, ZN => n1520);
   U816 : OAI22_X1 port map( A1 => n18701, A2 => n16888, B1 => n16941, B2 => 
                           n16886, ZN => n1519);
   U817 : OAI22_X1 port map( A1 => n18954, A2 => n16888, B1 => n16942, B2 => 
                           n16887, ZN => n1518);
   U818 : OAI22_X1 port map( A1 => n18702, A2 => n16888, B1 => n16943, B2 => 
                           n16886, ZN => n1517);
   U819 : OAI22_X1 port map( A1 => n19464, A2 => n16888, B1 => n16944, B2 => 
                           n16886, ZN => n1516);
   U820 : OAI22_X1 port map( A1 => n18955, A2 => n16888, B1 => n16945, B2 => 
                           n16887, ZN => n1515);
   U821 : OAI22_X1 port map( A1 => n19211, A2 => n16888, B1 => n16946, B2 => 
                           n16886, ZN => n1514);
   U822 : OAI22_X1 port map( A1 => n19212, A2 => n16888, B1 => n16947, B2 => 
                           n16887, ZN => n1513);
   U823 : OAI22_X1 port map( A1 => n19213, A2 => n16888, B1 => n16948, B2 => 
                           n16886, ZN => n1512);
   U824 : OAI22_X1 port map( A1 => n19465, A2 => n16888, B1 => n16949, B2 => 
                           n16887, ZN => n1511);
   U825 : OAI22_X1 port map( A1 => n19214, A2 => n16888, B1 => n16950, B2 => 
                           n16886, ZN => n1510);
   U826 : OAI22_X1 port map( A1 => n19215, A2 => n16888, B1 => n16951, B2 => 
                           n16886, ZN => n1509);
   U827 : OAI22_X1 port map( A1 => n19216, A2 => n16888, B1 => n16952, B2 => 
                           n16886, ZN => n1508);
   U828 : OAI22_X1 port map( A1 => n19466, A2 => n16888, B1 => n16953, B2 => 
                           n16886, ZN => n1507);
   U829 : OAI22_X1 port map( A1 => n19217, A2 => n16888, B1 => n16954, B2 => 
                           n16886, ZN => n1506);
   U830 : OAI22_X1 port map( A1 => n19467, A2 => n16888, B1 => n16955, B2 => 
                           n16886, ZN => n1505);
   U831 : OAI22_X1 port map( A1 => n18956, A2 => n16888, B1 => n16957, B2 => 
                           n16886, ZN => n1504);
   U832 : OAI22_X1 port map( A1 => n18703, A2 => n16888, B1 => n16958, B2 => 
                           n16887, ZN => n1503);
   U833 : OAI22_X1 port map( A1 => n19218, A2 => n16888, B1 => n16959, B2 => 
                           n16887, ZN => n1502);
   U834 : OAI22_X1 port map( A1 => n19219, A2 => n16888, B1 => n16960, B2 => 
                           n16887, ZN => n1501);
   U835 : OAI22_X1 port map( A1 => n19468, A2 => n16888, B1 => n16961, B2 => 
                           n16887, ZN => n1500);
   U836 : OAI22_X1 port map( A1 => n19220, A2 => n16888, B1 => n16962, B2 => 
                           n16887, ZN => n1499);
   U837 : OAI22_X1 port map( A1 => n18704, A2 => n16888, B1 => n16963, B2 => 
                           n16887, ZN => n1498);
   U838 : OAI22_X1 port map( A1 => n19469, A2 => n16888, B1 => n16964, B2 => 
                           n16887, ZN => n1497);
   U839 : OAI22_X1 port map( A1 => n19221, A2 => n16888, B1 => n16965, B2 => 
                           n16887, ZN => n1496);
   U840 : OAI22_X1 port map( A1 => n19222, A2 => n16888, B1 => n16967, B2 => 
                           n16887, ZN => n1495);
   U841 : NAND2_X1 port map( A1 => n16923, A2 => n16895, ZN => n16889);
   U842 : CLKBUF_X1 port map( A => n16889, Z => n16890);
   U843 : OAI22_X1 port map( A1 => n18790, A2 => n16891, B1 => n16896, B2 => 
                           n16890, ZN => n1494);
   U844 : OAI22_X1 port map( A1 => n19223, A2 => n16891, B1 => n16935, B2 => 
                           n16889, ZN => n1493);
   U845 : OAI22_X1 port map( A1 => n19470, A2 => n16891, B1 => n16936, B2 => 
                           n16890, ZN => n1492);
   U846 : OAI22_X1 port map( A1 => n19471, A2 => n16891, B1 => n16937, B2 => 
                           n16889, ZN => n1491);
   U847 : OAI22_X1 port map( A1 => n19224, A2 => n16891, B1 => n16938, B2 => 
                           n16890, ZN => n1490);
   U848 : OAI22_X1 port map( A1 => n19225, A2 => n16891, B1 => n16939, B2 => 
                           n16889, ZN => n1489);
   U849 : OAI22_X1 port map( A1 => n19226, A2 => n16891, B1 => n16940, B2 => 
                           n16890, ZN => n1488);
   U850 : OAI22_X1 port map( A1 => n19227, A2 => n16891, B1 => n16941, B2 => 
                           n16889, ZN => n1487);
   U851 : OAI22_X1 port map( A1 => n19472, A2 => n16891, B1 => n16942, B2 => 
                           n16890, ZN => n1486);
   U852 : OAI22_X1 port map( A1 => n19473, A2 => n16891, B1 => n16943, B2 => 
                           n16889, ZN => n1485);
   U853 : OAI22_X1 port map( A1 => n19474, A2 => n16891, B1 => n16944, B2 => 
                           n16889, ZN => n1484);
   U854 : OAI22_X1 port map( A1 => n19475, A2 => n16891, B1 => n16945, B2 => 
                           n16890, ZN => n1483);
   U855 : OAI22_X1 port map( A1 => n18957, A2 => n16891, B1 => n16946, B2 => 
                           n16889, ZN => n1482);
   U856 : OAI22_X1 port map( A1 => n19476, A2 => n16891, B1 => n16947, B2 => 
                           n16890, ZN => n1481);
   U857 : OAI22_X1 port map( A1 => n19477, A2 => n16891, B1 => n16948, B2 => 
                           n16889, ZN => n1480);
   U858 : OAI22_X1 port map( A1 => n19478, A2 => n16891, B1 => n16949, B2 => 
                           n16890, ZN => n1479);
   U859 : OAI22_X1 port map( A1 => n19479, A2 => n16891, B1 => n16950, B2 => 
                           n16889, ZN => n1478);
   U860 : OAI22_X1 port map( A1 => n19480, A2 => n16891, B1 => n16951, B2 => 
                           n16889, ZN => n1477);
   U861 : OAI22_X1 port map( A1 => n19228, A2 => n16891, B1 => n16952, B2 => 
                           n16889, ZN => n1476);
   U862 : OAI22_X1 port map( A1 => n19481, A2 => n16891, B1 => n16953, B2 => 
                           n16889, ZN => n1475);
   U863 : OAI22_X1 port map( A1 => n19229, A2 => n16891, B1 => n16954, B2 => 
                           n16889, ZN => n1474);
   U864 : OAI22_X1 port map( A1 => n19230, A2 => n16891, B1 => n16955, B2 => 
                           n16889, ZN => n1473);
   U865 : OAI22_X1 port map( A1 => n19231, A2 => n16891, B1 => n16957, B2 => 
                           n16889, ZN => n1472);
   U866 : OAI22_X1 port map( A1 => n19482, A2 => n16891, B1 => n16958, B2 => 
                           n16890, ZN => n1471);
   U867 : OAI22_X1 port map( A1 => n19232, A2 => n16891, B1 => n16959, B2 => 
                           n16890, ZN => n1470);
   U868 : OAI22_X1 port map( A1 => n18705, A2 => n16891, B1 => n16960, B2 => 
                           n16890, ZN => n1469);
   U869 : OAI22_X1 port map( A1 => n19483, A2 => n16891, B1 => n16961, B2 => 
                           n16890, ZN => n1468);
   U870 : OAI22_X1 port map( A1 => n19233, A2 => n16891, B1 => n16962, B2 => 
                           n16890, ZN => n1467);
   U871 : OAI22_X1 port map( A1 => n19234, A2 => n16891, B1 => n16963, B2 => 
                           n16890, ZN => n1466);
   U872 : OAI22_X1 port map( A1 => n19484, A2 => n16891, B1 => n16964, B2 => 
                           n16890, ZN => n1465);
   U873 : OAI22_X1 port map( A1 => n18706, A2 => n16891, B1 => n16965, B2 => 
                           n16890, ZN => n1464);
   U874 : OAI22_X1 port map( A1 => n19485, A2 => n16891, B1 => n16967, B2 => 
                           n16890, ZN => n1463);
   U875 : NAND2_X1 port map( A1 => n16928, A2 => n16895, ZN => n16892);
   U876 : CLKBUF_X1 port map( A => n16892, Z => n16893);
   U877 : OAI22_X1 port map( A1 => n19047, A2 => n16894, B1 => n16896, B2 => 
                           n16893, ZN => n1462);
   U878 : OAI22_X1 port map( A1 => n19486, A2 => n16894, B1 => n16935, B2 => 
                           n16892, ZN => n1461);
   U879 : OAI22_X1 port map( A1 => n19487, A2 => n16894, B1 => n16936, B2 => 
                           n16893, ZN => n1460);
   U880 : OAI22_X1 port map( A1 => n19235, A2 => n16894, B1 => n16937, B2 => 
                           n16892, ZN => n1459);
   U881 : OAI22_X1 port map( A1 => n19236, A2 => n16894, B1 => n16938, B2 => 
                           n16893, ZN => n1458);
   U882 : OAI22_X1 port map( A1 => n19488, A2 => n16894, B1 => n16939, B2 => 
                           n16892, ZN => n1457);
   U883 : OAI22_X1 port map( A1 => n19237, A2 => n16894, B1 => n16940, B2 => 
                           n16893, ZN => n1456);
   U884 : OAI22_X1 port map( A1 => n19489, A2 => n16894, B1 => n16941, B2 => 
                           n16892, ZN => n1455);
   U885 : OAI22_X1 port map( A1 => n19490, A2 => n16894, B1 => n16942, B2 => 
                           n16893, ZN => n1454);
   U886 : OAI22_X1 port map( A1 => n19491, A2 => n16894, B1 => n16943, B2 => 
                           n16892, ZN => n1453);
   U887 : OAI22_X1 port map( A1 => n19492, A2 => n16894, B1 => n16944, B2 => 
                           n16892, ZN => n1452);
   U888 : OAI22_X1 port map( A1 => n19493, A2 => n16894, B1 => n16945, B2 => 
                           n16893, ZN => n1451);
   U889 : OAI22_X1 port map( A1 => n19494, A2 => n16894, B1 => n16946, B2 => 
                           n16892, ZN => n1450);
   U890 : OAI22_X1 port map( A1 => n19238, A2 => n16894, B1 => n16947, B2 => 
                           n16893, ZN => n1449);
   U891 : OAI22_X1 port map( A1 => n19239, A2 => n16894, B1 => n16948, B2 => 
                           n16892, ZN => n1448);
   U892 : OAI22_X1 port map( A1 => n19240, A2 => n16894, B1 => n16949, B2 => 
                           n16893, ZN => n1447);
   U893 : OAI22_X1 port map( A1 => n19495, A2 => n16894, B1 => n16950, B2 => 
                           n16892, ZN => n1446);
   U894 : OAI22_X1 port map( A1 => n19496, A2 => n16894, B1 => n16951, B2 => 
                           n16892, ZN => n1445);
   U895 : OAI22_X1 port map( A1 => n19497, A2 => n16894, B1 => n16952, B2 => 
                           n16892, ZN => n1444);
   U896 : OAI22_X1 port map( A1 => n19241, A2 => n16894, B1 => n16953, B2 => 
                           n16892, ZN => n1443);
   U897 : OAI22_X1 port map( A1 => n19242, A2 => n16894, B1 => n16954, B2 => 
                           n16892, ZN => n1442);
   U898 : OAI22_X1 port map( A1 => n19243, A2 => n16894, B1 => n16955, B2 => 
                           n16892, ZN => n1441);
   U899 : OAI22_X1 port map( A1 => n19244, A2 => n16894, B1 => n16957, B2 => 
                           n16892, ZN => n1440);
   U900 : OAI22_X1 port map( A1 => n19245, A2 => n16894, B1 => n16958, B2 => 
                           n16893, ZN => n1439);
   U901 : OAI22_X1 port map( A1 => n19498, A2 => n16894, B1 => n16959, B2 => 
                           n16893, ZN => n1438);
   U902 : OAI22_X1 port map( A1 => n19499, A2 => n16894, B1 => n16960, B2 => 
                           n16893, ZN => n1437);
   U903 : OAI22_X1 port map( A1 => n19246, A2 => n16894, B1 => n16961, B2 => 
                           n16893, ZN => n1436);
   U904 : OAI22_X1 port map( A1 => n19500, A2 => n16894, B1 => n16962, B2 => 
                           n16893, ZN => n1435);
   U905 : OAI22_X1 port map( A1 => n19501, A2 => n16894, B1 => n16963, B2 => 
                           n16893, ZN => n1434);
   U906 : OAI22_X1 port map( A1 => n19502, A2 => n16894, B1 => n16964, B2 => 
                           n16893, ZN => n1433);
   U907 : OAI22_X1 port map( A1 => n19247, A2 => n16894, B1 => n16965, B2 => 
                           n16893, ZN => n1432);
   U908 : OAI22_X1 port map( A1 => n19503, A2 => n16894, B1 => n16967, B2 => 
                           n16893, ZN => n1431);
   U909 : NAND2_X1 port map( A1 => n16933, A2 => n16895, ZN => n16897);
   U910 : CLKBUF_X1 port map( A => n16897, Z => n16898);
   U911 : OAI22_X1 port map( A1 => n19048, A2 => n16899, B1 => n16896, B2 => 
                           n16898, ZN => n1430);
   U912 : OAI22_X1 port map( A1 => n19248, A2 => n16899, B1 => n16935, B2 => 
                           n16897, ZN => n1429);
   U913 : OAI22_X1 port map( A1 => n18958, A2 => n16899, B1 => n16936, B2 => 
                           n16898, ZN => n1428);
   U914 : OAI22_X1 port map( A1 => n18707, A2 => n16899, B1 => n16937, B2 => 
                           n16897, ZN => n1427);
   U915 : OAI22_X1 port map( A1 => n18959, A2 => n16899, B1 => n16938, B2 => 
                           n16898, ZN => n1426);
   U916 : OAI22_X1 port map( A1 => n18960, A2 => n16899, B1 => n16939, B2 => 
                           n16897, ZN => n1425);
   U917 : OAI22_X1 port map( A1 => n18961, A2 => n16899, B1 => n16940, B2 => 
                           n16898, ZN => n1424);
   U918 : OAI22_X1 port map( A1 => n18962, A2 => n16899, B1 => n16941, B2 => 
                           n16897, ZN => n1423);
   U919 : OAI22_X1 port map( A1 => n19504, A2 => n16899, B1 => n16942, B2 => 
                           n16898, ZN => n1422);
   U920 : OAI22_X1 port map( A1 => n18963, A2 => n16899, B1 => n16943, B2 => 
                           n16897, ZN => n1421);
   U921 : OAI22_X1 port map( A1 => n18708, A2 => n16899, B1 => n16944, B2 => 
                           n16897, ZN => n1420);
   U922 : OAI22_X1 port map( A1 => n18964, A2 => n16899, B1 => n16945, B2 => 
                           n16898, ZN => n1419);
   U923 : OAI22_X1 port map( A1 => n18965, A2 => n16899, B1 => n16946, B2 => 
                           n16897, ZN => n1418);
   U924 : OAI22_X1 port map( A1 => n19505, A2 => n16899, B1 => n16947, B2 => 
                           n16898, ZN => n1417);
   U925 : OAI22_X1 port map( A1 => n19249, A2 => n16899, B1 => n16948, B2 => 
                           n16897, ZN => n1416);
   U926 : OAI22_X1 port map( A1 => n19506, A2 => n16899, B1 => n16949, B2 => 
                           n16898, ZN => n1415);
   U927 : OAI22_X1 port map( A1 => n18966, A2 => n16899, B1 => n16950, B2 => 
                           n16897, ZN => n1414);
   U928 : OAI22_X1 port map( A1 => n18709, A2 => n16899, B1 => n16951, B2 => 
                           n16897, ZN => n1413);
   U929 : OAI22_X1 port map( A1 => n19507, A2 => n16899, B1 => n16952, B2 => 
                           n16897, ZN => n1412);
   U930 : OAI22_X1 port map( A1 => n18710, A2 => n16899, B1 => n16953, B2 => 
                           n16897, ZN => n1411);
   U931 : OAI22_X1 port map( A1 => n18967, A2 => n16899, B1 => n16954, B2 => 
                           n16897, ZN => n1410);
   U932 : OAI22_X1 port map( A1 => n18711, A2 => n16899, B1 => n16955, B2 => 
                           n16897, ZN => n1409);
   U933 : OAI22_X1 port map( A1 => n18968, A2 => n16899, B1 => n16957, B2 => 
                           n16897, ZN => n1408);
   U934 : OAI22_X1 port map( A1 => n18969, A2 => n16899, B1 => n16958, B2 => 
                           n16898, ZN => n1407);
   U935 : OAI22_X1 port map( A1 => n18712, A2 => n16899, B1 => n16959, B2 => 
                           n16898, ZN => n1406);
   U936 : OAI22_X1 port map( A1 => n18970, A2 => n16899, B1 => n16960, B2 => 
                           n16898, ZN => n1405);
   U937 : OAI22_X1 port map( A1 => n18971, A2 => n16899, B1 => n16961, B2 => 
                           n16898, ZN => n1404);
   U938 : OAI22_X1 port map( A1 => n18713, A2 => n16899, B1 => n16962, B2 => 
                           n16898, ZN => n1403);
   U939 : OAI22_X1 port map( A1 => n19508, A2 => n16899, B1 => n16963, B2 => 
                           n16898, ZN => n1402);
   U940 : OAI22_X1 port map( A1 => n18972, A2 => n16899, B1 => n16964, B2 => 
                           n16898, ZN => n1401);
   U941 : OAI22_X1 port map( A1 => n18973, A2 => n16899, B1 => n16965, B2 => 
                           n16898, ZN => n1400);
   U942 : OAI22_X1 port map( A1 => n18714, A2 => n16899, B1 => n16967, B2 => 
                           n16898, ZN => n1399);
   U943 : NOR2_X1 port map( A1 => n16901, A2 => n16900, ZN => n16932);
   U944 : NAND2_X1 port map( A1 => n16902, A2 => n16932, ZN => n16903);
   U945 : CLKBUF_X1 port map( A => n16903, Z => n16904);
   U946 : OAI22_X1 port map( A1 => n18791, A2 => n16905, B1 => n16934, B2 => 
                           n16904, ZN => n1398);
   U947 : OAI22_X1 port map( A1 => n18974, A2 => n16905, B1 => n16935, B2 => 
                           n16903, ZN => n1397);
   U948 : OAI22_X1 port map( A1 => n18715, A2 => n16905, B1 => n16936, B2 => 
                           n16904, ZN => n1396);
   U949 : OAI22_X1 port map( A1 => n18975, A2 => n16905, B1 => n16937, B2 => 
                           n16903, ZN => n1395);
   U950 : OAI22_X1 port map( A1 => n18976, A2 => n16905, B1 => n16938, B2 => 
                           n16904, ZN => n1394);
   U951 : OAI22_X1 port map( A1 => n18977, A2 => n16905, B1 => n16939, B2 => 
                           n16903, ZN => n1393);
   U952 : OAI22_X1 port map( A1 => n18716, A2 => n16905, B1 => n16940, B2 => 
                           n16904, ZN => n1392);
   U953 : OAI22_X1 port map( A1 => n18717, A2 => n16905, B1 => n16941, B2 => 
                           n16903, ZN => n1391);
   U954 : OAI22_X1 port map( A1 => n18718, A2 => n16905, B1 => n16942, B2 => 
                           n16904, ZN => n1390);
   U955 : OAI22_X1 port map( A1 => n18978, A2 => n16905, B1 => n16943, B2 => 
                           n16903, ZN => n1389);
   U956 : OAI22_X1 port map( A1 => n18979, A2 => n16905, B1 => n16944, B2 => 
                           n16903, ZN => n1388);
   U957 : OAI22_X1 port map( A1 => n18980, A2 => n16905, B1 => n16945, B2 => 
                           n16904, ZN => n1387);
   U958 : OAI22_X1 port map( A1 => n18981, A2 => n16905, B1 => n16946, B2 => 
                           n16903, ZN => n1386);
   U959 : OAI22_X1 port map( A1 => n18982, A2 => n16905, B1 => n16947, B2 => 
                           n16904, ZN => n1385);
   U960 : OAI22_X1 port map( A1 => n18719, A2 => n16905, B1 => n16948, B2 => 
                           n16903, ZN => n1384);
   U961 : OAI22_X1 port map( A1 => n18983, A2 => n16905, B1 => n16949, B2 => 
                           n16904, ZN => n1383);
   U962 : OAI22_X1 port map( A1 => n18984, A2 => n16905, B1 => n16950, B2 => 
                           n16903, ZN => n1382);
   U963 : OAI22_X1 port map( A1 => n18985, A2 => n16905, B1 => n16951, B2 => 
                           n16903, ZN => n1381);
   U964 : OAI22_X1 port map( A1 => n18720, A2 => n16905, B1 => n16952, B2 => 
                           n16903, ZN => n1380);
   U965 : OAI22_X1 port map( A1 => n18986, A2 => n16905, B1 => n16953, B2 => 
                           n16903, ZN => n1379);
   U966 : OAI22_X1 port map( A1 => n18987, A2 => n16905, B1 => n16954, B2 => 
                           n16903, ZN => n1378);
   U967 : OAI22_X1 port map( A1 => n19250, A2 => n16905, B1 => n16955, B2 => 
                           n16903, ZN => n1377);
   U968 : OAI22_X1 port map( A1 => n18721, A2 => n16905, B1 => n16957, B2 => 
                           n16903, ZN => n1376);
   U969 : OAI22_X1 port map( A1 => n18722, A2 => n16905, B1 => n16958, B2 => 
                           n16904, ZN => n1375);
   U970 : OAI22_X1 port map( A1 => n18723, A2 => n16905, B1 => n16959, B2 => 
                           n16904, ZN => n1374);
   U971 : OAI22_X1 port map( A1 => n19509, A2 => n16905, B1 => n16960, B2 => 
                           n16904, ZN => n1373);
   U972 : OAI22_X1 port map( A1 => n18724, A2 => n16905, B1 => n16961, B2 => 
                           n16904, ZN => n1372);
   U973 : OAI22_X1 port map( A1 => n18725, A2 => n16905, B1 => n16962, B2 => 
                           n16904, ZN => n1371);
   U974 : OAI22_X1 port map( A1 => n18726, A2 => n16905, B1 => n16963, B2 => 
                           n16904, ZN => n1370);
   U975 : OAI22_X1 port map( A1 => n18727, A2 => n16905, B1 => n16964, B2 => 
                           n16904, ZN => n1369);
   U976 : OAI22_X1 port map( A1 => n18728, A2 => n16905, B1 => n16965, B2 => 
                           n16904, ZN => n1368);
   U977 : OAI22_X1 port map( A1 => n18988, A2 => n16905, B1 => n16967, B2 => 
                           n16904, ZN => n1367);
   U978 : NAND2_X1 port map( A1 => n16906, A2 => n16932, ZN => n16907);
   U979 : CLKBUF_X1 port map( A => n16910, Z => n16908);
   U980 : CLKBUF_X1 port map( A => n16907, Z => n16909);
   U981 : OAI22_X1 port map( A1 => n18792, A2 => n16908, B1 => n16934, B2 => 
                           n16909, ZN => n1366);
   U982 : OAI22_X1 port map( A1 => n18729, A2 => n16910, B1 => n16935, B2 => 
                           n16907, ZN => n1365);
   U983 : OAI22_X1 port map( A1 => n19251, A2 => n16908, B1 => n16936, B2 => 
                           n16909, ZN => n1364);
   U984 : OAI22_X1 port map( A1 => n19252, A2 => n16910, B1 => n16937, B2 => 
                           n16907, ZN => n1363);
   U985 : OAI22_X1 port map( A1 => n19253, A2 => n16908, B1 => n16938, B2 => 
                           n16909, ZN => n1362);
   U986 : OAI22_X1 port map( A1 => n19510, A2 => n16910, B1 => n16939, B2 => 
                           n16907, ZN => n1361);
   U987 : OAI22_X1 port map( A1 => n19254, A2 => n16908, B1 => n16940, B2 => 
                           n16909, ZN => n1360);
   U988 : OAI22_X1 port map( A1 => n19511, A2 => n16910, B1 => n16941, B2 => 
                           n16907, ZN => n1359);
   U989 : OAI22_X1 port map( A1 => n19255, A2 => n16908, B1 => n16942, B2 => 
                           n16909, ZN => n1358);
   U990 : OAI22_X1 port map( A1 => n19256, A2 => n16910, B1 => n16943, B2 => 
                           n16907, ZN => n1357);
   U991 : OAI22_X1 port map( A1 => n18989, A2 => n16910, B1 => n16944, B2 => 
                           n16907, ZN => n1356);
   U992 : OAI22_X1 port map( A1 => n19257, A2 => n16910, B1 => n16945, B2 => 
                           n16909, ZN => n1355);
   U993 : OAI22_X1 port map( A1 => n19512, A2 => n16908, B1 => n16946, B2 => 
                           n16907, ZN => n1354);
   U994 : OAI22_X1 port map( A1 => n18730, A2 => n16908, B1 => n16947, B2 => 
                           n16909, ZN => n1353);
   U995 : OAI22_X1 port map( A1 => n19258, A2 => n16908, B1 => n16948, B2 => 
                           n16907, ZN => n1352);
   U996 : OAI22_X1 port map( A1 => n18731, A2 => n16908, B1 => n16949, B2 => 
                           n16909, ZN => n1351);
   U997 : OAI22_X1 port map( A1 => n19259, A2 => n16908, B1 => n16950, B2 => 
                           n16907, ZN => n1350);
   U998 : OAI22_X1 port map( A1 => n19260, A2 => n16908, B1 => n16951, B2 => 
                           n16907, ZN => n1349);
   U999 : OAI22_X1 port map( A1 => n19513, A2 => n16908, B1 => n16952, B2 => 
                           n16907, ZN => n1348);
   U1000 : OAI22_X1 port map( A1 => n18990, A2 => n16908, B1 => n16953, B2 => 
                           n16907, ZN => n1347);
   U1001 : OAI22_X1 port map( A1 => n18991, A2 => n16908, B1 => n16954, B2 => 
                           n16907, ZN => n1346);
   U1002 : OAI22_X1 port map( A1 => n18992, A2 => n16908, B1 => n16955, B2 => 
                           n16907, ZN => n1345);
   U1003 : OAI22_X1 port map( A1 => n19261, A2 => n16908, B1 => n16957, B2 => 
                           n16907, ZN => n1344);
   U1004 : OAI22_X1 port map( A1 => n19514, A2 => n16908, B1 => n16958, B2 => 
                           n16909, ZN => n1343);
   U1005 : OAI22_X1 port map( A1 => n19262, A2 => n16910, B1 => n16959, B2 => 
                           n16909, ZN => n1342);
   U1006 : OAI22_X1 port map( A1 => n19263, A2 => n16910, B1 => n16960, B2 => 
                           n16909, ZN => n1341);
   U1007 : OAI22_X1 port map( A1 => n19515, A2 => n16910, B1 => n16961, B2 => 
                           n16909, ZN => n1340);
   U1008 : OAI22_X1 port map( A1 => n19516, A2 => n16910, B1 => n16962, B2 => 
                           n16909, ZN => n1339);
   U1009 : OAI22_X1 port map( A1 => n19264, A2 => n16910, B1 => n16963, B2 => 
                           n16909, ZN => n1338);
   U1010 : OAI22_X1 port map( A1 => n19265, A2 => n16910, B1 => n16964, B2 => 
                           n16909, ZN => n1337);
   U1011 : OAI22_X1 port map( A1 => n19517, A2 => n16910, B1 => n16965, B2 => 
                           n16909, ZN => n1336);
   U1012 : OAI22_X1 port map( A1 => n19518, A2 => n16910, B1 => n16967, B2 => 
                           n16909, ZN => n1335);
   U1013 : NAND2_X1 port map( A1 => n16911, A2 => n16932, ZN => n16912);
   U1014 : CLKBUF_X1 port map( A => n16912, Z => n16913);
   U1015 : OAI22_X1 port map( A1 => n18793, A2 => n16914, B1 => n16934, B2 => 
                           n16913, ZN => n1334);
   U1016 : OAI22_X1 port map( A1 => n18993, A2 => n16914, B1 => n16935, B2 => 
                           n16912, ZN => n1333);
   U1017 : OAI22_X1 port map( A1 => n19519, A2 => n16914, B1 => n16936, B2 => 
                           n16913, ZN => n1332);
   U1018 : OAI22_X1 port map( A1 => n19520, A2 => n16914, B1 => n16937, B2 => 
                           n16912, ZN => n1331);
   U1019 : OAI22_X1 port map( A1 => n18994, A2 => n16914, B1 => n16938, B2 => 
                           n16913, ZN => n1330);
   U1020 : OAI22_X1 port map( A1 => n19521, A2 => n16914, B1 => n16939, B2 => 
                           n16912, ZN => n1329);
   U1021 : OAI22_X1 port map( A1 => n19522, A2 => n16914, B1 => n16940, B2 => 
                           n16913, ZN => n1328);
   U1022 : OAI22_X1 port map( A1 => n19523, A2 => n16914, B1 => n16941, B2 => 
                           n16912, ZN => n1327);
   U1023 : OAI22_X1 port map( A1 => n19266, A2 => n16914, B1 => n16942, B2 => 
                           n16913, ZN => n1326);
   U1024 : OAI22_X1 port map( A1 => n19267, A2 => n16914, B1 => n16943, B2 => 
                           n16912, ZN => n1325);
   U1025 : OAI22_X1 port map( A1 => n18732, A2 => n16914, B1 => n16944, B2 => 
                           n16912, ZN => n1324);
   U1026 : OAI22_X1 port map( A1 => n18733, A2 => n16914, B1 => n16945, B2 => 
                           n16913, ZN => n1323);
   U1027 : OAI22_X1 port map( A1 => n19268, A2 => n16914, B1 => n16946, B2 => 
                           n16912, ZN => n1322);
   U1028 : OAI22_X1 port map( A1 => n19269, A2 => n16914, B1 => n16947, B2 => 
                           n16913, ZN => n1321);
   U1029 : OAI22_X1 port map( A1 => n18995, A2 => n16914, B1 => n16948, B2 => 
                           n16912, ZN => n1320);
   U1030 : OAI22_X1 port map( A1 => n18734, A2 => n16914, B1 => n16949, B2 => 
                           n16913, ZN => n1319);
   U1031 : OAI22_X1 port map( A1 => n19270, A2 => n16914, B1 => n16950, B2 => 
                           n16912, ZN => n1318);
   U1032 : OAI22_X1 port map( A1 => n18735, A2 => n16914, B1 => n16951, B2 => 
                           n16912, ZN => n1317);
   U1033 : OAI22_X1 port map( A1 => n18996, A2 => n16914, B1 => n16952, B2 => 
                           n16912, ZN => n1316);
   U1034 : OAI22_X1 port map( A1 => n19271, A2 => n16914, B1 => n16953, B2 => 
                           n16912, ZN => n1315);
   U1035 : OAI22_X1 port map( A1 => n19524, A2 => n16914, B1 => n16954, B2 => 
                           n16912, ZN => n1314);
   U1036 : OAI22_X1 port map( A1 => n19272, A2 => n16914, B1 => n16955, B2 => 
                           n16912, ZN => n1313);
   U1037 : OAI22_X1 port map( A1 => n19525, A2 => n16914, B1 => n16957, B2 => 
                           n16912, ZN => n1312);
   U1038 : OAI22_X1 port map( A1 => n19273, A2 => n16914, B1 => n16958, B2 => 
                           n16913, ZN => n1311);
   U1039 : OAI22_X1 port map( A1 => n18736, A2 => n16914, B1 => n16959, B2 => 
                           n16913, ZN => n1310);
   U1040 : OAI22_X1 port map( A1 => n18737, A2 => n16914, B1 => n16960, B2 => 
                           n16913, ZN => n1309);
   U1041 : OAI22_X1 port map( A1 => n18997, A2 => n16914, B1 => n16961, B2 => 
                           n16913, ZN => n1308);
   U1042 : OAI22_X1 port map( A1 => n19526, A2 => n16914, B1 => n16962, B2 => 
                           n16913, ZN => n1307);
   U1043 : OAI22_X1 port map( A1 => n18738, A2 => n16914, B1 => n16963, B2 => 
                           n16913, ZN => n1306);
   U1044 : OAI22_X1 port map( A1 => n19274, A2 => n16914, B1 => n16964, B2 => 
                           n16913, ZN => n1305);
   U1045 : OAI22_X1 port map( A1 => n18998, A2 => n16914, B1 => n16965, B2 => 
                           n16913, ZN => n1304);
   U1046 : OAI22_X1 port map( A1 => n19527, A2 => n16914, B1 => n16967, B2 => 
                           n16913, ZN => n1303);
   U1047 : NAND2_X1 port map( A1 => n16915, A2 => n16932, ZN => n16916);
   U1048 : CLKBUF_X1 port map( A => n16916, Z => n16917);
   U1049 : OAI22_X1 port map( A1 => n19049, A2 => n16918, B1 => n16934, B2 => 
                           n16917, ZN => n1302);
   U1050 : OAI22_X1 port map( A1 => n19528, A2 => n16918, B1 => n16935, B2 => 
                           n16916, ZN => n1301);
   U1051 : OAI22_X1 port map( A1 => n19529, A2 => n16918, B1 => n16936, B2 => 
                           n16917, ZN => n1300);
   U1052 : OAI22_X1 port map( A1 => n19275, A2 => n16918, B1 => n16937, B2 => 
                           n16916, ZN => n1299);
   U1053 : OAI22_X1 port map( A1 => n19530, A2 => n16918, B1 => n16938, B2 => 
                           n16917, ZN => n1298);
   U1054 : OAI22_X1 port map( A1 => n19531, A2 => n16918, B1 => n16939, B2 => 
                           n16916, ZN => n1297);
   U1055 : OAI22_X1 port map( A1 => n19276, A2 => n16918, B1 => n16940, B2 => 
                           n16917, ZN => n1296);
   U1056 : OAI22_X1 port map( A1 => n18739, A2 => n16918, B1 => n16941, B2 => 
                           n16916, ZN => n1295);
   U1057 : OAI22_X1 port map( A1 => n19532, A2 => n16918, B1 => n16942, B2 => 
                           n16917, ZN => n1294);
   U1058 : OAI22_X1 port map( A1 => n19533, A2 => n16918, B1 => n16943, B2 => 
                           n16916, ZN => n1293);
   U1059 : OAI22_X1 port map( A1 => n19277, A2 => n16918, B1 => n16944, B2 => 
                           n16916, ZN => n1292);
   U1060 : OAI22_X1 port map( A1 => n19534, A2 => n16918, B1 => n16945, B2 => 
                           n16917, ZN => n1291);
   U1061 : OAI22_X1 port map( A1 => n19278, A2 => n16918, B1 => n16946, B2 => 
                           n16916, ZN => n1290);
   U1062 : OAI22_X1 port map( A1 => n18999, A2 => n16918, B1 => n16947, B2 => 
                           n16917, ZN => n1289);
   U1063 : OAI22_X1 port map( A1 => n19535, A2 => n16918, B1 => n16948, B2 => 
                           n16916, ZN => n1288);
   U1064 : OAI22_X1 port map( A1 => n19536, A2 => n16918, B1 => n16949, B2 => 
                           n16917, ZN => n1287);
   U1065 : OAI22_X1 port map( A1 => n18740, A2 => n16918, B1 => n16950, B2 => 
                           n16916, ZN => n1286);
   U1066 : OAI22_X1 port map( A1 => n19537, A2 => n16918, B1 => n16951, B2 => 
                           n16916, ZN => n1285);
   U1067 : OAI22_X1 port map( A1 => n18741, A2 => n16918, B1 => n16952, B2 => 
                           n16916, ZN => n1284);
   U1068 : OAI22_X1 port map( A1 => n19000, A2 => n16918, B1 => n16953, B2 => 
                           n16916, ZN => n1283);
   U1069 : OAI22_X1 port map( A1 => n19279, A2 => n16918, B1 => n16954, B2 => 
                           n16916, ZN => n1282);
   U1070 : OAI22_X1 port map( A1 => n18742, A2 => n16918, B1 => n16955, B2 => 
                           n16916, ZN => n1281);
   U1071 : OAI22_X1 port map( A1 => n19280, A2 => n16918, B1 => n16957, B2 => 
                           n16916, ZN => n1280);
   U1072 : OAI22_X1 port map( A1 => n19538, A2 => n16918, B1 => n16958, B2 => 
                           n16917, ZN => n1279);
   U1073 : OAI22_X1 port map( A1 => n19281, A2 => n16918, B1 => n16959, B2 => 
                           n16917, ZN => n1278);
   U1074 : OAI22_X1 port map( A1 => n19282, A2 => n16918, B1 => n16960, B2 => 
                           n16917, ZN => n1277);
   U1075 : OAI22_X1 port map( A1 => n19283, A2 => n16918, B1 => n16961, B2 => 
                           n16917, ZN => n1276);
   U1076 : OAI22_X1 port map( A1 => n19539, A2 => n16918, B1 => n16962, B2 => 
                           n16917, ZN => n1275);
   U1077 : OAI22_X1 port map( A1 => n18743, A2 => n16918, B1 => n16963, B2 => 
                           n16917, ZN => n1274);
   U1078 : OAI22_X1 port map( A1 => n19284, A2 => n16918, B1 => n16964, B2 => 
                           n16917, ZN => n1273);
   U1079 : OAI22_X1 port map( A1 => n19285, A2 => n16918, B1 => n16965, B2 => 
                           n16917, ZN => n1272);
   U1080 : OAI22_X1 port map( A1 => n19286, A2 => n16918, B1 => n16967, B2 => 
                           n16917, ZN => n1271);
   U1081 : NAND2_X1 port map( A1 => n16919, A2 => n16932, ZN => n16920);
   U1082 : CLKBUF_X1 port map( A => n16920, Z => n16921);
   U1083 : OAI22_X1 port map( A1 => n19050, A2 => n16922, B1 => n16934, B2 => 
                           n16921, ZN => n1270);
   U1084 : OAI22_X1 port map( A1 => n19540, A2 => n16922, B1 => n16935, B2 => 
                           n16920, ZN => n1269);
   U1085 : OAI22_X1 port map( A1 => n19541, A2 => n16922, B1 => n16936, B2 => 
                           n16921, ZN => n1268);
   U1086 : OAI22_X1 port map( A1 => n18744, A2 => n16922, B1 => n16937, B2 => 
                           n16920, ZN => n1267);
   U1087 : OAI22_X1 port map( A1 => n19287, A2 => n16922, B1 => n16938, B2 => 
                           n16921, ZN => n1266);
   U1088 : OAI22_X1 port map( A1 => n19288, A2 => n16922, B1 => n16939, B2 => 
                           n16920, ZN => n1265);
   U1089 : OAI22_X1 port map( A1 => n19289, A2 => n16922, B1 => n16940, B2 => 
                           n16921, ZN => n1264);
   U1090 : OAI22_X1 port map( A1 => n19290, A2 => n16922, B1 => n16941, B2 => 
                           n16920, ZN => n1263);
   U1091 : OAI22_X1 port map( A1 => n19291, A2 => n16922, B1 => n16942, B2 => 
                           n16921, ZN => n1262);
   U1092 : OAI22_X1 port map( A1 => n19292, A2 => n16922, B1 => n16943, B2 => 
                           n16920, ZN => n1261);
   U1093 : OAI22_X1 port map( A1 => n19293, A2 => n16922, B1 => n16944, B2 => 
                           n16920, ZN => n1260);
   U1094 : OAI22_X1 port map( A1 => n19294, A2 => n16922, B1 => n16945, B2 => 
                           n16921, ZN => n1259);
   U1095 : OAI22_X1 port map( A1 => n19295, A2 => n16922, B1 => n16946, B2 => 
                           n16920, ZN => n1258);
   U1096 : OAI22_X1 port map( A1 => n19296, A2 => n16922, B1 => n16947, B2 => 
                           n16921, ZN => n1257);
   U1097 : OAI22_X1 port map( A1 => n19542, A2 => n16922, B1 => n16948, B2 => 
                           n16920, ZN => n1256);
   U1098 : OAI22_X1 port map( A1 => n19297, A2 => n16922, B1 => n16949, B2 => 
                           n16921, ZN => n1255);
   U1099 : OAI22_X1 port map( A1 => n18745, A2 => n16922, B1 => n16950, B2 => 
                           n16920, ZN => n1254);
   U1100 : OAI22_X1 port map( A1 => n19001, A2 => n16922, B1 => n16951, B2 => 
                           n16920, ZN => n1253);
   U1101 : OAI22_X1 port map( A1 => n19002, A2 => n16922, B1 => n16952, B2 => 
                           n16920, ZN => n1252);
   U1102 : OAI22_X1 port map( A1 => n19543, A2 => n16922, B1 => n16953, B2 => 
                           n16920, ZN => n1251);
   U1103 : OAI22_X1 port map( A1 => n19544, A2 => n16922, B1 => n16954, B2 => 
                           n16920, ZN => n1250);
   U1104 : OAI22_X1 port map( A1 => n19545, A2 => n16922, B1 => n16955, B2 => 
                           n16920, ZN => n1249);
   U1105 : OAI22_X1 port map( A1 => n19298, A2 => n16922, B1 => n16957, B2 => 
                           n16920, ZN => n1248);
   U1106 : OAI22_X1 port map( A1 => n19546, A2 => n16922, B1 => n16958, B2 => 
                           n16921, ZN => n1247);
   U1107 : OAI22_X1 port map( A1 => n19003, A2 => n16922, B1 => n16959, B2 => 
                           n16921, ZN => n1246);
   U1108 : OAI22_X1 port map( A1 => n19299, A2 => n16922, B1 => n16960, B2 => 
                           n16921, ZN => n1245);
   U1109 : OAI22_X1 port map( A1 => n18746, A2 => n16922, B1 => n16961, B2 => 
                           n16921, ZN => n1244);
   U1110 : OAI22_X1 port map( A1 => n19004, A2 => n16922, B1 => n16962, B2 => 
                           n16921, ZN => n1243);
   U1111 : OAI22_X1 port map( A1 => n19547, A2 => n16922, B1 => n16963, B2 => 
                           n16921, ZN => n1242);
   U1112 : OAI22_X1 port map( A1 => n19300, A2 => n16922, B1 => n16964, B2 => 
                           n16921, ZN => n1241);
   U1113 : OAI22_X1 port map( A1 => n19301, A2 => n16922, B1 => n16965, B2 => 
                           n16921, ZN => n1240);
   U1114 : OAI22_X1 port map( A1 => n19548, A2 => n16922, B1 => n16967, B2 => 
                           n16921, ZN => n1239);
   U1115 : NAND2_X1 port map( A1 => n16923, A2 => n16932, ZN => n16924);
   U1116 : CLKBUF_X1 port map( A => n16927, Z => n16925);
   U1117 : CLKBUF_X1 port map( A => n16924, Z => n16926);
   U1118 : OAI22_X1 port map( A1 => n18535, A2 => n16925, B1 => n16934, B2 => 
                           n16926, ZN => n1238);
   U1119 : OAI22_X1 port map( A1 => n18747, A2 => n16927, B1 => n16935, B2 => 
                           n16924, ZN => n1237);
   U1120 : OAI22_X1 port map( A1 => n19005, A2 => n16925, B1 => n16936, B2 => 
                           n16926, ZN => n1236);
   U1121 : OAI22_X1 port map( A1 => n18748, A2 => n16927, B1 => n16937, B2 => 
                           n16924, ZN => n1235);
   U1122 : OAI22_X1 port map( A1 => n19006, A2 => n16925, B1 => n16938, B2 => 
                           n16926, ZN => n1234);
   U1123 : OAI22_X1 port map( A1 => n19007, A2 => n16927, B1 => n16939, B2 => 
                           n16924, ZN => n1233);
   U1124 : OAI22_X1 port map( A1 => n19008, A2 => n16925, B1 => n16940, B2 => 
                           n16926, ZN => n1232);
   U1125 : OAI22_X1 port map( A1 => n19009, A2 => n16927, B1 => n16941, B2 => 
                           n16924, ZN => n1231);
   U1126 : OAI22_X1 port map( A1 => n19010, A2 => n16925, B1 => n16942, B2 => 
                           n16926, ZN => n1230);
   U1127 : OAI22_X1 port map( A1 => n18749, A2 => n16927, B1 => n16943, B2 => 
                           n16924, ZN => n1229);
   U1128 : OAI22_X1 port map( A1 => n19011, A2 => n16927, B1 => n16944, B2 => 
                           n16924, ZN => n1228);
   U1129 : OAI22_X1 port map( A1 => n18750, A2 => n16927, B1 => n16945, B2 => 
                           n16926, ZN => n1227);
   U1130 : OAI22_X1 port map( A1 => n18751, A2 => n16925, B1 => n16946, B2 => 
                           n16924, ZN => n1226);
   U1131 : OAI22_X1 port map( A1 => n19012, A2 => n16925, B1 => n16947, B2 => 
                           n16926, ZN => n1225);
   U1132 : OAI22_X1 port map( A1 => n19013, A2 => n16925, B1 => n16948, B2 => 
                           n16924, ZN => n1224);
   U1133 : OAI22_X1 port map( A1 => n19014, A2 => n16925, B1 => n16949, B2 => 
                           n16926, ZN => n1223);
   U1134 : OAI22_X1 port map( A1 => n18752, A2 => n16925, B1 => n16950, B2 => 
                           n16924, ZN => n1222);
   U1135 : OAI22_X1 port map( A1 => n19015, A2 => n16925, B1 => n16951, B2 => 
                           n16924, ZN => n1221);
   U1136 : OAI22_X1 port map( A1 => n19016, A2 => n16925, B1 => n16952, B2 => 
                           n16924, ZN => n1220);
   U1137 : OAI22_X1 port map( A1 => n19017, A2 => n16925, B1 => n16953, B2 => 
                           n16924, ZN => n1219);
   U1138 : OAI22_X1 port map( A1 => n19018, A2 => n16925, B1 => n16954, B2 => 
                           n16924, ZN => n1218);
   U1139 : OAI22_X1 port map( A1 => n18753, A2 => n16925, B1 => n16955, B2 => 
                           n16924, ZN => n1217);
   U1140 : OAI22_X1 port map( A1 => n18754, A2 => n16925, B1 => n16957, B2 => 
                           n16924, ZN => n1216);
   U1141 : OAI22_X1 port map( A1 => n18755, A2 => n16925, B1 => n16958, B2 => 
                           n16926, ZN => n1215);
   U1142 : OAI22_X1 port map( A1 => n19019, A2 => n16927, B1 => n16959, B2 => 
                           n16926, ZN => n1214);
   U1143 : OAI22_X1 port map( A1 => n19020, A2 => n16927, B1 => n16960, B2 => 
                           n16926, ZN => n1213);
   U1144 : OAI22_X1 port map( A1 => n18756, A2 => n16927, B1 => n16961, B2 => 
                           n16926, ZN => n1212);
   U1145 : OAI22_X1 port map( A1 => n19021, A2 => n16927, B1 => n16962, B2 => 
                           n16926, ZN => n1211);
   U1146 : OAI22_X1 port map( A1 => n19022, A2 => n16927, B1 => n16963, B2 => 
                           n16926, ZN => n1210);
   U1147 : OAI22_X1 port map( A1 => n18757, A2 => n16927, B1 => n16964, B2 => 
                           n16926, ZN => n1209);
   U1148 : OAI22_X1 port map( A1 => n19023, A2 => n16927, B1 => n16965, B2 => 
                           n16926, ZN => n1208);
   U1149 : OAI22_X1 port map( A1 => n18758, A2 => n16927, B1 => n16967, B2 => 
                           n16926, ZN => n1207);
   U1150 : NAND2_X1 port map( A1 => n16928, A2 => n16932, ZN => n16929);
   U1151 : CLKBUF_X1 port map( A => n16929, Z => n16930);
   U1152 : OAI22_X1 port map( A1 => n19051, A2 => n16931, B1 => n16934, B2 => 
                           n16930, ZN => n1206);
   U1153 : OAI22_X1 port map( A1 => n18759, A2 => n16931, B1 => n16935, B2 => 
                           n16929, ZN => n1205);
   U1154 : OAI22_X1 port map( A1 => n19549, A2 => n16931, B1 => n16936, B2 => 
                           n16930, ZN => n1204);
   U1155 : OAI22_X1 port map( A1 => n19550, A2 => n16931, B1 => n16937, B2 => 
                           n16929, ZN => n1203);
   U1156 : OAI22_X1 port map( A1 => n18760, A2 => n16931, B1 => n16938, B2 => 
                           n16930, ZN => n1202);
   U1157 : OAI22_X1 port map( A1 => n18761, A2 => n16931, B1 => n16939, B2 => 
                           n16929, ZN => n1201);
   U1158 : OAI22_X1 port map( A1 => n18762, A2 => n16931, B1 => n16940, B2 => 
                           n16930, ZN => n1200);
   U1159 : OAI22_X1 port map( A1 => n19024, A2 => n16931, B1 => n16941, B2 => 
                           n16929, ZN => n1199);
   U1160 : OAI22_X1 port map( A1 => n18763, A2 => n16931, B1 => n16942, B2 => 
                           n16930, ZN => n1198);
   U1161 : OAI22_X1 port map( A1 => n19302, A2 => n16931, B1 => n16943, B2 => 
                           n16929, ZN => n1197);
   U1162 : OAI22_X1 port map( A1 => n19303, A2 => n16931, B1 => n16944, B2 => 
                           n16929, ZN => n1196);
   U1163 : OAI22_X1 port map( A1 => n18764, A2 => n16931, B1 => n16945, B2 => 
                           n16930, ZN => n1195);
   U1164 : OAI22_X1 port map( A1 => n19025, A2 => n16931, B1 => n16946, B2 => 
                           n16929, ZN => n1194);
   U1165 : OAI22_X1 port map( A1 => n19026, A2 => n16931, B1 => n16947, B2 => 
                           n16930, ZN => n1193);
   U1166 : OAI22_X1 port map( A1 => n19027, A2 => n16931, B1 => n16948, B2 => 
                           n16929, ZN => n1192);
   U1167 : OAI22_X1 port map( A1 => n18765, A2 => n16931, B1 => n16949, B2 => 
                           n16930, ZN => n1191);
   U1168 : OAI22_X1 port map( A1 => n19551, A2 => n16931, B1 => n16950, B2 => 
                           n16929, ZN => n1190);
   U1169 : OAI22_X1 port map( A1 => n19028, A2 => n16931, B1 => n16951, B2 => 
                           n16929, ZN => n1189);
   U1170 : OAI22_X1 port map( A1 => n19552, A2 => n16931, B1 => n16952, B2 => 
                           n16929, ZN => n1188);
   U1171 : OAI22_X1 port map( A1 => n18766, A2 => n16931, B1 => n16953, B2 => 
                           n16929, ZN => n1187);
   U1172 : OAI22_X1 port map( A1 => n18767, A2 => n16931, B1 => n16954, B2 => 
                           n16929, ZN => n1186);
   U1173 : OAI22_X1 port map( A1 => n18768, A2 => n16931, B1 => n16955, B2 => 
                           n16929, ZN => n1185);
   U1174 : OAI22_X1 port map( A1 => n19553, A2 => n16931, B1 => n16957, B2 => 
                           n16929, ZN => n1184);
   U1175 : OAI22_X1 port map( A1 => n19029, A2 => n16931, B1 => n16958, B2 => 
                           n16930, ZN => n1183);
   U1176 : OAI22_X1 port map( A1 => n19030, A2 => n16931, B1 => n16959, B2 => 
                           n16930, ZN => n1182);
   U1177 : OAI22_X1 port map( A1 => n19031, A2 => n16931, B1 => n16960, B2 => 
                           n16930, ZN => n1181);
   U1178 : OAI22_X1 port map( A1 => n18769, A2 => n16931, B1 => n16961, B2 => 
                           n16930, ZN => n1180);
   U1179 : OAI22_X1 port map( A1 => n19032, A2 => n16931, B1 => n16962, B2 => 
                           n16930, ZN => n1179);
   U1180 : OAI22_X1 port map( A1 => n18770, A2 => n16931, B1 => n16963, B2 => 
                           n16930, ZN => n1178);
   U1181 : OAI22_X1 port map( A1 => n19033, A2 => n16931, B1 => n16964, B2 => 
                           n16930, ZN => n1177);
   U1182 : OAI22_X1 port map( A1 => n19554, A2 => n16931, B1 => n16965, B2 => 
                           n16930, ZN => n1176);
   U1183 : OAI22_X1 port map( A1 => n18771, A2 => n16931, B1 => n16967, B2 => 
                           n16930, ZN => n1175);
   U1184 : NAND2_X1 port map( A1 => n16933, A2 => n16932, ZN => n16956);
   U1185 : CLKBUF_X1 port map( A => n16956, Z => n16966);
   U1186 : OAI22_X1 port map( A1 => n18536, A2 => n16968, B1 => n16934, B2 => 
                           n16966, ZN => n1174);
   U1187 : OAI22_X1 port map( A1 => n18772, A2 => n16968, B1 => n16935, B2 => 
                           n16956, ZN => n1173);
   U1188 : OAI22_X1 port map( A1 => n18773, A2 => n16968, B1 => n16936, B2 => 
                           n16966, ZN => n1172);
   U1189 : OAI22_X1 port map( A1 => n19034, A2 => n16968, B1 => n16937, B2 => 
                           n16956, ZN => n1171);
   U1190 : OAI22_X1 port map( A1 => n19035, A2 => n16968, B1 => n16938, B2 => 
                           n16966, ZN => n1170);
   U1191 : OAI22_X1 port map( A1 => n18774, A2 => n16968, B1 => n16939, B2 => 
                           n16956, ZN => n1169);
   U1192 : OAI22_X1 port map( A1 => n19036, A2 => n16968, B1 => n16940, B2 => 
                           n16966, ZN => n1168);
   U1193 : OAI22_X1 port map( A1 => n18775, A2 => n16968, B1 => n16941, B2 => 
                           n16956, ZN => n1167);
   U1194 : OAI22_X1 port map( A1 => n19037, A2 => n16968, B1 => n16942, B2 => 
                           n16966, ZN => n1166);
   U1195 : OAI22_X1 port map( A1 => n19038, A2 => n16968, B1 => n16943, B2 => 
                           n16956, ZN => n1165);
   U1196 : OAI22_X1 port map( A1 => n18776, A2 => n16968, B1 => n16944, B2 => 
                           n16956, ZN => n1164);
   U1197 : OAI22_X1 port map( A1 => n18777, A2 => n16968, B1 => n16945, B2 => 
                           n16966, ZN => n1163);
   U1198 : OAI22_X1 port map( A1 => n19039, A2 => n16968, B1 => n16946, B2 => 
                           n16956, ZN => n1162);
   U1199 : OAI22_X1 port map( A1 => n19040, A2 => n16968, B1 => n16947, B2 => 
                           n16966, ZN => n1161);
   U1200 : OAI22_X1 port map( A1 => n18778, A2 => n16968, B1 => n16948, B2 => 
                           n16956, ZN => n1160);
   U1201 : OAI22_X1 port map( A1 => n18779, A2 => n16968, B1 => n16949, B2 => 
                           n16966, ZN => n1159);
   U1202 : OAI22_X1 port map( A1 => n19041, A2 => n16968, B1 => n16950, B2 => 
                           n16956, ZN => n1158);
   U1203 : OAI22_X1 port map( A1 => n18780, A2 => n16968, B1 => n16951, B2 => 
                           n16956, ZN => n1157);
   U1204 : OAI22_X1 port map( A1 => n18781, A2 => n16968, B1 => n16952, B2 => 
                           n16956, ZN => n1156);
   U1205 : OAI22_X1 port map( A1 => n19042, A2 => n16968, B1 => n16953, B2 => 
                           n16956, ZN => n1155);
   U1206 : OAI22_X1 port map( A1 => n18782, A2 => n16968, B1 => n16954, B2 => 
                           n16956, ZN => n1154);
   U1207 : OAI22_X1 port map( A1 => n19043, A2 => n16968, B1 => n16955, B2 => 
                           n16956, ZN => n1153);
   U1208 : OAI22_X1 port map( A1 => n19044, A2 => n16968, B1 => n16957, B2 => 
                           n16956, ZN => n1152);
   U1209 : OAI22_X1 port map( A1 => n18783, A2 => n16968, B1 => n16958, B2 => 
                           n16966, ZN => n1151);
   U1210 : OAI22_X1 port map( A1 => n18784, A2 => n16968, B1 => n16959, B2 => 
                           n16966, ZN => n1150);
   U1211 : OAI22_X1 port map( A1 => n19045, A2 => n16968, B1 => n16960, B2 => 
                           n16966, ZN => n1149);
   U1212 : OAI22_X1 port map( A1 => n19555, A2 => n16968, B1 => n16961, B2 => 
                           n16966, ZN => n1148);
   U1213 : OAI22_X1 port map( A1 => n18785, A2 => n16968, B1 => n16962, B2 => 
                           n16966, ZN => n1147);
   U1214 : OAI22_X1 port map( A1 => n19046, A2 => n16968, B1 => n16963, B2 => 
                           n16966, ZN => n1146);
   U1215 : OAI22_X1 port map( A1 => n18786, A2 => n16968, B1 => n16964, B2 => 
                           n16966, ZN => n1145);
   U1216 : OAI22_X1 port map( A1 => n18787, A2 => n16968, B1 => n16965, B2 => 
                           n16966, ZN => n1144);
   U1217 : OAI22_X1 port map( A1 => n19304, A2 => n16968, B1 => n16967, B2 => 
                           n16966, ZN => n1143);
   U1218 : NAND3_X1 port map( A1 => n16783, A2 => ENABLE, A3 => RD2, ZN => 
                           n17749);
   U1219 : INV_X1 port map( A => ADD_RD2(0), ZN => n16969);
   U1220 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), A3 => n16969,
                           ZN => n16986);
   U1221 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n16976)
                           ;
   U1222 : NOR2_X1 port map( A1 => n16986, A2 => n16976, ZN => n17476);
   U1223 : INV_X1 port map( A => ADD_RD2(3), ZN => n16994);
   U1224 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n16994, ZN => n16977);
   U1225 : INV_X1 port map( A => ADD_RD2(2), ZN => n16974);
   U1226 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => n16969, A3 => n16974, ZN 
                           => n16985);
   U1227 : NOR2_X1 port map( A1 => n16977, A2 => n16985, ZN => n17453);
   U1228 : CLKBUF_X1 port map( A => n17453, Z => n17711);
   U1229 : AOI22_X1 port map( A1 => REGISTERS_30_31_port, A2 => n17476, B1 => 
                           REGISTERS_18_31_port, B2 => n17711, ZN => n16973);
   U1230 : NOR2_X1 port map( A1 => n16976, A2 => n16985, ZN => n17698);
   U1231 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n16974,
                           ZN => n16987);
   U1232 : NOR2_X1 port map( A1 => n16977, A2 => n16987, ZN => n17477);
   U1233 : CLKBUF_X1 port map( A => n17477, Z => n17713);
   U1234 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n17698, B1 => 
                           REGISTERS_19_31_port, B2 => n17713, ZN => n16972);
   U1235 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), ZN => n16975);
   U1236 : NAND2_X1 port map( A1 => n16975, A2 => n16969, ZN => n16989);
   U1237 : NOR2_X1 port map( A1 => n16976, A2 => n16989, ZN => n17542);
   U1238 : OR3_X1 port map( A1 => n16974, A2 => n16969, A3 => ADD_RD2(1), ZN =>
                           n17190);
   U1239 : NOR2_X1 port map( A1 => n17190, A2 => n16976, ZN => n17699);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n17542, B1 => 
                           REGISTERS_29_31_port, B2 => n17699, ZN => n16971);
   U1241 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(1), ZN => n16988);
   U1242 : NOR2_X1 port map( A1 => n16977, A2 => n16988, ZN => n17291);
   U1243 : NOR2_X1 port map( A1 => n16976, A2 => n16988, ZN => n17700);
   U1244 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n17291, B1 => 
                           REGISTERS_31_31_port, B2 => n17700, ZN => n16970);
   U1245 : NAND4_X1 port map( A1 => n16973, A2 => n16972, A3 => n16971, A4 => 
                           n16970, ZN => n16983);
   U1246 : OR3_X1 port map( A1 => n16974, A2 => ADD_RD2(0), A3 => ADD_RD2(1), 
                           ZN => n17017);
   U1247 : NOR2_X1 port map( A1 => n16976, A2 => n17017, ZN => n17594);
   U1248 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n16975, ZN => n16984);
   U1249 : NOR2_X1 port map( A1 => n16976, A2 => n16984, ZN => n17452);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n17594, B1 => 
                           REGISTERS_25_31_port, B2 => n17452, ZN => n16981);
   U1251 : NOR2_X1 port map( A1 => n16977, A2 => n16986, ZN => n17710);
   U1252 : NOR2_X1 port map( A1 => n16977, A2 => n17190, ZN => n17666);
   U1253 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n17710, B1 => 
                           REGISTERS_21_31_port, B2 => n17666, ZN => n16980);
   U1254 : NOR2_X1 port map( A1 => n16977, A2 => n17017, ZN => n17615);
   U1255 : NOR2_X1 port map( A1 => n16977, A2 => n16984, ZN => n17701);
   U1256 : CLKBUF_X1 port map( A => n17701, Z => n17671);
   U1257 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n17615, B1 => 
                           REGISTERS_17_31_port, B2 => n17671, ZN => n16979);
   U1258 : NOR2_X1 port map( A1 => n16976, A2 => n16987, ZN => n17614);
   U1259 : NOR2_X1 port map( A1 => n16977, A2 => n16989, ZN => n17709);
   U1260 : CLKBUF_X1 port map( A => n17709, Z => n17613);
   U1261 : AOI22_X1 port map( A1 => REGISTERS_27_31_port, A2 => n17614, B1 => 
                           REGISTERS_16_31_port, B2 => n17613, ZN => n16978);
   U1262 : NAND4_X1 port map( A1 => n16981, A2 => n16980, A3 => n16979, A4 => 
                           n16978, ZN => n16982);
   U1263 : NOR2_X1 port map( A1 => n16983, A2 => n16982, ZN => n17002);
   U1264 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n17694, 
                           ZN => n17746);
   U1265 : CLKBUF_X1 port map( A => n17746, Z => n17563);
   U1266 : INV_X1 port map( A => n16984, ZN => n17733);
   U1267 : CLKBUF_X1 port map( A => n17733, Z => n17723);
   U1268 : INV_X1 port map( A => n16985, ZN => n17731);
   U1269 : CLKBUF_X1 port map( A => n17731, Z => n17724);
   U1270 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_31_port, B1 => 
                           n17724, B2 => REGISTERS_2_31_port, ZN => n16993);
   U1271 : INV_X1 port map( A => n16986, ZN => n17649);
   U1272 : CLKBUF_X1 port map( A => n17649, Z => n17439);
   U1273 : INV_X1 port map( A => n17190, ZN => n17679);
   U1274 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_31_port, B1 => 
                           n17679, B2 => REGISTERS_5_31_port, ZN => n16992);
   U1275 : INV_X1 port map( A => n16987, ZN => n17738);
   U1276 : CLKBUF_X1 port map( A => n17738, Z => n17726);
   U1277 : INV_X1 port map( A => n16988, ZN => n17650);
   U1278 : CLKBUF_X1 port map( A => n17650, Z => n17438);
   U1279 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_31_port, B1 => 
                           n17438, B2 => REGISTERS_7_31_port, ZN => n16991);
   U1280 : INV_X1 port map( A => n17017, ZN => n17656);
   U1281 : INV_X1 port map( A => n16989, ZN => n17737);
   U1282 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_4_31_port, B1 => 
                           n17737, B2 => REGISTERS_0_31_port, ZN => n16990);
   U1283 : NAND4_X1 port map( A1 => n16993, A2 => n16992, A3 => n16991, A4 => 
                           n16990, ZN => n17000);
   U1284 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n16994, A3 => n17694, ZN 
                           => n17744);
   U1285 : CLKBUF_X1 port map( A => n17744, Z => n17585);
   U1286 : INV_X1 port map( A => n17190, ZN => n17721);
   U1287 : CLKBUF_X1 port map( A => n17737, Z => n17685);
   U1288 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_31_port, B1 => 
                           n17685, B2 => REGISTERS_8_31_port, ZN => n16998);
   U1289 : INV_X1 port map( A => n17017, ZN => n17736);
   U1290 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_31_port, B1 => 
                           n17736, B2 => REGISTERS_12_31_port, ZN => n16997);
   U1291 : CLKBUF_X1 port map( A => n17738, Z => n17651);
   U1292 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_31_port, B1 => 
                           n17651, B2 => REGISTERS_11_31_port, ZN => n16996);
   U1293 : AOI22_X1 port map( A1 => n17724, A2 => REGISTERS_10_31_port, B1 => 
                           n17438, B2 => REGISTERS_15_31_port, ZN => n16995);
   U1294 : NAND4_X1 port map( A1 => n16998, A2 => n16997, A3 => n16996, A4 => 
                           n16995, ZN => n16999);
   U1295 : AOI22_X1 port map( A1 => n17563, A2 => n17000, B1 => n17585, B2 => 
                           n16999, ZN => n17001);
   U1296 : OAI21_X1 port map( B1 => n17694, B2 => n17002, A => n17001, ZN => 
                           N448);
   U1297 : CLKBUF_X1 port map( A => n17291, Z => n17695);
   U1298 : CLKBUF_X1 port map( A => n17699, Z => n17496);
   U1299 : AOI22_X1 port map( A1 => n17695, A2 => REGISTERS_23_30_port, B1 => 
                           n17496, B2 => REGISTERS_29_30_port, ZN => n17006);
   U1300 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_30_port, B1 => 
                           n17698, B2 => REGISTERS_26_30_port, ZN => n17005);
   U1301 : CLKBUF_X1 port map( A => n17614, Z => n17696);
   U1302 : CLKBUF_X1 port map( A => n17476, Z => n17697);
   U1303 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_30_port, B1 => 
                           n17697, B2 => REGISTERS_30_30_port, ZN => n17004);
   U1304 : CLKBUF_X1 port map( A => n17700, Z => n17665);
   U1305 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_30_port, B1 => 
                           n17665, B2 => REGISTERS_31_30_port, ZN => n17003);
   U1306 : NAND4_X1 port map( A1 => n17006, A2 => n17005, A3 => n17004, A4 => 
                           n17003, ZN => n17012);
   U1307 : CLKBUF_X1 port map( A => n17710, Z => n17497);
   U1308 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_30_port, B1 => 
                           n17452, B2 => REGISTERS_25_30_port, ZN => n17010);
   U1309 : CLKBUF_X1 port map( A => n17594, Z => n17712);
   U1310 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_30_port, B1 => 
                           n17701, B2 => REGISTERS_17_30_port, ZN => n17009);
   U1311 : CLKBUF_X1 port map( A => n17542, Z => n17707);
   U1312 : AOI22_X1 port map( A1 => n17666, A2 => REGISTERS_21_30_port, B1 => 
                           n17707, B2 => REGISTERS_24_30_port, ZN => n17008);
   U1313 : CLKBUF_X1 port map( A => n17615, Z => n17702);
   U1314 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_30_port, B1 => 
                           n17711, B2 => REGISTERS_18_30_port, ZN => n17007);
   U1315 : NAND4_X1 port map( A1 => n17010, A2 => n17009, A3 => n17008, A4 => 
                           n17007, ZN => n17011);
   U1316 : NOR2_X1 port map( A1 => n17012, A2 => n17011, ZN => n17025);
   U1317 : CLKBUF_X1 port map( A => n17737, Z => n17722);
   U1318 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_0_30_port, B1 => 
                           n17438, B2 => REGISTERS_7_30_port, ZN => n17016);
   U1319 : CLKBUF_X1 port map( A => n17731, Z => n17678);
   U1320 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_4_30_port, B1 => 
                           n17678, B2 => REGISTERS_2_30_port, ZN => n17015);
   U1321 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_30_port, B1 => 
                           n17651, B2 => REGISTERS_3_30_port, ZN => n17014);
   U1322 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_30_port, B1 => 
                           n17679, B2 => REGISTERS_5_30_port, ZN => n17013);
   U1323 : NAND4_X1 port map( A1 => n17016, A2 => n17015, A3 => n17014, A4 => 
                           n17013, ZN => n17023);
   U1324 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_30_port, B1 => 
                           n17651, B2 => REGISTERS_11_30_port, ZN => n17021);
   U1325 : INV_X1 port map( A => n17017, ZN => n17725);
   U1326 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_30_port, B1 => 
                           n17438, B2 => REGISTERS_15_30_port, ZN => n17020);
   U1327 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_30_port, B1 => 
                           n17679, B2 => REGISTERS_13_30_port, ZN => n17019);
   U1328 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_8_30_port, B1 => 
                           n17678, B2 => REGISTERS_10_30_port, ZN => n17018);
   U1329 : NAND4_X1 port map( A1 => n17021, A2 => n17020, A3 => n17019, A4 => 
                           n17018, ZN => n17022);
   U1330 : AOI22_X1 port map( A1 => n17563, A2 => n17023, B1 => n17585, B2 => 
                           n17022, ZN => n17024);
   U1331 : OAI21_X1 port map( B1 => n17694, B2 => n17025, A => n17024, ZN => 
                           N447);
   U1332 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_29_port, B1 => 
                           n17713, B2 => REGISTERS_19_29_port, ZN => n17029);
   U1333 : AOI22_X1 port map( A1 => n17666, A2 => REGISTERS_21_29_port, B1 => 
                           n17695, B2 => REGISTERS_23_29_port, ZN => n17028);
   U1334 : CLKBUF_X1 port map( A => n17452, Z => n17714);
   U1335 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_29_port, B1 => 
                           n17700, B2 => REGISTERS_31_29_port, ZN => n17027);
   U1336 : CLKBUF_X1 port map( A => n17698, Z => n17638);
   U1337 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_29_port, B1 => 
                           n17453, B2 => REGISTERS_18_29_port, ZN => n17026);
   U1338 : NAND4_X1 port map( A1 => n17029, A2 => n17028, A3 => n17027, A4 => 
                           n17026, ZN => n17035);
   U1339 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_29_port, B1 => 
                           n17701, B2 => REGISTERS_17_29_port, ZN => n17033);
   U1340 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_29_port, B1 => 
                           n17496, B2 => REGISTERS_29_29_port, ZN => n17032);
   U1341 : AOI22_X1 port map( A1 => n17697, A2 => REGISTERS_30_29_port, B1 => 
                           n17542, B2 => REGISTERS_24_29_port, ZN => n17031);
   U1342 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_29_port, B1 => 
                           n17615, B2 => REGISTERS_20_29_port, ZN => n17030);
   U1343 : NAND4_X1 port map( A1 => n17033, A2 => n17032, A3 => n17031, A4 => 
                           n17030, ZN => n17034);
   U1344 : NOR2_X1 port map( A1 => n17035, A2 => n17034, ZN => n17047);
   U1345 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_29_port, B1 => 
                           n17678, B2 => REGISTERS_2_29_port, ZN => n17039);
   U1346 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_29_port, B1 => 
                           n17438, B2 => REGISTERS_7_29_port, ZN => n17038);
   U1347 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_29_port, B1 => 
                           n17723, B2 => REGISTERS_1_29_port, ZN => n17037);
   U1348 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_29_port, B1 => 
                           n17685, B2 => REGISTERS_0_29_port, ZN => n17036);
   U1349 : NAND4_X1 port map( A1 => n17039, A2 => n17038, A3 => n17037, A4 => 
                           n17036, ZN => n17045);
   U1350 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_29_port, B1 => 
                           n17438, B2 => REGISTERS_15_29_port, ZN => n17043);
   U1351 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_29_port, B1 => 
                           n17685, B2 => REGISTERS_8_29_port, ZN => n17042);
   U1352 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_29_port, B1 => 
                           n17736, B2 => REGISTERS_12_29_port, ZN => n17041);
   U1353 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_29_port, B1 => 
                           n17678, B2 => REGISTERS_10_29_port, ZN => n17040);
   U1354 : NAND4_X1 port map( A1 => n17043, A2 => n17042, A3 => n17041, A4 => 
                           n17040, ZN => n17044);
   U1355 : AOI22_X1 port map( A1 => n17563, A2 => n17045, B1 => n17585, B2 => 
                           n17044, ZN => n17046);
   U1356 : OAI21_X1 port map( B1 => n17694, B2 => n17047, A => n17046, ZN => 
                           N446);
   U1357 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_28_port, B1 => 
                           n17291, B2 => REGISTERS_23_28_port, ZN => n17051);
   U1358 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_28_port, B1 => 
                           n17700, B2 => REGISTERS_31_28_port, ZN => n17050);
   U1359 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_28_port, B1 => 
                           n17496, B2 => REGISTERS_29_28_port, ZN => n17049);
   U1360 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_28_port, B1 => 
                           n17453, B2 => REGISTERS_18_28_port, ZN => n17048);
   U1361 : NAND4_X1 port map( A1 => n17051, A2 => n17050, A3 => n17049, A4 => 
                           n17048, ZN => n17057);
   U1362 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_28_port, B1 => 
                           n17701, B2 => REGISTERS_17_28_port, ZN => n17055);
   U1363 : AOI22_X1 port map( A1 => n17697, A2 => REGISTERS_30_28_port, B1 => 
                           n17542, B2 => REGISTERS_24_28_port, ZN => n17054);
   U1364 : AOI22_X1 port map( A1 => n17614, A2 => REGISTERS_27_28_port, B1 => 
                           n17709, B2 => REGISTERS_16_28_port, ZN => n17053);
   U1365 : AOI22_X1 port map( A1 => n17666, A2 => REGISTERS_21_28_port, B1 => 
                           n17594, B2 => REGISTERS_28_28_port, ZN => n17052);
   U1366 : NAND4_X1 port map( A1 => n17055, A2 => n17054, A3 => n17053, A4 => 
                           n17052, ZN => n17056);
   U1367 : NOR2_X1 port map( A1 => n17057, A2 => n17056, ZN => n17069);
   U1368 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_28_port, B1 => 
                           n17651, B2 => REGISTERS_3_28_port, ZN => n17061);
   U1369 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_28_port, B1 => 
                           n17685, B2 => REGISTERS_0_28_port, ZN => n17060);
   U1370 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_28_port, B1 => 
                           n17438, B2 => REGISTERS_7_28_port, ZN => n17059);
   U1371 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_28_port, B1 => 
                           n17678, B2 => REGISTERS_2_28_port, ZN => n17058);
   U1372 : NAND4_X1 port map( A1 => n17061, A2 => n17060, A3 => n17059, A4 => 
                           n17058, ZN => n17067);
   U1373 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_28_port, B1 => 
                           n17438, B2 => REGISTERS_15_28_port, ZN => n17065);
   U1374 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_28_port, B1 => 
                           n17731, B2 => REGISTERS_10_28_port, ZN => n17064);
   U1375 : CLKBUF_X1 port map( A => n17733, Z => n17684);
   U1376 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_28_port, B1 => 
                           n17684, B2 => REGISTERS_9_28_port, ZN => n17063);
   U1377 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_28_port, B1 => 
                           n17685, B2 => REGISTERS_8_28_port, ZN => n17062);
   U1378 : NAND4_X1 port map( A1 => n17065, A2 => n17064, A3 => n17063, A4 => 
                           n17062, ZN => n17066);
   U1379 : AOI22_X1 port map( A1 => n17563, A2 => n17067, B1 => n17585, B2 => 
                           n17066, ZN => n17068);
   U1380 : OAI21_X1 port map( B1 => n17694, B2 => n17069, A => n17068, ZN => 
                           N445);
   U1381 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_27_port, B1 => 
                           n17698, B2 => REGISTERS_26_27_port, ZN => n17073);
   U1382 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_27_port, B1 => 
                           n17291, B2 => REGISTERS_23_27_port, ZN => n17072);
   U1383 : AOI22_X1 port map( A1 => n17594, A2 => REGISTERS_28_27_port, B1 => 
                           n17476, B2 => REGISTERS_30_27_port, ZN => n17071);
   U1384 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_27_port, B1 => 
                           n17453, B2 => REGISTERS_18_27_port, ZN => n17070);
   U1385 : NAND4_X1 port map( A1 => n17073, A2 => n17072, A3 => n17071, A4 => 
                           n17070, ZN => n17079);
   U1386 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_27_port, B1 => 
                           n17700, B2 => REGISTERS_31_27_port, ZN => n17077);
   U1387 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_27_port, B1 => 
                           n17542, B2 => REGISTERS_24_27_port, ZN => n17076);
   U1388 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_27_port, B1 => 
                           n17496, B2 => REGISTERS_29_27_port, ZN => n17075);
   U1389 : AOI22_X1 port map( A1 => n17666, A2 => REGISTERS_21_27_port, B1 => 
                           n17477, B2 => REGISTERS_19_27_port, ZN => n17074);
   U1390 : NAND4_X1 port map( A1 => n17077, A2 => n17076, A3 => n17075, A4 => 
                           n17074, ZN => n17078);
   U1391 : NOR2_X1 port map( A1 => n17079, A2 => n17078, ZN => n17091);
   U1392 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_27_port, B1 => 
                           n17438, B2 => REGISTERS_7_27_port, ZN => n17083);
   U1393 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_27_port, B1 => 
                           n17684, B2 => REGISTERS_1_27_port, ZN => n17082);
   U1394 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_27_port, B1 => 
                           n17651, B2 => REGISTERS_3_27_port, ZN => n17081);
   U1395 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_0_27_port, B1 => 
                           n17678, B2 => REGISTERS_2_27_port, ZN => n17080);
   U1396 : NAND4_X1 port map( A1 => n17083, A2 => n17082, A3 => n17081, A4 => 
                           n17080, ZN => n17089);
   U1397 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_27_port, B1 => 
                           n17651, B2 => REGISTERS_11_27_port, ZN => n17087);
   U1398 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_27_port, B1 => 
                           n17731, B2 => REGISTERS_10_27_port, ZN => n17086);
   U1399 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_27_port, B1 => 
                           n17721, B2 => REGISTERS_13_27_port, ZN => n17085);
   U1400 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_8_27_port, B1 => 
                           n17438, B2 => REGISTERS_15_27_port, ZN => n17084);
   U1401 : NAND4_X1 port map( A1 => n17087, A2 => n17086, A3 => n17085, A4 => 
                           n17084, ZN => n17088);
   U1402 : AOI22_X1 port map( A1 => n17563, A2 => n17089, B1 => n17585, B2 => 
                           n17088, ZN => n17090);
   U1403 : OAI21_X1 port map( B1 => n17694, B2 => n17091, A => n17090, ZN => 
                           N444);
   U1404 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_26_port, B1 => 
                           n17476, B2 => REGISTERS_30_26_port, ZN => n17095);
   U1405 : CLKBUF_X1 port map( A => n17666, Z => n17708);
   U1406 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_26_port, B1 => 
                           n17477, B2 => REGISTERS_19_26_port, ZN => n17094);
   U1407 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_26_port, B1 => 
                           n17615, B2 => REGISTERS_20_26_port, ZN => n17093);
   U1408 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_26_port, B1 => 
                           n17700, B2 => REGISTERS_31_26_port, ZN => n17092);
   U1409 : NAND4_X1 port map( A1 => n17095, A2 => n17094, A3 => n17093, A4 => 
                           n17092, ZN => n17101);
   U1410 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_26_port, B1 => 
                           n17496, B2 => REGISTERS_29_26_port, ZN => n17099);
   U1411 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_26_port, B1 => 
                           n17291, B2 => REGISTERS_23_26_port, ZN => n17098);
   U1412 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_26_port, B1 => 
                           n17701, B2 => REGISTERS_17_26_port, ZN => n17097);
   U1413 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_26_port, B1 => 
                           n17542, B2 => REGISTERS_24_26_port, ZN => n17096);
   U1414 : NAND4_X1 port map( A1 => n17099, A2 => n17098, A3 => n17097, A4 => 
                           n17096, ZN => n17100);
   U1415 : NOR2_X1 port map( A1 => n17101, A2 => n17100, ZN => n17113);
   U1416 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_26_port, B1 => 
                           n17656, B2 => REGISTERS_4_26_port, ZN => n17105);
   U1417 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_26_port, B1 => 
                           n17438, B2 => REGISTERS_7_26_port, ZN => n17104);
   U1418 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_26_port, B1 => 
                           n17737, B2 => REGISTERS_0_26_port, ZN => n17103);
   U1419 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_26_port, B1 => 
                           n17678, B2 => REGISTERS_2_26_port, ZN => n17102);
   U1420 : NAND4_X1 port map( A1 => n17105, A2 => n17104, A3 => n17103, A4 => 
                           n17102, ZN => n17111);
   U1421 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_13_26_port, B1 => 
                           n17438, B2 => REGISTERS_15_26_port, ZN => n17109);
   U1422 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_26_port, B1 => 
                           n17738, B2 => REGISTERS_11_26_port, ZN => n17108);
   U1423 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_26_port, B1 => 
                           n17731, B2 => REGISTERS_10_26_port, ZN => n17107);
   U1424 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_26_port, B1 => 
                           n17685, B2 => REGISTERS_8_26_port, ZN => n17106);
   U1425 : NAND4_X1 port map( A1 => n17109, A2 => n17108, A3 => n17107, A4 => 
                           n17106, ZN => n17110);
   U1426 : AOI22_X1 port map( A1 => n17563, A2 => n17111, B1 => n17585, B2 => 
                           n17110, ZN => n17112);
   U1427 : OAI21_X1 port map( B1 => n17694, B2 => n17113, A => n17112, ZN => 
                           N443);
   U1428 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_25_port, B1 => 
                           n17476, B2 => REGISTERS_30_25_port, ZN => n17117);
   U1429 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_25_port, B1 => 
                           n17542, B2 => REGISTERS_24_25_port, ZN => n17116);
   U1430 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_25_port, B1 => 
                           n17477, B2 => REGISTERS_19_25_port, ZN => n17115);
   U1431 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_25_port, B1 => 
                           n17700, B2 => REGISTERS_31_25_port, ZN => n17114);
   U1432 : NAND4_X1 port map( A1 => n17117, A2 => n17116, A3 => n17115, A4 => 
                           n17114, ZN => n17123);
   U1433 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_25_port, B1 => 
                           n17615, B2 => REGISTERS_20_25_port, ZN => n17121);
   U1434 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_25_port, B1 => 
                           n17291, B2 => REGISTERS_23_25_port, ZN => n17120);
   U1435 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_25_port, B1 => 
                           n17671, B2 => REGISTERS_17_25_port, ZN => n17119);
   U1436 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_25_port, B1 => 
                           n17496, B2 => REGISTERS_29_25_port, ZN => n17118);
   U1437 : NAND4_X1 port map( A1 => n17121, A2 => n17120, A3 => n17119, A4 => 
                           n17118, ZN => n17122);
   U1438 : NOR2_X1 port map( A1 => n17123, A2 => n17122, ZN => n17135);
   U1439 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_25_port, B1 => 
                           n17737, B2 => REGISTERS_0_25_port, ZN => n17127);
   U1440 : AOI22_X1 port map( A1 => n17724, A2 => REGISTERS_2_25_port, B1 => 
                           n17438, B2 => REGISTERS_7_25_port, ZN => n17126);
   U1441 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_25_port, B1 => 
                           n17651, B2 => REGISTERS_3_25_port, ZN => n17125);
   U1442 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_25_port, B1 => 
                           n17684, B2 => REGISTERS_1_25_port, ZN => n17124);
   U1443 : NAND4_X1 port map( A1 => n17127, A2 => n17126, A3 => n17125, A4 => 
                           n17124, ZN => n17133);
   U1444 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_25_port, B1 => 
                           n17678, B2 => REGISTERS_10_25_port, ZN => n17131);
   U1445 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_13_25_port, B1 => 
                           n17738, B2 => REGISTERS_11_25_port, ZN => n17130);
   U1446 : CLKBUF_X1 port map( A => n17649, Z => n17734);
   U1447 : CLKBUF_X1 port map( A => n17650, Z => n17735);
   U1448 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_25_port, B1 => 
                           n17735, B2 => REGISTERS_15_25_port, ZN => n17129);
   U1449 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_25_port, B1 => 
                           n17685, B2 => REGISTERS_8_25_port, ZN => n17128);
   U1450 : NAND4_X1 port map( A1 => n17131, A2 => n17130, A3 => n17129, A4 => 
                           n17128, ZN => n17132);
   U1451 : AOI22_X1 port map( A1 => n17563, A2 => n17133, B1 => n17585, B2 => 
                           n17132, ZN => n17134);
   U1452 : OAI21_X1 port map( B1 => n17694, B2 => n17135, A => n17134, ZN => 
                           N442);
   U1453 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_24_port, B1 => 
                           n17615, B2 => REGISTERS_20_24_port, ZN => n17139);
   U1454 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_24_port, B1 => 
                           n17453, B2 => REGISTERS_18_24_port, ZN => n17138);
   U1455 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_24_port, B1 => 
                           n17614, B2 => REGISTERS_27_24_port, ZN => n17137);
   U1456 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_24_port, B1 => 
                           n17700, B2 => REGISTERS_31_24_port, ZN => n17136);
   U1457 : NAND4_X1 port map( A1 => n17139, A2 => n17138, A3 => n17137, A4 => 
                           n17136, ZN => n17145);
   U1458 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_24_port, B1 => 
                           n17291, B2 => REGISTERS_23_24_port, ZN => n17143);
   U1459 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_24_port, B1 => 
                           n17496, B2 => REGISTERS_29_24_port, ZN => n17142);
   U1460 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_24_port, B1 => 
                           n17476, B2 => REGISTERS_30_24_port, ZN => n17141);
   U1461 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_24_port, B1 => 
                           n17542, B2 => REGISTERS_24_24_port, ZN => n17140);
   U1462 : NAND4_X1 port map( A1 => n17143, A2 => n17142, A3 => n17141, A4 => 
                           n17140, ZN => n17144);
   U1463 : NOR2_X1 port map( A1 => n17145, A2 => n17144, ZN => n17157);
   U1464 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_24_port, B1 => 
                           n17684, B2 => REGISTERS_1_24_port, ZN => n17149);
   U1465 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_0_24_port, B1 => 
                           n17650, B2 => REGISTERS_7_24_port, ZN => n17148);
   U1466 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_24_port, B1 => 
                           n17731, B2 => REGISTERS_2_24_port, ZN => n17147);
   U1467 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_24_port, B1 => 
                           n17721, B2 => REGISTERS_5_24_port, ZN => n17146);
   U1468 : NAND4_X1 port map( A1 => n17149, A2 => n17148, A3 => n17147, A4 => 
                           n17146, ZN => n17155);
   U1469 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_9_24_port, B1 => 
                           n17438, B2 => REGISTERS_15_24_port, ZN => n17153);
   U1470 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_24_port, B1 => 
                           n17678, B2 => REGISTERS_10_24_port, ZN => n17152);
   U1471 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_24_port, B1 => 
                           n17651, B2 => REGISTERS_11_24_port, ZN => n17151);
   U1472 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_13_24_port, B1 => 
                           n17737, B2 => REGISTERS_8_24_port, ZN => n17150);
   U1473 : NAND4_X1 port map( A1 => n17153, A2 => n17152, A3 => n17151, A4 => 
                           n17150, ZN => n17154);
   U1474 : AOI22_X1 port map( A1 => n17563, A2 => n17155, B1 => n17585, B2 => 
                           n17154, ZN => n17156);
   U1475 : OAI21_X1 port map( B1 => n17694, B2 => n17157, A => n17156, ZN => 
                           N441);
   U1476 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_23_port, B1 => 
                           n17453, B2 => REGISTERS_18_23_port, ZN => n17161);
   U1477 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_23_port, B1 => 
                           n17476, B2 => REGISTERS_30_23_port, ZN => n17160);
   U1478 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_23_port, B1 => 
                           n17477, B2 => REGISTERS_19_23_port, ZN => n17159);
   U1479 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_23_port, B1 => 
                           n17542, B2 => REGISTERS_24_23_port, ZN => n17158);
   U1480 : NAND4_X1 port map( A1 => n17161, A2 => n17160, A3 => n17159, A4 => 
                           n17158, ZN => n17167);
   U1481 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_23_port, B1 => 
                           n17709, B2 => REGISTERS_16_23_port, ZN => n17165);
   U1482 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_23_port, B1 => 
                           n17615, B2 => REGISTERS_20_23_port, ZN => n17164);
   U1483 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_23_port, B1 => 
                           n17700, B2 => REGISTERS_31_23_port, ZN => n17163);
   U1484 : AOI22_X1 port map( A1 => n17695, A2 => REGISTERS_23_23_port, B1 => 
                           n17496, B2 => REGISTERS_29_23_port, ZN => n17162);
   U1485 : NAND4_X1 port map( A1 => n17165, A2 => n17164, A3 => n17163, A4 => 
                           n17162, ZN => n17166);
   U1486 : NOR2_X1 port map( A1 => n17167, A2 => n17166, ZN => n17179);
   U1487 : AOI22_X1 port map( A1 => n17724, A2 => REGISTERS_2_23_port, B1 => 
                           n17735, B2 => REGISTERS_7_23_port, ZN => n17171);
   U1488 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_5_23_port, B1 => 
                           n17651, B2 => REGISTERS_3_23_port, ZN => n17170);
   U1489 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_6_23_port, B1 => 
                           n17684, B2 => REGISTERS_1_23_port, ZN => n17169);
   U1490 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_23_port, B1 => 
                           n17685, B2 => REGISTERS_0_23_port, ZN => n17168);
   U1491 : NAND4_X1 port map( A1 => n17171, A2 => n17170, A3 => n17169, A4 => 
                           n17168, ZN => n17177);
   U1492 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_23_port, B1 => 
                           n17731, B2 => REGISTERS_10_23_port, ZN => n17175);
   U1493 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_23_port, B1 => 
                           n17650, B2 => REGISTERS_15_23_port, ZN => n17174);
   U1494 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_14_23_port, B1 => 
                           n17721, B2 => REGISTERS_13_23_port, ZN => n17173);
   U1495 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_23_port, B1 => 
                           n17737, B2 => REGISTERS_8_23_port, ZN => n17172);
   U1496 : NAND4_X1 port map( A1 => n17175, A2 => n17174, A3 => n17173, A4 => 
                           n17172, ZN => n17176);
   U1497 : AOI22_X1 port map( A1 => n17563, A2 => n17177, B1 => n17585, B2 => 
                           n17176, ZN => n17178);
   U1498 : OAI21_X1 port map( B1 => n17749, B2 => n17179, A => n17178, ZN => 
                           N440);
   U1499 : AOI22_X1 port map( A1 => n17697, A2 => REGISTERS_30_22_port, B1 => 
                           n17291, B2 => REGISTERS_23_22_port, ZN => n17183);
   U1500 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_22_port, B1 => 
                           n17542, B2 => REGISTERS_24_22_port, ZN => n17182);
   U1501 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_22_port, B1 => 
                           n17496, B2 => REGISTERS_29_22_port, ZN => n17181);
   U1502 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_22_port, B1 => 
                           n17702, B2 => REGISTERS_20_22_port, ZN => n17180);
   U1503 : NAND4_X1 port map( A1 => n17183, A2 => n17182, A3 => n17181, A4 => 
                           n17180, ZN => n17189);
   U1504 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_22_port, B1 => 
                           n17700, B2 => REGISTERS_31_22_port, ZN => n17187);
   U1505 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_22_port, B1 => 
                           n17671, B2 => REGISTERS_17_22_port, ZN => n17186);
   U1506 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_22_port, B1 => 
                           n17709, B2 => REGISTERS_16_22_port, ZN => n17185);
   U1507 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_22_port, B1 => 
                           n17477, B2 => REGISTERS_19_22_port, ZN => n17184);
   U1508 : NAND4_X1 port map( A1 => n17187, A2 => n17186, A3 => n17185, A4 => 
                           n17184, ZN => n17188);
   U1509 : NOR2_X1 port map( A1 => n17189, A2 => n17188, ZN => n17202);
   U1510 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_22_port, B1 => 
                           n17685, B2 => REGISTERS_0_22_port, ZN => n17194);
   U1511 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_22_port, B1 => 
                           n17678, B2 => REGISTERS_2_22_port, ZN => n17193);
   U1512 : INV_X1 port map( A => n17190, ZN => n17732);
   U1513 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_22_port, B1 => 
                           n17733, B2 => REGISTERS_1_22_port, ZN => n17192);
   U1514 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_22_port, B1 => 
                           n17438, B2 => REGISTERS_7_22_port, ZN => n17191);
   U1515 : NAND4_X1 port map( A1 => n17194, A2 => n17193, A3 => n17192, A4 => 
                           n17191, ZN => n17200);
   U1516 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_22_port, B1 => 
                           n17656, B2 => REGISTERS_12_22_port, ZN => n17198);
   U1517 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_9_22_port, B1 => 
                           n17731, B2 => REGISTERS_10_22_port, ZN => n17197);
   U1518 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_13_22_port, B1 => 
                           n17737, B2 => REGISTERS_8_22_port, ZN => n17196);
   U1519 : AOI22_X1 port map( A1 => n17738, A2 => REGISTERS_11_22_port, B1 => 
                           n17735, B2 => REGISTERS_15_22_port, ZN => n17195);
   U1520 : NAND4_X1 port map( A1 => n17198, A2 => n17197, A3 => n17196, A4 => 
                           n17195, ZN => n17199);
   U1521 : AOI22_X1 port map( A1 => n17563, A2 => n17200, B1 => n17585, B2 => 
                           n17199, ZN => n17201);
   U1522 : OAI21_X1 port map( B1 => n17749, B2 => n17202, A => n17201, ZN => 
                           N439);
   U1523 : AOI22_X1 port map( A1 => n17709, A2 => REGISTERS_16_21_port, B1 => 
                           n17291, B2 => REGISTERS_23_21_port, ZN => n17206);
   U1524 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_21_port, B1 => 
                           n17477, B2 => REGISTERS_19_21_port, ZN => n17205);
   U1525 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_21_port, B1 => 
                           n17638, B2 => REGISTERS_26_21_port, ZN => n17204);
   U1526 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_21_port, B1 => 
                           n17452, B2 => REGISTERS_25_21_port, ZN => n17203);
   U1527 : NAND4_X1 port map( A1 => n17206, A2 => n17205, A3 => n17204, A4 => 
                           n17203, ZN => n17212);
   U1528 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_21_port, B1 => 
                           n17453, B2 => REGISTERS_18_21_port, ZN => n17210);
   U1529 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_21_port, B1 => 
                           n17707, B2 => REGISTERS_24_21_port, ZN => n17209);
   U1530 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_21_port, B1 => 
                           n17699, B2 => REGISTERS_29_21_port, ZN => n17208);
   U1531 : AOI22_X1 port map( A1 => n17697, A2 => REGISTERS_30_21_port, B1 => 
                           n17665, B2 => REGISTERS_31_21_port, ZN => n17207);
   U1532 : NAND4_X1 port map( A1 => n17210, A2 => n17209, A3 => n17208, A4 => 
                           n17207, ZN => n17211);
   U1533 : NOR2_X1 port map( A1 => n17212, A2 => n17211, ZN => n17224);
   U1534 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_21_port, B1 => 
                           n17731, B2 => REGISTERS_2_21_port, ZN => n17216);
   U1535 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_21_port, B1 => 
                           n17650, B2 => REGISTERS_7_21_port, ZN => n17215);
   U1536 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_5_21_port, B1 => 
                           n17738, B2 => REGISTERS_3_21_port, ZN => n17214);
   U1537 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_21_port, B1 => 
                           n17685, B2 => REGISTERS_0_21_port, ZN => n17213);
   U1538 : NAND4_X1 port map( A1 => n17216, A2 => n17215, A3 => n17214, A4 => 
                           n17213, ZN => n17222);
   U1539 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_21_port, B1 => 
                           n17737, B2 => REGISTERS_8_21_port, ZN => n17220);
   U1540 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_21_port, B1 => 
                           n17684, B2 => REGISTERS_9_21_port, ZN => n17219);
   U1541 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_21_port, B1 => 
                           n17678, B2 => REGISTERS_10_21_port, ZN => n17218);
   U1542 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_21_port, B1 => 
                           n17438, B2 => REGISTERS_15_21_port, ZN => n17217);
   U1543 : NAND4_X1 port map( A1 => n17220, A2 => n17219, A3 => n17218, A4 => 
                           n17217, ZN => n17221);
   U1544 : AOI22_X1 port map( A1 => n17563, A2 => n17222, B1 => n17585, B2 => 
                           n17221, ZN => n17223);
   U1545 : OAI21_X1 port map( B1 => n17749, B2 => n17224, A => n17223, ZN => 
                           N438);
   U1546 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_20_port, B1 => 
                           n17665, B2 => REGISTERS_31_20_port, ZN => n17228);
   U1547 : AOI22_X1 port map( A1 => n17477, A2 => REGISTERS_19_20_port, B1 => 
                           n17707, B2 => REGISTERS_24_20_port, ZN => n17227);
   U1548 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_20_port, B1 => 
                           n17453, B2 => REGISTERS_18_20_port, ZN => n17226);
   U1549 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_20_port, B1 => 
                           n17638, B2 => REGISTERS_26_20_port, ZN => n17225);
   U1550 : NAND4_X1 port map( A1 => n17228, A2 => n17227, A3 => n17226, A4 => 
                           n17225, ZN => n17234);
   U1551 : AOI22_X1 port map( A1 => n17709, A2 => REGISTERS_16_20_port, B1 => 
                           n17476, B2 => REGISTERS_30_20_port, ZN => n17232);
   U1552 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_20_port, B1 => 
                           n17702, B2 => REGISTERS_20_20_port, ZN => n17231);
   U1553 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_20_port, B1 => 
                           n17291, B2 => REGISTERS_23_20_port, ZN => n17230);
   U1554 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_20_port, B1 => 
                           n17699, B2 => REGISTERS_29_20_port, ZN => n17229);
   U1555 : NAND4_X1 port map( A1 => n17232, A2 => n17231, A3 => n17230, A4 => 
                           n17229, ZN => n17233);
   U1556 : NOR2_X1 port map( A1 => n17234, A2 => n17233, ZN => n17246);
   U1557 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_6_20_port, B1 => 
                           n17721, B2 => REGISTERS_5_20_port, ZN => n17238);
   U1558 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_1_20_port, B1 => 
                           n17737, B2 => REGISTERS_0_20_port, ZN => n17237);
   U1559 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_20_port, B1 => 
                           n17735, B2 => REGISTERS_7_20_port, ZN => n17236);
   U1560 : AOI22_X1 port map( A1 => n17738, A2 => REGISTERS_3_20_port, B1 => 
                           n17731, B2 => REGISTERS_2_20_port, ZN => n17235);
   U1561 : NAND4_X1 port map( A1 => n17238, A2 => n17237, A3 => n17236, A4 => 
                           n17235, ZN => n17244);
   U1562 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_8_20_port, B1 => 
                           n17678, B2 => REGISTERS_10_20_port, ZN => n17242);
   U1563 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_20_port, B1 => 
                           n17733, B2 => REGISTERS_9_20_port, ZN => n17241);
   U1564 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_20_port, B1 => 
                           n17651, B2 => REGISTERS_11_20_port, ZN => n17240);
   U1565 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_14_20_port, B1 => 
                           n17650, B2 => REGISTERS_15_20_port, ZN => n17239);
   U1566 : NAND4_X1 port map( A1 => n17242, A2 => n17241, A3 => n17240, A4 => 
                           n17239, ZN => n17243);
   U1567 : AOI22_X1 port map( A1 => n17563, A2 => n17244, B1 => n17744, B2 => 
                           n17243, ZN => n17245);
   U1568 : OAI21_X1 port map( B1 => n17749, B2 => n17246, A => n17245, ZN => 
                           N437);
   U1569 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_19_port, B1 => 
                           n17496, B2 => REGISTERS_29_19_port, ZN => n17250);
   U1570 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_19_port, B1 => 
                           n17695, B2 => REGISTERS_23_19_port, ZN => n17249);
   U1571 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_19_port, B1 => 
                           n17613, B2 => REGISTERS_16_19_port, ZN => n17248);
   U1572 : AOI22_X1 port map( A1 => n17701, A2 => REGISTERS_17_19_port, B1 => 
                           n17477, B2 => REGISTERS_19_19_port, ZN => n17247);
   U1573 : NAND4_X1 port map( A1 => n17250, A2 => n17249, A3 => n17248, A4 => 
                           n17247, ZN => n17256);
   U1574 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_19_port, B1 => 
                           n17666, B2 => REGISTERS_21_19_port, ZN => n17254);
   U1575 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_19_port, B1 => 
                           n17476, B2 => REGISTERS_30_19_port, ZN => n17253);
   U1576 : AOI22_X1 port map( A1 => n17698, A2 => REGISTERS_26_19_port, B1 => 
                           n17707, B2 => REGISTERS_24_19_port, ZN => n17252);
   U1577 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_19_port, B1 => 
                           n17665, B2 => REGISTERS_31_19_port, ZN => n17251);
   U1578 : NAND4_X1 port map( A1 => n17254, A2 => n17253, A3 => n17252, A4 => 
                           n17251, ZN => n17255);
   U1579 : NOR2_X1 port map( A1 => n17256, A2 => n17255, ZN => n17268);
   U1580 : CLKBUF_X1 port map( A => n17746, Z => n17587);
   U1581 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_19_port, B1 => 
                           n17731, B2 => REGISTERS_2_19_port, ZN => n17260);
   U1582 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_19_port, B1 => 
                           n17685, B2 => REGISTERS_0_19_port, ZN => n17259);
   U1583 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_19_port, B1 => 
                           n17438, B2 => REGISTERS_7_19_port, ZN => n17258);
   U1584 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_19_port, B1 => 
                           n17738, B2 => REGISTERS_3_19_port, ZN => n17257);
   U1585 : NAND4_X1 port map( A1 => n17260, A2 => n17259, A3 => n17258, A4 => 
                           n17257, ZN => n17266);
   U1586 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_19_port, B1 => 
                           n17721, B2 => REGISTERS_13_19_port, ZN => n17264);
   U1587 : AOI22_X1 port map( A1 => n17724, A2 => REGISTERS_10_19_port, B1 => 
                           n17735, B2 => REGISTERS_15_19_port, ZN => n17263);
   U1588 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_19_port, B1 => 
                           n17684, B2 => REGISTERS_9_19_port, ZN => n17262);
   U1589 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_19_port, B1 => 
                           n17737, B2 => REGISTERS_8_19_port, ZN => n17261);
   U1590 : NAND4_X1 port map( A1 => n17264, A2 => n17263, A3 => n17262, A4 => 
                           n17261, ZN => n17265);
   U1591 : AOI22_X1 port map( A1 => n17587, A2 => n17266, B1 => n17585, B2 => 
                           n17265, ZN => n17267);
   U1592 : OAI21_X1 port map( B1 => n17749, B2 => n17268, A => n17267, ZN => 
                           N436);
   U1593 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_18_port, B1 => 
                           n17496, B2 => REGISTERS_29_18_port, ZN => n17272);
   U1594 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_18_port, B1 => 
                           n17453, B2 => REGISTERS_18_18_port, ZN => n17271);
   U1595 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_18_port, B1 => 
                           n17477, B2 => REGISTERS_19_18_port, ZN => n17270);
   U1596 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_18_port, B1 => 
                           n17452, B2 => REGISTERS_25_18_port, ZN => n17269);
   U1597 : NAND4_X1 port map( A1 => n17272, A2 => n17271, A3 => n17270, A4 => 
                           n17269, ZN => n17278);
   U1598 : AOI22_X1 port map( A1 => n17291, A2 => REGISTERS_23_18_port, B1 => 
                           n17707, B2 => REGISTERS_24_18_port, ZN => n17276);
   U1599 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_18_port, B1 => 
                           n17614, B2 => REGISTERS_27_18_port, ZN => n17275);
   U1600 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_18_port, B1 => 
                           n17665, B2 => REGISTERS_31_18_port, ZN => n17274);
   U1601 : AOI22_X1 port map( A1 => n17701, A2 => REGISTERS_17_18_port, B1 => 
                           n17476, B2 => REGISTERS_30_18_port, ZN => n17273);
   U1602 : NAND4_X1 port map( A1 => n17276, A2 => n17275, A3 => n17274, A4 => 
                           n17273, ZN => n17277);
   U1603 : NOR2_X1 port map( A1 => n17278, A2 => n17277, ZN => n17290);
   U1604 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_18_port, B1 => 
                           n17650, B2 => REGISTERS_7_18_port, ZN => n17282);
   U1605 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_1_18_port, B1 => 
                           n17685, B2 => REGISTERS_0_18_port, ZN => n17281);
   U1606 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_18_port, B1 => 
                           n17651, B2 => REGISTERS_3_18_port, ZN => n17280);
   U1607 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_4_18_port, B1 => 
                           n17678, B2 => REGISTERS_2_18_port, ZN => n17279);
   U1608 : NAND4_X1 port map( A1 => n17282, A2 => n17281, A3 => n17280, A4 => 
                           n17279, ZN => n17288);
   U1609 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_18_port, B1 => 
                           n17733, B2 => REGISTERS_9_18_port, ZN => n17286);
   U1610 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_18_port, B1 => 
                           n17731, B2 => REGISTERS_10_18_port, ZN => n17285);
   U1611 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_18_port, B1 => 
                           n17737, B2 => REGISTERS_8_18_port, ZN => n17284);
   U1612 : AOI22_X1 port map( A1 => n17651, A2 => REGISTERS_11_18_port, B1 => 
                           n17438, B2 => REGISTERS_15_18_port, ZN => n17283);
   U1613 : NAND4_X1 port map( A1 => n17286, A2 => n17285, A3 => n17284, A4 => 
                           n17283, ZN => n17287);
   U1614 : AOI22_X1 port map( A1 => n17587, A2 => n17288, B1 => n17585, B2 => 
                           n17287, ZN => n17289);
   U1615 : OAI21_X1 port map( B1 => n17749, B2 => n17290, A => n17289, ZN => 
                           N435);
   U1616 : AOI22_X1 port map( A1 => n17291, A2 => REGISTERS_23_17_port, B1 => 
                           n17707, B2 => REGISTERS_24_17_port, ZN => n17295);
   U1617 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_17_port, B1 => 
                           n17711, B2 => REGISTERS_18_17_port, ZN => n17294);
   U1618 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_17_port, B1 => 
                           n17665, B2 => REGISTERS_31_17_port, ZN => n17293);
   U1619 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_17_port, B1 => 
                           n17713, B2 => REGISTERS_19_17_port, ZN => n17292);
   U1620 : NAND4_X1 port map( A1 => n17295, A2 => n17294, A3 => n17293, A4 => 
                           n17292, ZN => n17301);
   U1621 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_17_port, B1 => 
                           n17613, B2 => REGISTERS_16_17_port, ZN => n17299);
   U1622 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_17_port, B1 => 
                           n17496, B2 => REGISTERS_29_17_port, ZN => n17298);
   U1623 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_17_port, B1 => 
                           n17638, B2 => REGISTERS_26_17_port, ZN => n17297);
   U1624 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_17_port, B1 => 
                           n17697, B2 => REGISTERS_30_17_port, ZN => n17296);
   U1625 : NAND4_X1 port map( A1 => n17299, A2 => n17298, A3 => n17297, A4 => 
                           n17296, ZN => n17300);
   U1626 : NOR2_X1 port map( A1 => n17301, A2 => n17300, ZN => n17313);
   U1627 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_17_port, B1 => 
                           n17656, B2 => REGISTERS_4_17_port, ZN => n17305);
   U1628 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_17_port, B1 => 
                           n17685, B2 => REGISTERS_0_17_port, ZN => n17304);
   U1629 : AOI22_X1 port map( A1 => n17724, A2 => REGISTERS_2_17_port, B1 => 
                           n17438, B2 => REGISTERS_7_17_port, ZN => n17303);
   U1630 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_1_17_port, B1 => 
                           n17738, B2 => REGISTERS_3_17_port, ZN => n17302);
   U1631 : NAND4_X1 port map( A1 => n17305, A2 => n17304, A3 => n17303, A4 => 
                           n17302, ZN => n17311);
   U1632 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_17_port, B1 => 
                           n17651, B2 => REGISTERS_11_17_port, ZN => n17309);
   U1633 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_17_port, B1 => 
                           n17735, B2 => REGISTERS_15_17_port, ZN => n17308);
   U1634 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_8_17_port, B1 => 
                           n17731, B2 => REGISTERS_10_17_port, ZN => n17307);
   U1635 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_17_port, B1 => 
                           n17656, B2 => REGISTERS_12_17_port, ZN => n17306);
   U1636 : NAND4_X1 port map( A1 => n17309, A2 => n17308, A3 => n17307, A4 => 
                           n17306, ZN => n17310);
   U1637 : AOI22_X1 port map( A1 => n17587, A2 => n17311, B1 => n17585, B2 => 
                           n17310, ZN => n17312);
   U1638 : OAI21_X1 port map( B1 => n17749, B2 => n17313, A => n17312, ZN => 
                           N434);
   U1639 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_16_port, B1 => 
                           n17671, B2 => REGISTERS_17_16_port, ZN => n17317);
   U1640 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_16_port, B1 => 
                           n17452, B2 => REGISTERS_25_16_port, ZN => n17316);
   U1641 : AOI22_X1 port map( A1 => n17477, A2 => REGISTERS_19_16_port, B1 => 
                           n17665, B2 => REGISTERS_31_16_port, ZN => n17315);
   U1642 : AOI22_X1 port map( A1 => n17594, A2 => REGISTERS_28_16_port, B1 => 
                           n17697, B2 => REGISTERS_30_16_port, ZN => n17314);
   U1643 : NAND4_X1 port map( A1 => n17317, A2 => n17316, A3 => n17315, A4 => 
                           n17314, ZN => n17323);
   U1644 : AOI22_X1 port map( A1 => n17695, A2 => REGISTERS_23_16_port, B1 => 
                           n17707, B2 => REGISTERS_24_16_port, ZN => n17321);
   U1645 : AOI22_X1 port map( A1 => n17453, A2 => REGISTERS_18_16_port, B1 => 
                           n17496, B2 => REGISTERS_29_16_port, ZN => n17320);
   U1646 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_16_port, B1 => 
                           n17613, B2 => REGISTERS_16_16_port, ZN => n17319);
   U1647 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_16_port, B1 => 
                           n17698, B2 => REGISTERS_26_16_port, ZN => n17318);
   U1648 : NAND4_X1 port map( A1 => n17321, A2 => n17320, A3 => n17319, A4 => 
                           n17318, ZN => n17322);
   U1649 : NOR2_X1 port map( A1 => n17323, A2 => n17322, ZN => n17335);
   U1650 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_16_port, B1 => 
                           n17684, B2 => REGISTERS_1_16_port, ZN => n17327);
   U1651 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_5_16_port, B1 => 
                           n17738, B2 => REGISTERS_3_16_port, ZN => n17326);
   U1652 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_0_16_port, B1 => 
                           n17650, B2 => REGISTERS_7_16_port, ZN => n17325);
   U1653 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_4_16_port, B1 => 
                           n17724, B2 => REGISTERS_2_16_port, ZN => n17324);
   U1654 : NAND4_X1 port map( A1 => n17327, A2 => n17326, A3 => n17325, A4 => 
                           n17324, ZN => n17333);
   U1655 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_12_16_port, B1 => 
                           n17738, B2 => REGISTERS_11_16_port, ZN => n17331);
   U1656 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_16_port, B1 => 
                           n17731, B2 => REGISTERS_10_16_port, ZN => n17330);
   U1657 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_13_16_port, B1 => 
                           n17735, B2 => REGISTERS_15_16_port, ZN => n17329);
   U1658 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_9_16_port, B1 => 
                           n17737, B2 => REGISTERS_8_16_port, ZN => n17328);
   U1659 : NAND4_X1 port map( A1 => n17331, A2 => n17330, A3 => n17329, A4 => 
                           n17328, ZN => n17332);
   U1660 : AOI22_X1 port map( A1 => n17587, A2 => n17333, B1 => n17585, B2 => 
                           n17332, ZN => n17334);
   U1661 : OAI21_X1 port map( B1 => n17749, B2 => n17335, A => n17334, ZN => 
                           N433);
   U1662 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_15_port, B1 => 
                           n17496, B2 => REGISTERS_29_15_port, ZN => n17339);
   U1663 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_15_port, B1 => 
                           n17713, B2 => REGISTERS_19_15_port, ZN => n17338);
   U1664 : AOI22_X1 port map( A1 => n17452, A2 => REGISTERS_25_15_port, B1 => 
                           n17614, B2 => REGISTERS_27_15_port, ZN => n17337);
   U1665 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_15_port, B1 => 
                           n17594, B2 => REGISTERS_28_15_port, ZN => n17336);
   U1666 : NAND4_X1 port map( A1 => n17339, A2 => n17338, A3 => n17337, A4 => 
                           n17336, ZN => n17345);
   U1667 : AOI22_X1 port map( A1 => n17476, A2 => REGISTERS_30_15_port, B1 => 
                           n17665, B2 => REGISTERS_31_15_port, ZN => n17343);
   U1668 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_15_port, B1 => 
                           n17707, B2 => REGISTERS_24_15_port, ZN => n17342);
   U1669 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_15_port, B1 => 
                           n17695, B2 => REGISTERS_23_15_port, ZN => n17341);
   U1670 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_15_port, B1 => 
                           n17671, B2 => REGISTERS_17_15_port, ZN => n17340);
   U1671 : NAND4_X1 port map( A1 => n17343, A2 => n17342, A3 => n17341, A4 => 
                           n17340, ZN => n17344);
   U1672 : NOR2_X1 port map( A1 => n17345, A2 => n17344, ZN => n17357);
   U1673 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_15_port, B1 => 
                           n17721, B2 => REGISTERS_5_15_port, ZN => n17349);
   U1674 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_15_port, B1 => 
                           n17733, B2 => REGISTERS_1_15_port, ZN => n17348);
   U1675 : AOI22_X1 port map( A1 => n17724, A2 => REGISTERS_2_15_port, B1 => 
                           n17438, B2 => REGISTERS_7_15_port, ZN => n17347);
   U1676 : AOI22_X1 port map( A1 => n17651, A2 => REGISTERS_3_15_port, B1 => 
                           n17722, B2 => REGISTERS_0_15_port, ZN => n17346);
   U1677 : NAND4_X1 port map( A1 => n17349, A2 => n17348, A3 => n17347, A4 => 
                           n17346, ZN => n17355);
   U1678 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_15_port, B1 => 
                           n17735, B2 => REGISTERS_15_15_port, ZN => n17353);
   U1679 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_9_15_port, B1 => 
                           n17651, B2 => REGISTERS_11_15_port, ZN => n17352);
   U1680 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_15_port, B1 => 
                           n17656, B2 => REGISTERS_12_15_port, ZN => n17351);
   U1681 : AOI22_X1 port map( A1 => n17685, A2 => REGISTERS_8_15_port, B1 => 
                           n17678, B2 => REGISTERS_10_15_port, ZN => n17350);
   U1682 : NAND4_X1 port map( A1 => n17353, A2 => n17352, A3 => n17351, A4 => 
                           n17350, ZN => n17354);
   U1683 : AOI22_X1 port map( A1 => n17587, A2 => n17355, B1 => n17585, B2 => 
                           n17354, ZN => n17356);
   U1684 : OAI21_X1 port map( B1 => n17694, B2 => n17357, A => n17356, ZN => 
                           N432);
   U1685 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_14_port, B1 => 
                           n17713, B2 => REGISTERS_19_14_port, ZN => n17361);
   U1686 : AOI22_X1 port map( A1 => n17614, A2 => REGISTERS_27_14_port, B1 => 
                           n17638, B2 => REGISTERS_26_14_port, ZN => n17360);
   U1687 : AOI22_X1 port map( A1 => n17452, A2 => REGISTERS_25_14_port, B1 => 
                           n17695, B2 => REGISTERS_23_14_port, ZN => n17359);
   U1688 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_14_port, B1 => 
                           n17665, B2 => REGISTERS_31_14_port, ZN => n17358);
   U1689 : NAND4_X1 port map( A1 => n17361, A2 => n17360, A3 => n17359, A4 => 
                           n17358, ZN => n17367);
   U1690 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_14_port, B1 => 
                           n17697, B2 => REGISTERS_30_14_port, ZN => n17365);
   U1691 : AOI22_X1 port map( A1 => n17453, A2 => REGISTERS_18_14_port, B1 => 
                           n17496, B2 => REGISTERS_29_14_port, ZN => n17364);
   U1692 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_14_port, B1 => 
                           n17707, B2 => REGISTERS_24_14_port, ZN => n17363);
   U1693 : AOI22_X1 port map( A1 => n17666, A2 => REGISTERS_21_14_port, B1 => 
                           n17594, B2 => REGISTERS_28_14_port, ZN => n17362);
   U1694 : NAND4_X1 port map( A1 => n17365, A2 => n17364, A3 => n17363, A4 => 
                           n17362, ZN => n17366);
   U1695 : NOR2_X1 port map( A1 => n17367, A2 => n17366, ZN => n17379);
   U1696 : AOI22_X1 port map( A1 => n17738, A2 => REGISTERS_3_14_port, B1 => 
                           n17650, B2 => REGISTERS_7_14_port, ZN => n17371);
   U1697 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_14_port, B1 => 
                           n17721, B2 => REGISTERS_5_14_port, ZN => n17370);
   U1698 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_1_14_port, B1 => 
                           n17724, B2 => REGISTERS_2_14_port, ZN => n17369);
   U1699 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_14_port, B1 => 
                           n17722, B2 => REGISTERS_0_14_port, ZN => n17368);
   U1700 : NAND4_X1 port map( A1 => n17371, A2 => n17370, A3 => n17369, A4 => 
                           n17368, ZN => n17377);
   U1701 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_9_14_port, B1 => 
                           n17650, B2 => REGISTERS_15_14_port, ZN => n17375);
   U1702 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_14_14_port, B1 => 
                           n17656, B2 => REGISTERS_12_14_port, ZN => n17374);
   U1703 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_14_port, B1 => 
                           n17737, B2 => REGISTERS_8_14_port, ZN => n17373);
   U1704 : AOI22_X1 port map( A1 => n17651, A2 => REGISTERS_11_14_port, B1 => 
                           n17724, B2 => REGISTERS_10_14_port, ZN => n17372);
   U1705 : NAND4_X1 port map( A1 => n17375, A2 => n17374, A3 => n17373, A4 => 
                           n17372, ZN => n17376);
   U1706 : AOI22_X1 port map( A1 => n17587, A2 => n17377, B1 => n17585, B2 => 
                           n17376, ZN => n17378);
   U1707 : OAI21_X1 port map( B1 => n17749, B2 => n17379, A => n17378, ZN => 
                           N431);
   U1708 : AOI22_X1 port map( A1 => n17666, A2 => REGISTERS_21_13_port, B1 => 
                           n17614, B2 => REGISTERS_27_13_port, ZN => n17383);
   U1709 : AOI22_X1 port map( A1 => n17697, A2 => REGISTERS_30_13_port, B1 => 
                           n17707, B2 => REGISTERS_24_13_port, ZN => n17382);
   U1710 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_13_port, B1 => 
                           n17711, B2 => REGISTERS_18_13_port, ZN => n17381);
   U1711 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_13_port, B1 => 
                           n17665, B2 => REGISTERS_31_13_port, ZN => n17380);
   U1712 : NAND4_X1 port map( A1 => n17383, A2 => n17382, A3 => n17381, A4 => 
                           n17380, ZN => n17389);
   U1713 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_13_port, B1 => 
                           n17594, B2 => REGISTERS_28_13_port, ZN => n17387);
   U1714 : AOI22_X1 port map( A1 => n17695, A2 => REGISTERS_23_13_port, B1 => 
                           n17496, B2 => REGISTERS_29_13_port, ZN => n17386);
   U1715 : AOI22_X1 port map( A1 => n17615, A2 => REGISTERS_20_13_port, B1 => 
                           n17713, B2 => REGISTERS_19_13_port, ZN => n17385);
   U1716 : AOI22_X1 port map( A1 => n17452, A2 => REGISTERS_25_13_port, B1 => 
                           n17638, B2 => REGISTERS_26_13_port, ZN => n17384);
   U1717 : NAND4_X1 port map( A1 => n17387, A2 => n17386, A3 => n17385, A4 => 
                           n17384, ZN => n17388);
   U1718 : NOR2_X1 port map( A1 => n17389, A2 => n17388, ZN => n17401);
   U1719 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_1_13_port, B1 => 
                           n17685, B2 => REGISTERS_0_13_port, ZN => n17393);
   U1720 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_13_port, B1 => 
                           n17438, B2 => REGISTERS_7_13_port, ZN => n17392);
   U1721 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_6_13_port, B1 => 
                           n17678, B2 => REGISTERS_2_13_port, ZN => n17391);
   U1722 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_13_port, B1 => 
                           n17738, B2 => REGISTERS_3_13_port, ZN => n17390);
   U1723 : NAND4_X1 port map( A1 => n17393, A2 => n17392, A3 => n17391, A4 => 
                           n17390, ZN => n17399);
   U1724 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_13_port, B1 => 
                           n17684, B2 => REGISTERS_9_13_port, ZN => n17397);
   U1725 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_13_port, B1 => 
                           n17735, B2 => REGISTERS_15_13_port, ZN => n17396);
   U1726 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_8_13_port, B1 => 
                           n17731, B2 => REGISTERS_10_13_port, ZN => n17395);
   U1727 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_13_port, B1 => 
                           n17656, B2 => REGISTERS_12_13_port, ZN => n17394);
   U1728 : NAND4_X1 port map( A1 => n17397, A2 => n17396, A3 => n17395, A4 => 
                           n17394, ZN => n17398);
   U1729 : AOI22_X1 port map( A1 => n17587, A2 => n17399, B1 => n17585, B2 => 
                           n17398, ZN => n17400);
   U1730 : OAI21_X1 port map( B1 => n17694, B2 => n17401, A => n17400, ZN => 
                           N430);
   U1731 : AOI22_X1 port map( A1 => n17594, A2 => REGISTERS_28_12_port, B1 => 
                           n17697, B2 => REGISTERS_30_12_port, ZN => n17405);
   U1732 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_12_port, B1 => 
                           n17665, B2 => REGISTERS_31_12_port, ZN => n17404);
   U1733 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_12_port, B1 => 
                           n17711, B2 => REGISTERS_18_12_port, ZN => n17403);
   U1734 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_12_port, B1 => 
                           n17695, B2 => REGISTERS_23_12_port, ZN => n17402);
   U1735 : NAND4_X1 port map( A1 => n17405, A2 => n17404, A3 => n17403, A4 => 
                           n17402, ZN => n17411);
   U1736 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_12_port, B1 => 
                           n17614, B2 => REGISTERS_27_12_port, ZN => n17409);
   U1737 : AOI22_X1 port map( A1 => n17615, A2 => REGISTERS_20_12_port, B1 => 
                           n17707, B2 => REGISTERS_24_12_port, ZN => n17408);
   U1738 : AOI22_X1 port map( A1 => n17666, A2 => REGISTERS_21_12_port, B1 => 
                           n17452, B2 => REGISTERS_25_12_port, ZN => n17407);
   U1739 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_12_port, B1 => 
                           n17496, B2 => REGISTERS_29_12_port, ZN => n17406);
   U1740 : NAND4_X1 port map( A1 => n17409, A2 => n17408, A3 => n17407, A4 => 
                           n17406, ZN => n17410);
   U1741 : NOR2_X1 port map( A1 => n17411, A2 => n17410, ZN => n17423);
   U1742 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_4_12_port, B1 => 
                           n17731, B2 => REGISTERS_2_12_port, ZN => n17415);
   U1743 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_12_port, B1 => 
                           n17650, B2 => REGISTERS_7_12_port, ZN => n17414);
   U1744 : AOI22_X1 port map( A1 => n17651, A2 => REGISTERS_3_12_port, B1 => 
                           n17722, B2 => REGISTERS_0_12_port, ZN => n17413);
   U1745 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_12_port, B1 => 
                           n17733, B2 => REGISTERS_1_12_port, ZN => n17412);
   U1746 : NAND4_X1 port map( A1 => n17415, A2 => n17414, A3 => n17413, A4 => 
                           n17412, ZN => n17421);
   U1747 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_12_port, B1 => 
                           n17650, B2 => REGISTERS_15_12_port, ZN => n17419);
   U1748 : AOI22_X1 port map( A1 => n17737, A2 => REGISTERS_8_12_port, B1 => 
                           n17678, B2 => REGISTERS_10_12_port, ZN => n17418);
   U1749 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_14_12_port, B1 => 
                           n17656, B2 => REGISTERS_12_12_port, ZN => n17417);
   U1750 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_9_12_port, B1 => 
                           n17651, B2 => REGISTERS_11_12_port, ZN => n17416);
   U1751 : NAND4_X1 port map( A1 => n17419, A2 => n17418, A3 => n17417, A4 => 
                           n17416, ZN => n17420);
   U1752 : AOI22_X1 port map( A1 => n17587, A2 => n17421, B1 => n17585, B2 => 
                           n17420, ZN => n17422);
   U1753 : OAI21_X1 port map( B1 => n17749, B2 => n17423, A => n17422, ZN => 
                           N429);
   U1754 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_11_port, B1 => 
                           n17496, B2 => REGISTERS_29_11_port, ZN => n17427);
   U1755 : AOI22_X1 port map( A1 => n17614, A2 => REGISTERS_27_11_port, B1 => 
                           n17613, B2 => REGISTERS_16_11_port, ZN => n17426);
   U1756 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_11_port, B1 => 
                           n17671, B2 => REGISTERS_17_11_port, ZN => n17425);
   U1757 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_11_port, B1 => 
                           n17697, B2 => REGISTERS_30_11_port, ZN => n17424);
   U1758 : NAND4_X1 port map( A1 => n17427, A2 => n17426, A3 => n17425, A4 => 
                           n17424, ZN => n17433);
   U1759 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_11_port, B1 => 
                           n17707, B2 => REGISTERS_24_11_port, ZN => n17431);
   U1760 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_11_port, B1 => 
                           n17452, B2 => REGISTERS_25_11_port, ZN => n17430);
   U1761 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_11_port, B1 => 
                           n17665, B2 => REGISTERS_31_11_port, ZN => n17429);
   U1762 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_11_port, B1 => 
                           n17695, B2 => REGISTERS_23_11_port, ZN => n17428);
   U1763 : NAND4_X1 port map( A1 => n17431, A2 => n17430, A3 => n17429, A4 => 
                           n17428, ZN => n17432);
   U1764 : NOR2_X1 port map( A1 => n17433, A2 => n17432, ZN => n17447);
   U1765 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_11_port, B1 => 
                           n17731, B2 => REGISTERS_2_11_port, ZN => n17437);
   U1766 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_11_port, B1 => 
                           n17721, B2 => REGISTERS_5_11_port, ZN => n17436);
   U1767 : AOI22_X1 port map( A1 => n17737, A2 => REGISTERS_0_11_port, B1 => 
                           n17650, B2 => REGISTERS_7_11_port, ZN => n17435);
   U1768 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_11_port, B1 => 
                           n17738, B2 => REGISTERS_3_11_port, ZN => n17434);
   U1769 : NAND4_X1 port map( A1 => n17437, A2 => n17436, A3 => n17435, A4 => 
                           n17434, ZN => n17445);
   U1770 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_11_port, B1 => 
                           n17438, B2 => REGISTERS_15_11_port, ZN => n17443);
   U1771 : AOI22_X1 port map( A1 => n17439, A2 => REGISTERS_14_11_port, B1 => 
                           n17656, B2 => REGISTERS_12_11_port, ZN => n17442);
   U1772 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_11_port, B1 => 
                           n17722, B2 => REGISTERS_8_11_port, ZN => n17441);
   U1773 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_9_11_port, B1 => 
                           n17678, B2 => REGISTERS_10_11_port, ZN => n17440);
   U1774 : NAND4_X1 port map( A1 => n17443, A2 => n17442, A3 => n17441, A4 => 
                           n17440, ZN => n17444);
   U1775 : AOI22_X1 port map( A1 => n17587, A2 => n17445, B1 => n17585, B2 => 
                           n17444, ZN => n17446);
   U1776 : OAI21_X1 port map( B1 => n17749, B2 => n17447, A => n17446, ZN => 
                           N428);
   U1777 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_10_port, B1 => 
                           n17695, B2 => REGISTERS_23_10_port, ZN => n17451);
   U1778 : AOI22_X1 port map( A1 => n17542, A2 => REGISTERS_24_10_port, B1 => 
                           n17496, B2 => REGISTERS_29_10_port, ZN => n17450);
   U1779 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_10_port, B1 => 
                           n17614, B2 => REGISTERS_27_10_port, ZN => n17449);
   U1780 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_10_port, B1 => 
                           n17697, B2 => REGISTERS_30_10_port, ZN => n17448);
   U1781 : NAND4_X1 port map( A1 => n17451, A2 => n17450, A3 => n17449, A4 => 
                           n17448, ZN => n17459);
   U1782 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_10_port, B1 => 
                           n17671, B2 => REGISTERS_17_10_port, ZN => n17457);
   U1783 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_10_port, B1 => 
                           n17452, B2 => REGISTERS_25_10_port, ZN => n17456);
   U1784 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_10_port, B1 => 
                           n17713, B2 => REGISTERS_19_10_port, ZN => n17455);
   U1785 : AOI22_X1 port map( A1 => n17453, A2 => REGISTERS_18_10_port, B1 => 
                           n17665, B2 => REGISTERS_31_10_port, ZN => n17454);
   U1786 : NAND4_X1 port map( A1 => n17457, A2 => n17456, A3 => n17455, A4 => 
                           n17454, ZN => n17458);
   U1787 : NOR2_X1 port map( A1 => n17459, A2 => n17458, ZN => n17471);
   U1788 : AOI22_X1 port map( A1 => n17738, A2 => REGISTERS_3_10_port, B1 => 
                           n17735, B2 => REGISTERS_7_10_port, ZN => n17463);
   U1789 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_10_port, B1 => 
                           n17724, B2 => REGISTERS_2_10_port, ZN => n17462);
   U1790 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_10_port, B1 => 
                           n17684, B2 => REGISTERS_1_10_port, ZN => n17461);
   U1791 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_6_10_port, B1 => 
                           n17737, B2 => REGISTERS_0_10_port, ZN => n17460);
   U1792 : NAND4_X1 port map( A1 => n17463, A2 => n17462, A3 => n17461, A4 => 
                           n17460, ZN => n17469);
   U1793 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_14_10_port, B1 => 
                           n17724, B2 => REGISTERS_10_10_port, ZN => n17467);
   U1794 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_10_port, B1 => 
                           n17650, B2 => REGISTERS_15_10_port, ZN => n17466);
   U1795 : AOI22_X1 port map( A1 => n17738, A2 => REGISTERS_11_10_port, B1 => 
                           n17737, B2 => REGISTERS_8_10_port, ZN => n17465);
   U1796 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_10_port, B1 => 
                           n17733, B2 => REGISTERS_9_10_port, ZN => n17464);
   U1797 : NAND4_X1 port map( A1 => n17467, A2 => n17466, A3 => n17465, A4 => 
                           n17464, ZN => n17468);
   U1798 : AOI22_X1 port map( A1 => n17587, A2 => n17469, B1 => n17585, B2 => 
                           n17468, ZN => n17470);
   U1799 : OAI21_X1 port map( B1 => n17749, B2 => n17471, A => n17470, ZN => 
                           N427);
   U1800 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_9_port, B1 => 
                           n17701, B2 => REGISTERS_17_9_port, ZN => n17475);
   U1801 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_9_port, B1 => 
                           n17613, B2 => REGISTERS_16_9_port, ZN => n17474);
   U1802 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_9_port, B1 => 
                           n17496, B2 => REGISTERS_29_9_port, ZN => n17473);
   U1803 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_9_port, B1 => 
                           n17711, B2 => REGISTERS_18_9_port, ZN => n17472);
   U1804 : NAND4_X1 port map( A1 => n17475, A2 => n17474, A3 => n17473, A4 => 
                           n17472, ZN => n17483);
   U1805 : AOI22_X1 port map( A1 => n17476, A2 => REGISTERS_30_9_port, B1 => 
                           n17695, B2 => REGISTERS_23_9_port, ZN => n17481);
   U1806 : AOI22_X1 port map( A1 => n17477, A2 => REGISTERS_19_9_port, B1 => 
                           n17665, B2 => REGISTERS_31_9_port, ZN => n17480);
   U1807 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_9_port, B1 => 
                           n17615, B2 => REGISTERS_20_9_port, ZN => n17479);
   U1808 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_9_port, B1 => 
                           n17707, B2 => REGISTERS_24_9_port, ZN => n17478);
   U1809 : NAND4_X1 port map( A1 => n17481, A2 => n17480, A3 => n17479, A4 => 
                           n17478, ZN => n17482);
   U1810 : NOR2_X1 port map( A1 => n17483, A2 => n17482, ZN => n17495);
   U1811 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_1_9_port, B1 => 
                           n17726, B2 => REGISTERS_3_9_port, ZN => n17487);
   U1812 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_4_9_port, B1 => 
                           n17724, B2 => REGISTERS_2_9_port, ZN => n17486);
   U1813 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_9_port, B1 => 
                           n17737, B2 => REGISTERS_0_9_port, ZN => n17485);
   U1814 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_6_9_port, B1 => 
                           n17735, B2 => REGISTERS_7_9_port, ZN => n17484);
   U1815 : NAND4_X1 port map( A1 => n17487, A2 => n17486, A3 => n17485, A4 => 
                           n17484, ZN => n17493);
   U1816 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_9_9_port, B1 => 
                           n17738, B2 => REGISTERS_11_9_port, ZN => n17491);
   U1817 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_9_port, B1 => 
                           n17678, B2 => REGISTERS_10_9_port, ZN => n17490);
   U1818 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_14_9_port, B1 => 
                           n17722, B2 => REGISTERS_8_9_port, ZN => n17489);
   U1819 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_9_port, B1 => 
                           n17650, B2 => REGISTERS_15_9_port, ZN => n17488);
   U1820 : NAND4_X1 port map( A1 => n17491, A2 => n17490, A3 => n17489, A4 => 
                           n17488, ZN => n17492);
   U1821 : AOI22_X1 port map( A1 => n17587, A2 => n17493, B1 => n17585, B2 => 
                           n17492, ZN => n17494);
   U1822 : OAI21_X1 port map( B1 => n17694, B2 => n17495, A => n17494, ZN => 
                           N426);
   U1823 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_8_port, B1 => 
                           n17615, B2 => REGISTERS_20_8_port, ZN => n17501);
   U1824 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_8_port, B1 => 
                           n17496, B2 => REGISTERS_29_8_port, ZN => n17500);
   U1825 : AOI22_X1 port map( A1 => n17497, A2 => REGISTERS_22_8_port, B1 => 
                           n17711, B2 => REGISTERS_18_8_port, ZN => n17499);
   U1826 : AOI22_X1 port map( A1 => n17709, A2 => REGISTERS_16_8_port, B1 => 
                           n17665, B2 => REGISTERS_31_8_port, ZN => n17498);
   U1827 : NAND4_X1 port map( A1 => n17501, A2 => n17500, A3 => n17499, A4 => 
                           n17498, ZN => n17507);
   U1828 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_8_port, B1 => 
                           n17713, B2 => REGISTERS_19_8_port, ZN => n17505);
   U1829 : AOI22_X1 port map( A1 => n17701, A2 => REGISTERS_17_8_port, B1 => 
                           n17695, B2 => REGISTERS_23_8_port, ZN => n17504);
   U1830 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_8_port, B1 => 
                           n17697, B2 => REGISTERS_30_8_port, ZN => n17503);
   U1831 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_8_port, B1 => 
                           n17707, B2 => REGISTERS_24_8_port, ZN => n17502);
   U1832 : NAND4_X1 port map( A1 => n17505, A2 => n17504, A3 => n17503, A4 => 
                           n17502, ZN => n17506);
   U1833 : NOR2_X1 port map( A1 => n17507, A2 => n17506, ZN => n17519);
   U1834 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_8_port, B1 => 
                           n17651, B2 => REGISTERS_3_8_port, ZN => n17511);
   U1835 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_1_8_port, B1 => 
                           n17735, B2 => REGISTERS_7_8_port, ZN => n17510);
   U1836 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_6_8_port, B1 => 
                           n17685, B2 => REGISTERS_0_8_port, ZN => n17509);
   U1837 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_8_port, B1 => 
                           n17731, B2 => REGISTERS_2_8_port, ZN => n17508);
   U1838 : NAND4_X1 port map( A1 => n17511, A2 => n17510, A3 => n17509, A4 => 
                           n17508, ZN => n17517);
   U1839 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_12_8_port, B1 => 
                           n17651, B2 => REGISTERS_11_8_port, ZN => n17515);
   U1840 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_14_8_port, B1 => 
                           n17650, B2 => REGISTERS_15_8_port, ZN => n17514);
   U1841 : AOI22_X1 port map( A1 => n17685, A2 => REGISTERS_8_8_port, B1 => 
                           n17731, B2 => REGISTERS_10_8_port, ZN => n17513);
   U1842 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_8_port, B1 => 
                           n17733, B2 => REGISTERS_9_8_port, ZN => n17512);
   U1843 : NAND4_X1 port map( A1 => n17515, A2 => n17514, A3 => n17513, A4 => 
                           n17512, ZN => n17516);
   U1844 : AOI22_X1 port map( A1 => n17587, A2 => n17517, B1 => n17585, B2 => 
                           n17516, ZN => n17518);
   U1845 : OAI21_X1 port map( B1 => n17749, B2 => n17519, A => n17518, ZN => 
                           N425);
   U1846 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_7_port, B1 => 
                           n17665, B2 => REGISTERS_31_7_port, ZN => n17523);
   U1847 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_7_port, B1 => 
                           n17698, B2 => REGISTERS_26_7_port, ZN => n17522);
   U1848 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_7_port, B1 => 
                           n17695, B2 => REGISTERS_23_7_port, ZN => n17521);
   U1849 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_7_port, B1 => 
                           n17707, B2 => REGISTERS_24_7_port, ZN => n17520);
   U1850 : NAND4_X1 port map( A1 => n17523, A2 => n17522, A3 => n17521, A4 => 
                           n17520, ZN => n17529);
   U1851 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_7_port, B1 => 
                           n17697, B2 => REGISTERS_30_7_port, ZN => n17527);
   U1852 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_7_port, B1 => 
                           n17711, B2 => REGISTERS_18_7_port, ZN => n17526);
   U1853 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_7_port, B1 => 
                           n17594, B2 => REGISTERS_28_7_port, ZN => n17525);
   U1854 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_7_port, B1 => 
                           n17699, B2 => REGISTERS_29_7_port, ZN => n17524);
   U1855 : NAND4_X1 port map( A1 => n17527, A2 => n17526, A3 => n17525, A4 => 
                           n17524, ZN => n17528);
   U1856 : NOR2_X1 port map( A1 => n17529, A2 => n17528, ZN => n17541);
   U1857 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_7_port, B1 => 
                           n17724, B2 => REGISTERS_2_7_port, ZN => n17533);
   U1858 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_1_7_port, B1 => 
                           n17726, B2 => REGISTERS_3_7_port, ZN => n17532);
   U1859 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_7_port, B1 => 
                           n17685, B2 => REGISTERS_0_7_port, ZN => n17531);
   U1860 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_7_port, B1 => 
                           n17650, B2 => REGISTERS_7_7_port, ZN => n17530);
   U1861 : NAND4_X1 port map( A1 => n17533, A2 => n17532, A3 => n17531, A4 => 
                           n17530, ZN => n17539);
   U1862 : AOI22_X1 port map( A1 => n17737, A2 => REGISTERS_8_7_port, B1 => 
                           n17735, B2 => REGISTERS_15_7_port, ZN => n17537);
   U1863 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_9_7_port, B1 => 
                           n17724, B2 => REGISTERS_10_7_port, ZN => n17536);
   U1864 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_12_7_port, B1 => 
                           n17726, B2 => REGISTERS_11_7_port, ZN => n17535);
   U1865 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_7_port, B1 => 
                           n17679, B2 => REGISTERS_13_7_port, ZN => n17534);
   U1866 : NAND4_X1 port map( A1 => n17537, A2 => n17536, A3 => n17535, A4 => 
                           n17534, ZN => n17538);
   U1867 : AOI22_X1 port map( A1 => n17587, A2 => n17539, B1 => n17585, B2 => 
                           n17538, ZN => n17540);
   U1868 : OAI21_X1 port map( B1 => n17694, B2 => n17541, A => n17540, ZN => 
                           N424);
   U1869 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_6_port, B1 => 
                           n17709, B2 => REGISTERS_16_6_port, ZN => n17546);
   U1870 : AOI22_X1 port map( A1 => n17542, A2 => REGISTERS_24_6_port, B1 => 
                           n17699, B2 => REGISTERS_29_6_port, ZN => n17545);
   U1871 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_6_port, B1 => 
                           n17711, B2 => REGISTERS_18_6_port, ZN => n17544);
   U1872 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_6_port, B1 => 
                           n17698, B2 => REGISTERS_26_6_port, ZN => n17543);
   U1873 : NAND4_X1 port map( A1 => n17546, A2 => n17545, A3 => n17544, A4 => 
                           n17543, ZN => n17552);
   U1874 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_6_port, B1 => 
                           n17665, B2 => REGISTERS_31_6_port, ZN => n17550);
   U1875 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_6_port, B1 => 
                           n17695, B2 => REGISTERS_23_6_port, ZN => n17549);
   U1876 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_6_port, B1 => 
                           n17697, B2 => REGISTERS_30_6_port, ZN => n17548);
   U1877 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_6_port, B1 => 
                           n17666, B2 => REGISTERS_21_6_port, ZN => n17547);
   U1878 : NAND4_X1 port map( A1 => n17550, A2 => n17549, A3 => n17548, A4 => 
                           n17547, ZN => n17551);
   U1879 : NOR2_X1 port map( A1 => n17552, A2 => n17551, ZN => n17565);
   U1880 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_6_port, B1 => 
                           n17650, B2 => REGISTERS_7_6_port, ZN => n17556);
   U1881 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_6_port, B1 => 
                           n17721, B2 => REGISTERS_5_6_port, ZN => n17555);
   U1882 : AOI22_X1 port map( A1 => n17651, A2 => REGISTERS_3_6_port, B1 => 
                           n17737, B2 => REGISTERS_0_6_port, ZN => n17554);
   U1883 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_4_6_port, B1 => 
                           n17678, B2 => REGISTERS_2_6_port, ZN => n17553);
   U1884 : NAND4_X1 port map( A1 => n17556, A2 => n17555, A3 => n17554, A4 => 
                           n17553, ZN => n17562);
   U1885 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_6_port, B1 => 
                           n17731, B2 => REGISTERS_10_6_port, ZN => n17560);
   U1886 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_13_6_port, B1 => 
                           n17684, B2 => REGISTERS_9_6_port, ZN => n17559);
   U1887 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_6_port, B1 => 
                           n17685, B2 => REGISTERS_8_6_port, ZN => n17558);
   U1888 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_6_port, B1 => 
                           n17735, B2 => REGISTERS_15_6_port, ZN => n17557);
   U1889 : NAND4_X1 port map( A1 => n17560, A2 => n17559, A3 => n17558, A4 => 
                           n17557, ZN => n17561);
   U1890 : AOI22_X1 port map( A1 => n17563, A2 => n17562, B1 => n17585, B2 => 
                           n17561, ZN => n17564);
   U1891 : OAI21_X1 port map( B1 => n17749, B2 => n17565, A => n17564, ZN => 
                           N423);
   U1892 : AOI22_X1 port map( A1 => n17700, A2 => REGISTERS_31_5_port, B1 => 
                           n17699, B2 => REGISTERS_29_5_port, ZN => n17569);
   U1893 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_5_port, B1 => 
                           n17707, B2 => REGISTERS_24_5_port, ZN => n17568);
   U1894 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_5_port, B1 => 
                           n17697, B2 => REGISTERS_30_5_port, ZN => n17567);
   U1895 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_5_port, B1 => 
                           n17711, B2 => REGISTERS_18_5_port, ZN => n17566);
   U1896 : NAND4_X1 port map( A1 => n17569, A2 => n17568, A3 => n17567, A4 => 
                           n17566, ZN => n17575);
   U1897 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_5_port, B1 => 
                           n17698, B2 => REGISTERS_26_5_port, ZN => n17573);
   U1898 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_5_port, B1 => 
                           n17695, B2 => REGISTERS_23_5_port, ZN => n17572);
   U1899 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_5_port, B1 => 
                           n17594, B2 => REGISTERS_28_5_port, ZN => n17571);
   U1900 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_5_port, B1 => 
                           n17701, B2 => REGISTERS_17_5_port, ZN => n17570);
   U1901 : NAND4_X1 port map( A1 => n17573, A2 => n17572, A3 => n17571, A4 => 
                           n17570, ZN => n17574);
   U1902 : NOR2_X1 port map( A1 => n17575, A2 => n17574, ZN => n17589);
   U1903 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_5_port, B1 => 
                           n17684, B2 => REGISTERS_1_5_port, ZN => n17579);
   U1904 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_5_port, B1 => 
                           n17685, B2 => REGISTERS_0_5_port, ZN => n17578);
   U1905 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_5_port, B1 => 
                           n17731, B2 => REGISTERS_2_5_port, ZN => n17577);
   U1906 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_5_port, B1 => 
                           n17650, B2 => REGISTERS_7_5_port, ZN => n17576);
   U1907 : NAND4_X1 port map( A1 => n17579, A2 => n17578, A3 => n17577, A4 => 
                           n17576, ZN => n17586);
   U1908 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_5_port, B1 => 
                           n17723, B2 => REGISTERS_9_5_port, ZN => n17583);
   U1909 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_5_port, B1 => 
                           n17738, B2 => REGISTERS_11_5_port, ZN => n17582);
   U1910 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_8_5_port, B1 => 
                           n17724, B2 => REGISTERS_10_5_port, ZN => n17581);
   U1911 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_12_5_port, B1 => 
                           n17735, B2 => REGISTERS_15_5_port, ZN => n17580);
   U1912 : NAND4_X1 port map( A1 => n17583, A2 => n17582, A3 => n17581, A4 => 
                           n17580, ZN => n17584);
   U1913 : AOI22_X1 port map( A1 => n17587, A2 => n17586, B1 => n17585, B2 => 
                           n17584, ZN => n17588);
   U1914 : OAI21_X1 port map( B1 => n17694, B2 => n17589, A => n17588, ZN => 
                           N422);
   U1915 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_4_port, B1 => 
                           n17713, B2 => REGISTERS_19_4_port, ZN => n17593);
   U1916 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_4_port, B1 => 
                           n17665, B2 => REGISTERS_31_4_port, ZN => n17592);
   U1917 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_4_port, B1 => 
                           n17709, B2 => REGISTERS_16_4_port, ZN => n17591);
   U1918 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_4_port, B1 => 
                           n17695, B2 => REGISTERS_23_4_port, ZN => n17590);
   U1919 : NAND4_X1 port map( A1 => n17593, A2 => n17592, A3 => n17591, A4 => 
                           n17590, ZN => n17600);
   U1920 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_4_port, B1 => 
                           n17594, B2 => REGISTERS_28_4_port, ZN => n17598);
   U1921 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_4_port, B1 => 
                           n17699, B2 => REGISTERS_29_4_port, ZN => n17597);
   U1922 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_4_port, B1 => 
                           n17697, B2 => REGISTERS_30_4_port, ZN => n17596);
   U1923 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_4_port, B1 => 
                           n17707, B2 => REGISTERS_24_4_port, ZN => n17595);
   U1924 : NAND4_X1 port map( A1 => n17598, A2 => n17597, A3 => n17596, A4 => 
                           n17595, ZN => n17599);
   U1925 : NOR2_X1 port map( A1 => n17600, A2 => n17599, ZN => n17612);
   U1926 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_0_4_port, B1 => 
                           n17678, B2 => REGISTERS_2_4_port, ZN => n17604);
   U1927 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_4_port, B1 => 
                           n17650, B2 => REGISTERS_7_4_port, ZN => n17603);
   U1928 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_4_port, B1 => 
                           n17723, B2 => REGISTERS_1_4_port, ZN => n17602);
   U1929 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_4_port, B1 => 
                           n17656, B2 => REGISTERS_4_4_port, ZN => n17601);
   U1930 : NAND4_X1 port map( A1 => n17604, A2 => n17603, A3 => n17602, A4 => 
                           n17601, ZN => n17610);
   U1931 : AOI22_X1 port map( A1 => n17733, A2 => REGISTERS_9_4_port, B1 => 
                           n17735, B2 => REGISTERS_15_4_port, ZN => n17608);
   U1932 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_4_port, B1 => 
                           n17656, B2 => REGISTERS_12_4_port, ZN => n17607);
   U1933 : AOI22_X1 port map( A1 => n17738, A2 => REGISTERS_11_4_port, B1 => 
                           n17737, B2 => REGISTERS_8_4_port, ZN => n17606);
   U1934 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_4_port, B1 => 
                           n17724, B2 => REGISTERS_10_4_port, ZN => n17605);
   U1935 : NAND4_X1 port map( A1 => n17608, A2 => n17607, A3 => n17606, A4 => 
                           n17605, ZN => n17609);
   U1936 : AOI22_X1 port map( A1 => n17746, A2 => n17610, B1 => n17744, B2 => 
                           n17609, ZN => n17611);
   U1937 : OAI21_X1 port map( B1 => n17749, B2 => n17612, A => n17611, ZN => 
                           N421);
   U1938 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_3_port, B1 => 
                           n17697, B2 => REGISTERS_30_3_port, ZN => n17619);
   U1939 : AOI22_X1 port map( A1 => n17613, A2 => REGISTERS_16_3_port, B1 => 
                           n17698, B2 => REGISTERS_26_3_port, ZN => n17618);
   U1940 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_3_port, B1 => 
                           n17614, B2 => REGISTERS_27_3_port, ZN => n17617);
   U1941 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_3_port, B1 => 
                           n17615, B2 => REGISTERS_20_3_port, ZN => n17616);
   U1942 : NAND4_X1 port map( A1 => n17619, A2 => n17618, A3 => n17617, A4 => 
                           n17616, ZN => n17625);
   U1943 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_3_port, B1 => 
                           n17707, B2 => REGISTERS_24_3_port, ZN => n17623);
   U1944 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_3_port, B1 => 
                           n17699, B2 => REGISTERS_29_3_port, ZN => n17622);
   U1945 : AOI22_X1 port map( A1 => n17695, A2 => REGISTERS_23_3_port, B1 => 
                           n17665, B2 => REGISTERS_31_3_port, ZN => n17621);
   U1946 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_3_port, B1 => 
                           n17711, B2 => REGISTERS_18_3_port, ZN => n17620);
   U1947 : NAND4_X1 port map( A1 => n17623, A2 => n17622, A3 => n17621, A4 => 
                           n17620, ZN => n17624);
   U1948 : NOR2_X1 port map( A1 => n17625, A2 => n17624, ZN => n17637);
   U1949 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_3_port, B1 => 
                           n17650, B2 => REGISTERS_7_3_port, ZN => n17629);
   U1950 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_4_3_port, B1 => 
                           n17685, B2 => REGISTERS_0_3_port, ZN => n17628);
   U1951 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_3_3_port, B1 => 
                           n17724, B2 => REGISTERS_2_3_port, ZN => n17627);
   U1952 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_5_3_port, B1 => 
                           n17733, B2 => REGISTERS_1_3_port, ZN => n17626);
   U1953 : NAND4_X1 port map( A1 => n17629, A2 => n17628, A3 => n17627, A4 => 
                           n17626, ZN => n17635);
   U1954 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_9_3_port, B1 => 
                           n17726, B2 => REGISTERS_11_3_port, ZN => n17633);
   U1955 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_3_port, B1 => 
                           n17724, B2 => REGISTERS_10_3_port, ZN => n17632);
   U1956 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_8_3_port, B1 => 
                           n17735, B2 => REGISTERS_15_3_port, ZN => n17631);
   U1957 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_13_3_port, B1 => 
                           n17736, B2 => REGISTERS_12_3_port, ZN => n17630);
   U1958 : NAND4_X1 port map( A1 => n17633, A2 => n17632, A3 => n17631, A4 => 
                           n17630, ZN => n17634);
   U1959 : AOI22_X1 port map( A1 => n17746, A2 => n17635, B1 => n17744, B2 => 
                           n17634, ZN => n17636);
   U1960 : OAI21_X1 port map( B1 => n17694, B2 => n17637, A => n17636, ZN => 
                           N420);
   U1961 : AOI22_X1 port map( A1 => n17711, A2 => REGISTERS_18_2_port, B1 => 
                           n17665, B2 => REGISTERS_31_2_port, ZN => n17642);
   U1962 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_2_port, B1 => 
                           n17699, B2 => REGISTERS_29_2_port, ZN => n17641);
   U1963 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_2_port, B1 => 
                           n17713, B2 => REGISTERS_19_2_port, ZN => n17640);
   U1964 : AOI22_X1 port map( A1 => n17638, A2 => REGISTERS_26_2_port, B1 => 
                           n17707, B2 => REGISTERS_24_2_port, ZN => n17639);
   U1965 : NAND4_X1 port map( A1 => n17642, A2 => n17641, A3 => n17640, A4 => 
                           n17639, ZN => n17648);
   U1966 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_2_port, B1 => 
                           n17695, B2 => REGISTERS_23_2_port, ZN => n17646);
   U1967 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_2_port, B1 => 
                           n17701, B2 => REGISTERS_17_2_port, ZN => n17645);
   U1968 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_2_port, B1 => 
                           n17697, B2 => REGISTERS_30_2_port, ZN => n17644);
   U1969 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_2_port, B1 => 
                           n17709, B2 => REGISTERS_16_2_port, ZN => n17643);
   U1970 : NAND4_X1 port map( A1 => n17646, A2 => n17645, A3 => n17644, A4 => 
                           n17643, ZN => n17647);
   U1971 : NOR2_X1 port map( A1 => n17648, A2 => n17647, ZN => n17664);
   U1972 : AOI22_X1 port map( A1 => n17649, A2 => REGISTERS_6_2_port, B1 => 
                           n17733, B2 => REGISTERS_1_2_port, ZN => n17655);
   U1973 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_5_2_port, B1 => 
                           n17650, B2 => REGISTERS_7_2_port, ZN => n17654);
   U1974 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_0_2_port, B1 => 
                           n17678, B2 => REGISTERS_2_2_port, ZN => n17653);
   U1975 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_2_port, B1 => 
                           n17651, B2 => REGISTERS_3_2_port, ZN => n17652);
   U1976 : NAND4_X1 port map( A1 => n17655, A2 => n17654, A3 => n17653, A4 => 
                           n17652, ZN => n17662);
   U1977 : AOI22_X1 port map( A1 => n17684, A2 => REGISTERS_9_2_port, B1 => 
                           n17735, B2 => REGISTERS_15_2_port, ZN => n17660);
   U1978 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_13_2_port, B1 => 
                           n17724, B2 => REGISTERS_10_2_port, ZN => n17659);
   U1979 : AOI22_X1 port map( A1 => n17656, A2 => REGISTERS_12_2_port, B1 => 
                           n17738, B2 => REGISTERS_11_2_port, ZN => n17658);
   U1980 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_2_port, B1 => 
                           n17722, B2 => REGISTERS_8_2_port, ZN => n17657);
   U1981 : NAND4_X1 port map( A1 => n17660, A2 => n17659, A3 => n17658, A4 => 
                           n17657, ZN => n17661);
   U1982 : AOI22_X1 port map( A1 => n17746, A2 => n17662, B1 => n17744, B2 => 
                           n17661, ZN => n17663);
   U1983 : OAI21_X1 port map( B1 => n17749, B2 => n17664, A => n17663, ZN => 
                           N419);
   U1984 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_1_port, B1 => 
                           n17698, B2 => REGISTERS_26_1_port, ZN => n17670);
   U1985 : AOI22_X1 port map( A1 => n17713, A2 => REGISTERS_19_1_port, B1 => 
                           n17707, B2 => REGISTERS_24_1_port, ZN => n17669);
   U1986 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_1_port, B1 => 
                           n17665, B2 => REGISTERS_31_1_port, ZN => n17668);
   U1987 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_1_port, B1 => 
                           n17666, B2 => REGISTERS_21_1_port, ZN => n17667);
   U1988 : NAND4_X1 port map( A1 => n17670, A2 => n17669, A3 => n17668, A4 => 
                           n17667, ZN => n17677);
   U1989 : AOI22_X1 port map( A1 => n17671, A2 => REGISTERS_17_1_port, B1 => 
                           n17711, B2 => REGISTERS_18_1_port, ZN => n17675);
   U1990 : AOI22_X1 port map( A1 => n17697, A2 => REGISTERS_30_1_port, B1 => 
                           n17695, B2 => REGISTERS_23_1_port, ZN => n17674);
   U1991 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_1_port, B1 => 
                           n17709, B2 => REGISTERS_16_1_port, ZN => n17673);
   U1992 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_1_port, B1 => 
                           n17699, B2 => REGISTERS_29_1_port, ZN => n17672);
   U1993 : NAND4_X1 port map( A1 => n17675, A2 => n17674, A3 => n17673, A4 => 
                           n17672, ZN => n17676);
   U1994 : NOR2_X1 port map( A1 => n17677, A2 => n17676, ZN => n17693);
   U1995 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_6_1_port, B1 => 
                           n17736, B2 => REGISTERS_4_1_port, ZN => n17683);
   U1996 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_1_port, B1 => 
                           n17735, B2 => REGISTERS_7_1_port, ZN => n17682);
   U1997 : AOI22_X1 port map( A1 => n17722, A2 => REGISTERS_0_1_port, B1 => 
                           n17678, B2 => REGISTERS_2_1_port, ZN => n17681);
   U1998 : AOI22_X1 port map( A1 => n17679, A2 => REGISTERS_5_1_port, B1 => 
                           n17738, B2 => REGISTERS_3_1_port, ZN => n17680);
   U1999 : NAND4_X1 port map( A1 => n17683, A2 => n17682, A3 => n17681, A4 => 
                           n17680, ZN => n17691);
   U2000 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_1_port, B1 => 
                           n17724, B2 => REGISTERS_10_1_port, ZN => n17689);
   U2001 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_1_port, B1 => 
                           n17735, B2 => REGISTERS_15_1_port, ZN => n17688);
   U2002 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_1_port, B1 => 
                           n17684, B2 => REGISTERS_9_1_port, ZN => n17687);
   U2003 : AOI22_X1 port map( A1 => n17726, A2 => REGISTERS_11_1_port, B1 => 
                           n17685, B2 => REGISTERS_8_1_port, ZN => n17686);
   U2004 : NAND4_X1 port map( A1 => n17689, A2 => n17688, A3 => n17687, A4 => 
                           n17686, ZN => n17690);
   U2005 : AOI22_X1 port map( A1 => n17746, A2 => n17691, B1 => n17744, B2 => 
                           n17690, ZN => n17692);
   U2006 : OAI21_X1 port map( B1 => n17694, B2 => n17693, A => n17692, ZN => 
                           N418);
   U2007 : AOI22_X1 port map( A1 => n17696, A2 => REGISTERS_27_0_port, B1 => 
                           n17695, B2 => REGISTERS_23_0_port, ZN => n17706);
   U2008 : AOI22_X1 port map( A1 => n17698, A2 => REGISTERS_26_0_port, B1 => 
                           n17697, B2 => REGISTERS_30_0_port, ZN => n17705);
   U2009 : AOI22_X1 port map( A1 => n17700, A2 => REGISTERS_31_0_port, B1 => 
                           n17699, B2 => REGISTERS_29_0_port, ZN => n17704);
   U2010 : AOI22_X1 port map( A1 => n17702, A2 => REGISTERS_20_0_port, B1 => 
                           n17701, B2 => REGISTERS_17_0_port, ZN => n17703);
   U2011 : NAND4_X1 port map( A1 => n17706, A2 => n17705, A3 => n17704, A4 => 
                           n17703, ZN => n17720);
   U2012 : AOI22_X1 port map( A1 => n17708, A2 => REGISTERS_21_0_port, B1 => 
                           n17707, B2 => REGISTERS_24_0_port, ZN => n17718);
   U2013 : AOI22_X1 port map( A1 => n17710, A2 => REGISTERS_22_0_port, B1 => 
                           n17709, B2 => REGISTERS_16_0_port, ZN => n17717);
   U2014 : AOI22_X1 port map( A1 => n17712, A2 => REGISTERS_28_0_port, B1 => 
                           n17711, B2 => REGISTERS_18_0_port, ZN => n17716);
   U2015 : AOI22_X1 port map( A1 => n17714, A2 => REGISTERS_25_0_port, B1 => 
                           n17713, B2 => REGISTERS_19_0_port, ZN => n17715);
   U2016 : NAND4_X1 port map( A1 => n17718, A2 => n17717, A3 => n17716, A4 => 
                           n17715, ZN => n17719);
   U2017 : NOR2_X1 port map( A1 => n17720, A2 => n17719, ZN => n17748);
   U2018 : AOI22_X1 port map( A1 => n17721, A2 => REGISTERS_5_0_port, B1 => 
                           n17735, B2 => REGISTERS_7_0_port, ZN => n17730);
   U2019 : AOI22_X1 port map( A1 => n17723, A2 => REGISTERS_1_0_port, B1 => 
                           n17722, B2 => REGISTERS_0_0_port, ZN => n17729);
   U2020 : AOI22_X1 port map( A1 => n17725, A2 => REGISTERS_4_0_port, B1 => 
                           n17724, B2 => REGISTERS_2_0_port, ZN => n17728);
   U2021 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_6_0_port, B1 => 
                           n17726, B2 => REGISTERS_3_0_port, ZN => n17727);
   U2022 : NAND4_X1 port map( A1 => n17730, A2 => n17729, A3 => n17728, A4 => 
                           n17727, ZN => n17745);
   U2023 : AOI22_X1 port map( A1 => n17732, A2 => REGISTERS_13_0_port, B1 => 
                           n17731, B2 => REGISTERS_10_0_port, ZN => n17742);
   U2024 : AOI22_X1 port map( A1 => n17734, A2 => REGISTERS_14_0_port, B1 => 
                           n17733, B2 => REGISTERS_9_0_port, ZN => n17741);
   U2025 : AOI22_X1 port map( A1 => n17736, A2 => REGISTERS_12_0_port, B1 => 
                           n17735, B2 => REGISTERS_15_0_port, ZN => n17740);
   U2026 : AOI22_X1 port map( A1 => n17738, A2 => REGISTERS_11_0_port, B1 => 
                           n17737, B2 => REGISTERS_8_0_port, ZN => n17739);
   U2027 : NAND4_X1 port map( A1 => n17742, A2 => n17741, A3 => n17740, A4 => 
                           n17739, ZN => n17743);
   U2028 : AOI22_X1 port map( A1 => n17746, A2 => n17745, B1 => n17744, B2 => 
                           n17743, ZN => n17747);
   U2029 : OAI21_X1 port map( B1 => n17749, B2 => n17748, A => n17747, ZN => 
                           N417);
   U2030 : NAND3_X1 port map( A1 => n16783, A2 => ENABLE, A3 => RD1, ZN => 
                           n18531);
   U2031 : INV_X1 port map( A => ADD_RD1(3), ZN => n17772);
   U2032 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n17772, ZN => n17758);
   U2033 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), ZN => n17750);
   U2034 : INV_X1 port map( A => ADD_RD1(2), ZN => n17757);
   U2035 : NAND2_X1 port map( A1 => n17750, A2 => n17757, ZN => n17766);
   U2036 : NOR2_X1 port map( A1 => n17758, A2 => n17766, ZN => n18396);
   U2037 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n17759)
                           ;
   U2038 : INV_X1 port map( A => ADD_RD1(0), ZN => n17755);
   U2039 : OR3_X1 port map( A1 => n17757, A2 => n17755, A3 => ADD_RD1(1), ZN =>
                           n17909);
   U2040 : NOR2_X1 port map( A1 => n17759, A2 => n17909, ZN => n18420);
   U2041 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n18396, B1 => 
                           REGISTERS_29_31_port, B2 => n18420, ZN => n17754);
   U2042 : INV_X1 port map( A => ADD_RD1(1), ZN => n17756);
   U2043 : OR3_X1 port map( A1 => n17756, A2 => n17755, A3 => ADD_RD1(2), ZN =>
                           n17814);
   U2044 : NOR2_X1 port map( A1 => n17759, A2 => n17814, ZN => n18477);
   U2045 : CLKBUF_X1 port map( A => n18477, Z => n18368);
   U2046 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => n17750, ZN => n17767);
   U2047 : NOR2_X1 port map( A1 => n17758, A2 => n17767, ZN => n18443);
   U2048 : AOI22_X1 port map( A1 => REGISTERS_27_31_port, A2 => n18368, B1 => 
                           REGISTERS_20_31_port, B2 => n18443, ZN => n17753);
   U2049 : OR3_X1 port map( A1 => n17755, A2 => ADD_RD1(2), A3 => ADD_RD1(1), 
                           ZN => n17791);
   U2050 : NOR2_X1 port map( A1 => n17759, A2 => n17791, ZN => n18342);
   U2051 : CLKBUF_X1 port map( A => n18342, Z => n18496);
   U2052 : NOR2_X1 port map( A1 => n17758, A2 => n17814, ZN => n18205);
   U2053 : CLKBUF_X1 port map( A => n18205, Z => n18491);
   U2054 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n18496, B1 => 
                           REGISTERS_19_31_port, B2 => n18491, ZN => n17752);
   U2055 : OR3_X1 port map( A1 => n17756, A2 => n17757, A3 => ADD_RD1(0), ZN =>
                           n17837);
   U2056 : NOR2_X1 port map( A1 => n17837, A2 => n17758, ZN => n18441);
   U2057 : CLKBUF_X1 port map( A => n18441, Z => n18478);
   U2058 : NOR2_X1 port map( A1 => n17758, A2 => n17791, ZN => n18347);
   U2059 : CLKBUF_X1 port map( A => n18347, Z => n18480);
   U2060 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n18478, B1 => 
                           REGISTERS_17_31_port, B2 => n18480, ZN => n17751);
   U2061 : NAND4_X1 port map( A1 => n17754, A2 => n17753, A3 => n17752, A4 => 
                           n17751, ZN => n17765);
   U2062 : NOR2_X1 port map( A1 => n17759, A2 => n17767, ZN => n18272);
   U2063 : CLKBUF_X1 port map( A => n18272, Z => n18482);
   U2064 : OR3_X1 port map( A1 => n17756, A2 => ADD_RD1(2), A3 => ADD_RD1(0), 
                           ZN => n17932);
   U2065 : NOR2_X1 port map( A1 => n17758, A2 => n17932, ZN => n18295);
   U2066 : CLKBUF_X1 port map( A => n18295, Z => n18493);
   U2067 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n18482, B1 => 
                           REGISTERS_18_31_port, B2 => n18493, ZN => n17763);
   U2068 : NOR2_X1 port map( A1 => n17759, A2 => n17837, ZN => n18483);
   U2069 : CLKBUF_X1 port map( A => n18483, Z => n18449);
   U2070 : OR3_X1 port map( A1 => n17757, A2 => n17756, A3 => n17755, ZN => 
                           n17842);
   U2071 : NOR2_X1 port map( A1 => n17759, A2 => n17842, ZN => n18322);
   U2072 : CLKBUF_X1 port map( A => n18322, Z => n18479);
   U2073 : AOI22_X1 port map( A1 => REGISTERS_30_31_port, A2 => n18449, B1 => 
                           REGISTERS_31_31_port, B2 => n18479, ZN => n17762);
   U2074 : NOR2_X1 port map( A1 => n17758, A2 => n17909, ZN => n18484);
   U2075 : CLKBUF_X1 port map( A => n18484, Z => n18415);
   U2076 : NOR2_X1 port map( A1 => n17759, A2 => n17932, ZN => n18440);
   U2077 : CLKBUF_X1 port map( A => n18440, Z => n18490);
   U2078 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n18415, B1 => 
                           REGISTERS_26_31_port, B2 => n18490, ZN => n17761);
   U2079 : NOR2_X1 port map( A1 => n17842, A2 => n17758, ZN => n18489);
   U2080 : CLKBUF_X1 port map( A => n18489, Z => n18442);
   U2081 : NOR2_X1 port map( A1 => n17759, A2 => n17766, ZN => n18492);
   U2082 : CLKBUF_X1 port map( A => n18492, Z => n18448);
   U2083 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n18442, B1 => 
                           REGISTERS_24_31_port, B2 => n18448, ZN => n17760);
   U2084 : NAND4_X1 port map( A1 => n17763, A2 => n17762, A3 => n17761, A4 => 
                           n17760, ZN => n17764);
   U2085 : NOR2_X1 port map( A1 => n17765, A2 => n17764, ZN => n17780);
   U2086 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n18476, 
                           ZN => n18528);
   U2087 : CLKBUF_X1 port map( A => n18528, Z => n18339);
   U2088 : INV_X1 port map( A => n17814, ZN => n18507);
   U2089 : INV_X1 port map( A => n17766, ZN => n18464);
   U2090 : CLKBUF_X1 port map( A => n18464, Z => n18519);
   U2091 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n18507, B1 => 
                           REGISTERS_0_31_port, B2 => n18519, ZN => n17771);
   U2092 : INV_X1 port map( A => n17909, ZN => n18457);
   U2093 : INV_X1 port map( A => n17842, ZN => n18520);
   U2094 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n18457, B1 => 
                           REGISTERS_7_31_port, B2 => n18520, ZN => n17770);
   U2095 : INV_X1 port map( A => n17791, ZN => n18427);
   U2096 : INV_X1 port map( A => n17837, ZN => n18465);
   U2097 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n18427, B1 => 
                           REGISTERS_6_31_port, B2 => n18465, ZN => n17769);
   U2098 : INV_X1 port map( A => n17932, ZN => n18516);
   U2099 : INV_X1 port map( A => n17767, ZN => n18514);
   U2100 : CLKBUF_X1 port map( A => n18514, Z => n18466);
   U2101 : AOI22_X1 port map( A1 => REGISTERS_2_31_port, A2 => n18516, B1 => 
                           REGISTERS_4_31_port, B2 => n18466, ZN => n17768);
   U2102 : NAND4_X1 port map( A1 => n17771, A2 => n17770, A3 => n17769, A4 => 
                           n17768, ZN => n17778);
   U2103 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n17772, A3 => n18476, ZN 
                           => n18526);
   U2104 : CLKBUF_X1 port map( A => n18526, Z => n18363);
   U2105 : INV_X1 port map( A => n17791, ZN => n18459);
   U2106 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n18459, B1 => 
                           REGISTERS_15_31_port, B2 => n18520, ZN => n17776);
   U2107 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n18507, B1 => 
                           REGISTERS_10_31_port, B2 => n18516, ZN => n17775);
   U2108 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n18519, B1 => 
                           REGISTERS_13_31_port, B2 => n18457, ZN => n17774);
   U2109 : INV_X1 port map( A => n17837, ZN => n18517);
   U2110 : AOI22_X1 port map( A1 => REGISTERS_14_31_port, A2 => n18517, B1 => 
                           REGISTERS_12_31_port, B2 => n18466, ZN => n17773);
   U2111 : NAND4_X1 port map( A1 => n17776, A2 => n17775, A3 => n17774, A4 => 
                           n17773, ZN => n17777);
   U2112 : AOI22_X1 port map( A1 => n18339, A2 => n17778, B1 => n18363, B2 => 
                           n17777, ZN => n17779);
   U2113 : OAI21_X1 port map( B1 => n18476, B2 => n17780, A => n17779, ZN => 
                           N416);
   U2114 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n18480, B1 => 
                           REGISTERS_23_30_port, B2 => n18489, ZN => n17784);
   U2115 : CLKBUF_X1 port map( A => n18443, Z => n18495);
   U2116 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n18495, B1 => 
                           REGISTERS_21_30_port, B2 => n18484, ZN => n17783);
   U2117 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n18448, B1 => 
                           REGISTERS_29_30_port, B2 => n18420, ZN => n17782);
   U2118 : AOI22_X1 port map( A1 => REGISTERS_26_30_port, A2 => n18490, B1 => 
                           REGISTERS_31_30_port, B2 => n18322, ZN => n17781);
   U2119 : NAND4_X1 port map( A1 => n17784, A2 => n17783, A3 => n17782, A4 => 
                           n17781, ZN => n17790);
   U2120 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n18368, B1 => 
                           REGISTERS_30_30_port, B2 => n18449, ZN => n17788);
   U2121 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n18482, B1 => 
                           REGISTERS_25_30_port, B2 => n18496, ZN => n17787);
   U2122 : AOI22_X1 port map( A1 => REGISTERS_22_30_port, A2 => n18478, B1 => 
                           REGISTERS_18_30_port, B2 => n18295, ZN => n17786);
   U2123 : CLKBUF_X1 port map( A => n18396, Z => n18494);
   U2124 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n18494, B1 => 
                           REGISTERS_19_30_port, B2 => n18205, ZN => n17785);
   U2125 : NAND4_X1 port map( A1 => n17788, A2 => n17787, A3 => n17786, A4 => 
                           n17785, ZN => n17789);
   U2126 : NOR2_X1 port map( A1 => n17790, A2 => n17789, ZN => n17803);
   U2127 : INV_X1 port map( A => n17791, ZN => n18515);
   U2128 : AOI22_X1 port map( A1 => REGISTERS_2_30_port, A2 => n18516, B1 => 
                           REGISTERS_1_30_port, B2 => n18515, ZN => n17795);
   U2129 : INV_X1 port map( A => n17814, ZN => n18513);
   U2130 : AOI22_X1 port map( A1 => REGISTERS_7_30_port, A2 => n18520, B1 => 
                           REGISTERS_3_30_port, B2 => n18513, ZN => n17794);
   U2131 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n18519, B1 => 
                           REGISTERS_6_30_port, B2 => n18517, ZN => n17793);
   U2132 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n18514, B1 => 
                           REGISTERS_5_30_port, B2 => n18457, ZN => n17792);
   U2133 : NAND4_X1 port map( A1 => n17795, A2 => n17794, A3 => n17793, A4 => 
                           n17792, ZN => n17801);
   U2134 : INV_X1 port map( A => n17842, ZN => n18504);
   U2135 : CLKBUF_X1 port map( A => n18464, Z => n18503);
   U2136 : AOI22_X1 port map( A1 => REGISTERS_15_30_port, A2 => n18504, B1 => 
                           REGISTERS_8_30_port, B2 => n18503, ZN => n17799);
   U2137 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n18427, B1 => 
                           REGISTERS_10_30_port, B2 => n18516, ZN => n17798);
   U2138 : AOI22_X1 port map( A1 => REGISTERS_11_30_port, A2 => n18513, B1 => 
                           REGISTERS_14_30_port, B2 => n18517, ZN => n17797);
   U2139 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n18466, B1 => 
                           REGISTERS_13_30_port, B2 => n18457, ZN => n17796);
   U2140 : NAND4_X1 port map( A1 => n17799, A2 => n17798, A3 => n17797, A4 => 
                           n17796, ZN => n17800);
   U2141 : AOI22_X1 port map( A1 => n18339, A2 => n17801, B1 => n18363, B2 => 
                           n17800, ZN => n17802);
   U2142 : OAI21_X1 port map( B1 => n18476, B2 => n17803, A => n17802, ZN => 
                           N415);
   U2143 : AOI22_X1 port map( A1 => REGISTERS_21_29_port, A2 => n18415, B1 => 
                           REGISTERS_31_29_port, B2 => n18322, ZN => n17807);
   U2144 : AOI22_X1 port map( A1 => REGISTERS_30_29_port, A2 => n18449, B1 => 
                           REGISTERS_16_29_port, B2 => n18396, ZN => n17806);
   U2145 : CLKBUF_X1 port map( A => n18420, Z => n18481);
   U2146 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n18481, B1 => 
                           REGISTERS_24_29_port, B2 => n18492, ZN => n17805);
   U2147 : AOI22_X1 port map( A1 => REGISTERS_26_29_port, A2 => n18490, B1 => 
                           REGISTERS_18_29_port, B2 => n18295, ZN => n17804);
   U2148 : NAND4_X1 port map( A1 => n17807, A2 => n17806, A3 => n17805, A4 => 
                           n17804, ZN => n17813);
   U2149 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n18482, B1 => 
                           REGISTERS_19_29_port, B2 => n18205, ZN => n17811);
   U2150 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n18368, B1 => 
                           REGISTERS_17_29_port, B2 => n18480, ZN => n17810);
   U2151 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n18442, B1 => 
                           REGISTERS_25_29_port, B2 => n18342, ZN => n17809);
   U2152 : AOI22_X1 port map( A1 => REGISTERS_22_29_port, A2 => n18478, B1 => 
                           REGISTERS_20_29_port, B2 => n18443, ZN => n17808);
   U2153 : NAND4_X1 port map( A1 => n17811, A2 => n17810, A3 => n17809, A4 => 
                           n17808, ZN => n17812);
   U2154 : NOR2_X1 port map( A1 => n17813, A2 => n17812, ZN => n17826);
   U2155 : AOI22_X1 port map( A1 => REGISTERS_5_29_port, A2 => n18457, B1 => 
                           REGISTERS_7_29_port, B2 => n18520, ZN => n17818);
   U2156 : INV_X1 port map( A => n17814, ZN => n18383);
   U2157 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n18383, B1 => 
                           REGISTERS_2_29_port, B2 => n18516, ZN => n17817);
   U2158 : AOI22_X1 port map( A1 => REGISTERS_1_29_port, A2 => n18459, B1 => 
                           REGISTERS_0_29_port, B2 => n18503, ZN => n17816);
   U2159 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n18514, B1 => 
                           REGISTERS_6_29_port, B2 => n18517, ZN => n17815);
   U2160 : NAND4_X1 port map( A1 => n17818, A2 => n17817, A3 => n17816, A4 => 
                           n17815, ZN => n17824);
   U2161 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n18520, B1 => 
                           REGISTERS_14_29_port, B2 => n18517, ZN => n17822);
   U2162 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n18507, B1 => 
                           REGISTERS_8_29_port, B2 => n18503, ZN => n17821);
   U2163 : INV_X1 port map( A => n17932, ZN => n18508);
   U2164 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n18514, B1 => 
                           REGISTERS_10_29_port, B2 => n18508, ZN => n17820);
   U2165 : INV_X1 port map( A => n17909, ZN => n18505);
   U2166 : AOI22_X1 port map( A1 => REGISTERS_9_29_port, A2 => n18515, B1 => 
                           REGISTERS_13_29_port, B2 => n18505, ZN => n17819);
   U2167 : NAND4_X1 port map( A1 => n17822, A2 => n17821, A3 => n17820, A4 => 
                           n17819, ZN => n17823);
   U2168 : AOI22_X1 port map( A1 => n18339, A2 => n17824, B1 => n18363, B2 => 
                           n17823, ZN => n17825);
   U2169 : OAI21_X1 port map( B1 => n18476, B2 => n17826, A => n17825, ZN => 
                           N414);
   U2170 : AOI22_X1 port map( A1 => REGISTERS_31_28_port, A2 => n18479, B1 => 
                           REGISTERS_18_28_port, B2 => n18295, ZN => n17830);
   U2171 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n18448, B1 => 
                           REGISTERS_22_28_port, B2 => n18441, ZN => n17829);
   U2172 : AOI22_X1 port map( A1 => REGISTERS_21_28_port, A2 => n18415, B1 => 
                           REGISTERS_27_28_port, B2 => n18368, ZN => n17828);
   U2173 : AOI22_X1 port map( A1 => REGISTERS_26_28_port, A2 => n18490, B1 => 
                           REGISTERS_23_28_port, B2 => n18489, ZN => n17827);
   U2174 : NAND4_X1 port map( A1 => n17830, A2 => n17829, A3 => n17828, A4 => 
                           n17827, ZN => n17836);
   U2175 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n18494, B1 => 
                           REGISTERS_29_28_port, B2 => n18420, ZN => n17834);
   U2176 : AOI22_X1 port map( A1 => REGISTERS_30_28_port, A2 => n18449, B1 => 
                           REGISTERS_25_28_port, B2 => n18342, ZN => n17833);
   U2177 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n18480, B1 => 
                           REGISTERS_28_28_port, B2 => n18482, ZN => n17832);
   U2178 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n18443, B1 => 
                           REGISTERS_19_28_port, B2 => n18205, ZN => n17831);
   U2179 : NAND4_X1 port map( A1 => n17834, A2 => n17833, A3 => n17832, A4 => 
                           n17831, ZN => n17835);
   U2180 : NOR2_X1 port map( A1 => n17836, A2 => n17835, ZN => n17850);
   U2181 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n18507, B1 => 
                           REGISTERS_4_28_port, B2 => n18514, ZN => n17841);
   U2182 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n18427, B1 => 
                           REGISTERS_2_28_port, B2 => n18508, ZN => n17840);
   U2183 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n18519, B1 => 
                           REGISTERS_7_28_port, B2 => n18520, ZN => n17839);
   U2184 : INV_X1 port map( A => n17837, ZN => n18456);
   U2185 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n18457, B1 => 
                           REGISTERS_6_28_port, B2 => n18456, ZN => n17838);
   U2186 : NAND4_X1 port map( A1 => n17841, A2 => n17840, A3 => n17839, A4 => 
                           n17838, ZN => n17848);
   U2187 : INV_X1 port map( A => n17842, ZN => n18458);
   U2188 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n18458, B1 => 
                           REGISTERS_13_28_port, B2 => n18505, ZN => n17846);
   U2189 : AOI22_X1 port map( A1 => REGISTERS_10_28_port, A2 => n18516, B1 => 
                           REGISTERS_8_28_port, B2 => n18503, ZN => n17845);
   U2190 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n18459, B1 => 
                           REGISTERS_12_28_port, B2 => n18466, ZN => n17844);
   U2191 : AOI22_X1 port map( A1 => REGISTERS_14_28_port, A2 => n18465, B1 => 
                           REGISTERS_11_28_port, B2 => n18513, ZN => n17843);
   U2192 : NAND4_X1 port map( A1 => n17846, A2 => n17845, A3 => n17844, A4 => 
                           n17843, ZN => n17847);
   U2193 : AOI22_X1 port map( A1 => n18339, A2 => n17848, B1 => n18363, B2 => 
                           n17847, ZN => n17849);
   U2194 : OAI21_X1 port map( B1 => n18476, B2 => n17850, A => n17849, ZN => 
                           N413);
   U2195 : AOI22_X1 port map( A1 => REGISTERS_26_27_port, A2 => n18490, B1 => 
                           REGISTERS_28_27_port, B2 => n18272, ZN => n17854);
   U2196 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n18443, B1 => 
                           REGISTERS_30_27_port, B2 => n18483, ZN => n17853);
   U2197 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n18368, B1 => 
                           REGISTERS_19_27_port, B2 => n18205, ZN => n17852);
   U2198 : AOI22_X1 port map( A1 => REGISTERS_23_27_port, A2 => n18442, B1 => 
                           REGISTERS_22_27_port, B2 => n18441, ZN => n17851);
   U2199 : NAND4_X1 port map( A1 => n17854, A2 => n17853, A3 => n17852, A4 => 
                           n17851, ZN => n17860);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n18448, B1 => 
                           REGISTERS_25_27_port, B2 => n18342, ZN => n17858);
   U2201 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n18480, B1 => 
                           REGISTERS_21_27_port, B2 => n18484, ZN => n17857);
   U2202 : AOI22_X1 port map( A1 => REGISTERS_31_27_port, A2 => n18479, B1 => 
                           REGISTERS_16_27_port, B2 => n18396, ZN => n17856);
   U2203 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n18481, B1 => 
                           REGISTERS_18_27_port, B2 => n18295, ZN => n17855);
   U2204 : NAND4_X1 port map( A1 => n17858, A2 => n17857, A3 => n17856, A4 => 
                           n17855, ZN => n17859);
   U2205 : NOR2_X1 port map( A1 => n17860, A2 => n17859, ZN => n17872);
   U2206 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n18457, B1 => 
                           REGISTERS_1_27_port, B2 => n18427, ZN => n17864);
   U2207 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n18520, B1 => 
                           REGISTERS_6_27_port, B2 => n18456, ZN => n17863);
   U2208 : CLKBUF_X1 port map( A => n18514, Z => n18506);
   U2209 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n18506, B1 => 
                           REGISTERS_2_27_port, B2 => n18508, ZN => n17862);
   U2210 : AOI22_X1 port map( A1 => REGISTERS_3_27_port, A2 => n18507, B1 => 
                           REGISTERS_0_27_port, B2 => n18503, ZN => n17861);
   U2211 : NAND4_X1 port map( A1 => n17864, A2 => n17863, A3 => n17862, A4 => 
                           n17861, ZN => n17870);
   U2212 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n18507, B1 => 
                           REGISTERS_9_27_port, B2 => n18427, ZN => n17868);
   U2213 : AOI22_X1 port map( A1 => REGISTERS_13_27_port, A2 => n18457, B1 => 
                           REGISTERS_15_27_port, B2 => n18458, ZN => n17867);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_14_27_port, A2 => n18517, B1 => 
                           REGISTERS_8_27_port, B2 => n18464, ZN => n17866);
   U2215 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n18466, B1 => 
                           REGISTERS_10_27_port, B2 => n18508, ZN => n17865);
   U2216 : NAND4_X1 port map( A1 => n17868, A2 => n17867, A3 => n17866, A4 => 
                           n17865, ZN => n17869);
   U2217 : AOI22_X1 port map( A1 => n18339, A2 => n17870, B1 => n18363, B2 => 
                           n17869, ZN => n17871);
   U2218 : OAI21_X1 port map( B1 => n18476, B2 => n17872, A => n17871, ZN => 
                           N412);
   U2219 : AOI22_X1 port map( A1 => REGISTERS_22_26_port, A2 => n18478, B1 => 
                           REGISTERS_19_26_port, B2 => n18205, ZN => n17876);
   U2220 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n18481, B1 => 
                           REGISTERS_21_26_port, B2 => n18415, ZN => n17875);
   U2221 : AOI22_X1 port map( A1 => REGISTERS_23_26_port, A2 => n18442, B1 => 
                           REGISTERS_20_26_port, B2 => n18495, ZN => n17874);
   U2222 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n18494, B1 => 
                           REGISTERS_30_26_port, B2 => n18483, ZN => n17873);
   U2223 : NAND4_X1 port map( A1 => n17876, A2 => n17875, A3 => n17874, A4 => 
                           n17873, ZN => n17882);
   U2224 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n18448, B1 => 
                           REGISTERS_17_26_port, B2 => n18347, ZN => n17880);
   U2225 : AOI22_X1 port map( A1 => REGISTERS_26_26_port, A2 => n18490, B1 => 
                           REGISTERS_31_26_port, B2 => n18322, ZN => n17879);
   U2226 : AOI22_X1 port map( A1 => REGISTERS_25_26_port, A2 => n18496, B1 => 
                           REGISTERS_28_26_port, B2 => n18272, ZN => n17878);
   U2227 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n18477, B1 => 
                           REGISTERS_18_26_port, B2 => n18295, ZN => n17877);
   U2228 : NAND4_X1 port map( A1 => n17880, A2 => n17879, A3 => n17878, A4 => 
                           n17877, ZN => n17881);
   U2229 : NOR2_X1 port map( A1 => n17882, A2 => n17881, ZN => n17894);
   U2230 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n18457, B1 => 
                           REGISTERS_2_26_port, B2 => n18508, ZN => n17886);
   U2231 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n18506, B1 => 
                           REGISTERS_3_26_port, B2 => n18507, ZN => n17885);
   U2232 : AOI22_X1 port map( A1 => REGISTERS_6_26_port, A2 => n18465, B1 => 
                           REGISTERS_0_26_port, B2 => n18503, ZN => n17884);
   U2233 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n18520, B1 => 
                           REGISTERS_1_26_port, B2 => n18427, ZN => n17883);
   U2234 : NAND4_X1 port map( A1 => n17886, A2 => n17885, A3 => n17884, A4 => 
                           n17883, ZN => n17892);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n18457, B1 => 
                           REGISTERS_12_26_port, B2 => n18466, ZN => n17890);
   U2236 : AOI22_X1 port map( A1 => REGISTERS_10_26_port, A2 => n18516, B1 => 
                           REGISTERS_14_26_port, B2 => n18456, ZN => n17889);
   U2237 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n18458, B1 => 
                           REGISTERS_11_26_port, B2 => n18513, ZN => n17888);
   U2238 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n18519, B1 => 
                           REGISTERS_9_26_port, B2 => n18427, ZN => n17887);
   U2239 : NAND4_X1 port map( A1 => n17890, A2 => n17889, A3 => n17888, A4 => 
                           n17887, ZN => n17891);
   U2240 : AOI22_X1 port map( A1 => n18339, A2 => n17892, B1 => n18363, B2 => 
                           n17891, ZN => n17893);
   U2241 : OAI21_X1 port map( B1 => n18476, B2 => n17894, A => n17893, ZN => 
                           N411);
   U2242 : AOI22_X1 port map( A1 => REGISTERS_18_25_port, A2 => n18493, B1 => 
                           REGISTERS_19_25_port, B2 => n18205, ZN => n17898);
   U2243 : AOI22_X1 port map( A1 => REGISTERS_23_25_port, A2 => n18442, B1 => 
                           REGISTERS_27_25_port, B2 => n18368, ZN => n17897);
   U2244 : AOI22_X1 port map( A1 => REGISTERS_26_25_port, A2 => n18490, B1 => 
                           REGISTERS_24_25_port, B2 => n18492, ZN => n17896);
   U2245 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n18481, B1 => 
                           REGISTERS_22_25_port, B2 => n18441, ZN => n17895);
   U2246 : NAND4_X1 port map( A1 => n17898, A2 => n17897, A3 => n17896, A4 => 
                           n17895, ZN => n17904);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n18494, B1 => 
                           REGISTERS_28_25_port, B2 => n18272, ZN => n17902);
   U2248 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n18443, B1 => 
                           REGISTERS_21_25_port, B2 => n18415, ZN => n17901);
   U2249 : AOI22_X1 port map( A1 => REGISTERS_31_25_port, A2 => n18479, B1 => 
                           REGISTERS_25_25_port, B2 => n18342, ZN => n17900);
   U2250 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n18480, B1 => 
                           REGISTERS_30_25_port, B2 => n18483, ZN => n17899);
   U2251 : NAND4_X1 port map( A1 => n17902, A2 => n17901, A3 => n17900, A4 => 
                           n17899, ZN => n17903);
   U2252 : NOR2_X1 port map( A1 => n17904, A2 => n17903, ZN => n17917);
   U2253 : AOI22_X1 port map( A1 => REGISTERS_7_25_port, A2 => n18520, B1 => 
                           REGISTERS_3_25_port, B2 => n18383, ZN => n17908);
   U2254 : AOI22_X1 port map( A1 => REGISTERS_6_25_port, A2 => n18517, B1 => 
                           REGISTERS_4_25_port, B2 => n18466, ZN => n17907);
   U2255 : AOI22_X1 port map( A1 => REGISTERS_2_25_port, A2 => n18508, B1 => 
                           REGISTERS_5_25_port, B2 => n18505, ZN => n17906);
   U2256 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n18519, B1 => 
                           REGISTERS_1_25_port, B2 => n18459, ZN => n17905);
   U2257 : NAND4_X1 port map( A1 => n17908, A2 => n17907, A3 => n17906, A4 => 
                           n17905, ZN => n17915);
   U2258 : INV_X1 port map( A => n17909, ZN => n18518);
   U2259 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n18514, B1 => 
                           REGISTERS_13_25_port, B2 => n18518, ZN => n17913);
   U2260 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n18507, B1 => 
                           REGISTERS_14_25_port, B2 => n18456, ZN => n17912);
   U2261 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n18520, B1 => 
                           REGISTERS_8_25_port, B2 => n18464, ZN => n17911);
   U2262 : AOI22_X1 port map( A1 => REGISTERS_10_25_port, A2 => n18516, B1 => 
                           REGISTERS_9_25_port, B2 => n18459, ZN => n17910);
   U2263 : NAND4_X1 port map( A1 => n17913, A2 => n17912, A3 => n17911, A4 => 
                           n17910, ZN => n17914);
   U2264 : AOI22_X1 port map( A1 => n18339, A2 => n17915, B1 => n18363, B2 => 
                           n17914, ZN => n17916);
   U2265 : OAI21_X1 port map( B1 => n18476, B2 => n17917, A => n17916, ZN => 
                           N410);
   U2266 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n18494, B1 => 
                           REGISTERS_31_24_port, B2 => n18322, ZN => n17921);
   U2267 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n18481, B1 => 
                           REGISTERS_24_24_port, B2 => n18492, ZN => n17920);
   U2268 : AOI22_X1 port map( A1 => REGISTERS_30_24_port, A2 => n18449, B1 => 
                           REGISTERS_28_24_port, B2 => n18272, ZN => n17919);
   U2269 : AOI22_X1 port map( A1 => REGISTERS_26_24_port, A2 => n18490, B1 => 
                           REGISTERS_21_24_port, B2 => n18415, ZN => n17918);
   U2270 : NAND4_X1 port map( A1 => n17921, A2 => n17920, A3 => n17919, A4 => 
                           n17918, ZN => n17927);
   U2271 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n18442, B1 => 
                           REGISTERS_19_24_port, B2 => n18205, ZN => n17925);
   U2272 : AOI22_X1 port map( A1 => REGISTERS_25_24_port, A2 => n18496, B1 => 
                           REGISTERS_17_24_port, B2 => n18347, ZN => n17924);
   U2273 : AOI22_X1 port map( A1 => REGISTERS_22_24_port, A2 => n18478, B1 => 
                           REGISTERS_27_24_port, B2 => n18368, ZN => n17923);
   U2274 : AOI22_X1 port map( A1 => REGISTERS_18_24_port, A2 => n18493, B1 => 
                           REGISTERS_20_24_port, B2 => n18495, ZN => n17922);
   U2275 : NAND4_X1 port map( A1 => n17925, A2 => n17924, A3 => n17923, A4 => 
                           n17922, ZN => n17926);
   U2276 : NOR2_X1 port map( A1 => n17927, A2 => n17926, ZN => n17940);
   U2277 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n18515, B1 => 
                           REGISTERS_0_24_port, B2 => n18503, ZN => n17931);
   U2278 : AOI22_X1 port map( A1 => REGISTERS_2_24_port, A2 => n18516, B1 => 
                           REGISTERS_5_24_port, B2 => n18518, ZN => n17930);
   U2279 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n18507, B1 => 
                           REGISTERS_6_24_port, B2 => n18456, ZN => n17929);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n18506, B1 => 
                           REGISTERS_7_24_port, B2 => n18458, ZN => n17928);
   U2281 : NAND4_X1 port map( A1 => n17931, A2 => n17930, A3 => n17929, A4 => 
                           n17928, ZN => n17938);
   U2282 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n18515, B1 => 
                           REGISTERS_15_24_port, B2 => n18458, ZN => n17936);
   U2283 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n18507, B1 => 
                           REGISTERS_13_24_port, B2 => n18518, ZN => n17935);
   U2284 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n18514, B1 => 
                           REGISTERS_8_24_port, B2 => n18464, ZN => n17934);
   U2285 : INV_X1 port map( A => n17932, ZN => n18467);
   U2286 : AOI22_X1 port map( A1 => REGISTERS_14_24_port, A2 => n18465, B1 => 
                           REGISTERS_10_24_port, B2 => n18467, ZN => n17933);
   U2287 : NAND4_X1 port map( A1 => n17936, A2 => n17935, A3 => n17934, A4 => 
                           n17933, ZN => n17937);
   U2288 : AOI22_X1 port map( A1 => n18339, A2 => n17938, B1 => n18363, B2 => 
                           n17937, ZN => n17939);
   U2289 : OAI21_X1 port map( B1 => n18476, B2 => n17940, A => n17939, ZN => 
                           N409);
   U2290 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n18481, B1 => 
                           REGISTERS_17_23_port, B2 => n18347, ZN => n17944);
   U2291 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n18415, B1 => 
                           REGISTERS_28_23_port, B2 => n18482, ZN => n17943);
   U2292 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n18495, B1 => 
                           REGISTERS_18_23_port, B2 => n18295, ZN => n17942);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n18494, B1 => 
                           REGISTERS_19_23_port, B2 => n18205, ZN => n17941);
   U2294 : NAND4_X1 port map( A1 => n17944, A2 => n17943, A3 => n17942, A4 => 
                           n17941, ZN => n17950);
   U2295 : AOI22_X1 port map( A1 => REGISTERS_23_23_port, A2 => n18442, B1 => 
                           REGISTERS_24_23_port, B2 => n18492, ZN => n17948);
   U2296 : AOI22_X1 port map( A1 => REGISTERS_31_23_port, A2 => n18479, B1 => 
                           REGISTERS_25_23_port, B2 => n18496, ZN => n17947);
   U2297 : AOI22_X1 port map( A1 => REGISTERS_27_23_port, A2 => n18477, B1 => 
                           REGISTERS_30_23_port, B2 => n18449, ZN => n17946);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_22_23_port, A2 => n18478, B1 => 
                           REGISTERS_26_23_port, B2 => n18490, ZN => n17945);
   U2299 : NAND4_X1 port map( A1 => n17948, A2 => n17947, A3 => n17946, A4 => 
                           n17945, ZN => n17949);
   U2300 : NOR2_X1 port map( A1 => n17950, A2 => n17949, ZN => n17962);
   U2301 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n18457, B1 => 
                           REGISTERS_3_23_port, B2 => n18383, ZN => n17954);
   U2302 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n18459, B1 => 
                           REGISTERS_0_23_port, B2 => n18503, ZN => n17953);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n18458, B1 => 
                           REGISTERS_4_23_port, B2 => n18514, ZN => n17952);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_2_23_port, A2 => n18516, B1 => 
                           REGISTERS_6_23_port, B2 => n18456, ZN => n17951);
   U2305 : NAND4_X1 port map( A1 => n17954, A2 => n17953, A3 => n17952, A4 => 
                           n17951, ZN => n17960);
   U2306 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n18520, B1 => 
                           REGISTERS_14_23_port, B2 => n18456, ZN => n17958);
   U2307 : AOI22_X1 port map( A1 => REGISTERS_10_23_port, A2 => n18516, B1 => 
                           REGISTERS_11_23_port, B2 => n18513, ZN => n17957);
   U2308 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n18506, B1 => 
                           REGISTERS_8_23_port, B2 => n18464, ZN => n17956);
   U2309 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n18457, B1 => 
                           REGISTERS_9_23_port, B2 => n18459, ZN => n17955);
   U2310 : NAND4_X1 port map( A1 => n17958, A2 => n17957, A3 => n17956, A4 => 
                           n17955, ZN => n17959);
   U2311 : AOI22_X1 port map( A1 => n18339, A2 => n17960, B1 => n18363, B2 => 
                           n17959, ZN => n17961);
   U2312 : OAI21_X1 port map( B1 => n18531, B2 => n17962, A => n17961, ZN => 
                           N408);
   U2313 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n18415, B1 => 
                           REGISTERS_20_22_port, B2 => n18495, ZN => n17966);
   U2314 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n18448, B1 => 
                           REGISTERS_29_22_port, B2 => n18481, ZN => n17965);
   U2315 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n18480, B1 => 
                           REGISTERS_19_22_port, B2 => n18491, ZN => n17964);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n18442, B1 => 
                           REGISTERS_28_22_port, B2 => n18272, ZN => n17963);
   U2317 : NAND4_X1 port map( A1 => n17966, A2 => n17965, A3 => n17964, A4 => 
                           n17963, ZN => n17972);
   U2318 : AOI22_X1 port map( A1 => REGISTERS_27_22_port, A2 => n18368, B1 => 
                           REGISTERS_16_22_port, B2 => n18494, ZN => n17970);
   U2319 : AOI22_X1 port map( A1 => REGISTERS_31_22_port, A2 => n18479, B1 => 
                           REGISTERS_25_22_port, B2 => n18342, ZN => n17969);
   U2320 : AOI22_X1 port map( A1 => REGISTERS_22_22_port, A2 => n18478, B1 => 
                           REGISTERS_30_22_port, B2 => n18483, ZN => n17968);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_18_22_port, A2 => n18493, B1 => 
                           REGISTERS_26_22_port, B2 => n18440, ZN => n17967);
   U2322 : NAND4_X1 port map( A1 => n17970, A2 => n17969, A3 => n17968, A4 => 
                           n17967, ZN => n17971);
   U2323 : NOR2_X1 port map( A1 => n17972, A2 => n17971, ZN => n17984);
   U2324 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n18520, B1 => 
                           REGISTERS_3_22_port, B2 => n18507, ZN => n17976);
   U2325 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n18519, B1 => 
                           REGISTERS_2_22_port, B2 => n18467, ZN => n17975);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_6_22_port, A2 => n18465, B1 => 
                           REGISTERS_1_22_port, B2 => n18459, ZN => n17974);
   U2327 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n18466, B1 => 
                           REGISTERS_5_22_port, B2 => n18518, ZN => n17973);
   U2328 : NAND4_X1 port map( A1 => n17976, A2 => n17975, A3 => n17974, A4 => 
                           n17973, ZN => n17982);
   U2329 : AOI22_X1 port map( A1 => REGISTERS_14_22_port, A2 => n18465, B1 => 
                           REGISTERS_8_22_port, B2 => n18503, ZN => n17980);
   U2330 : AOI22_X1 port map( A1 => REGISTERS_9_22_port, A2 => n18515, B1 => 
                           REGISTERS_11_22_port, B2 => n18383, ZN => n17979);
   U2331 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n18518, B1 => 
                           REGISTERS_15_22_port, B2 => n18458, ZN => n17978);
   U2332 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n18514, B1 => 
                           REGISTERS_10_22_port, B2 => n18467, ZN => n17977);
   U2333 : NAND4_X1 port map( A1 => n17980, A2 => n17979, A3 => n17978, A4 => 
                           n17977, ZN => n17981);
   U2334 : AOI22_X1 port map( A1 => n18339, A2 => n17982, B1 => n18363, B2 => 
                           n17981, ZN => n17983);
   U2335 : OAI21_X1 port map( B1 => n18531, B2 => n17984, A => n17983, ZN => 
                           N407);
   U2336 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n18415, B1 => 
                           REGISTERS_31_21_port, B2 => n18322, ZN => n17988);
   U2337 : AOI22_X1 port map( A1 => REGISTERS_17_21_port, A2 => n18347, B1 => 
                           REGISTERS_23_21_port, B2 => n18489, ZN => n17987);
   U2338 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n18495, B1 => 
                           REGISTERS_28_21_port, B2 => n18272, ZN => n17986);
   U2339 : AOI22_X1 port map( A1 => REGISTERS_18_21_port, A2 => n18295, B1 => 
                           REGISTERS_19_21_port, B2 => n18491, ZN => n17985);
   U2340 : NAND4_X1 port map( A1 => n17988, A2 => n17987, A3 => n17986, A4 => 
                           n17985, ZN => n17994);
   U2341 : AOI22_X1 port map( A1 => REGISTERS_25_21_port, A2 => n18496, B1 => 
                           REGISTERS_27_21_port, B2 => n18368, ZN => n17992);
   U2342 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n18481, B1 => 
                           REGISTERS_26_21_port, B2 => n18440, ZN => n17991);
   U2343 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n18478, B1 => 
                           REGISTERS_16_21_port, B2 => n18494, ZN => n17990);
   U2344 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n18448, B1 => 
                           REGISTERS_30_21_port, B2 => n18483, ZN => n17989);
   U2345 : NAND4_X1 port map( A1 => n17992, A2 => n17991, A3 => n17990, A4 => 
                           n17989, ZN => n17993);
   U2346 : NOR2_X1 port map( A1 => n17994, A2 => n17993, ZN => n18006);
   U2347 : AOI22_X1 port map( A1 => REGISTERS_6_21_port, A2 => n18465, B1 => 
                           REGISTERS_1_21_port, B2 => n18459, ZN => n17998);
   U2348 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n18505, B1 => 
                           REGISTERS_3_21_port, B2 => n18513, ZN => n17997);
   U2349 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n18458, B1 => 
                           REGISTERS_4_21_port, B2 => n18514, ZN => n17996);
   U2350 : AOI22_X1 port map( A1 => REGISTERS_2_21_port, A2 => n18467, B1 => 
                           REGISTERS_0_21_port, B2 => n18464, ZN => n17995);
   U2351 : NAND4_X1 port map( A1 => n17998, A2 => n17997, A3 => n17996, A4 => 
                           n17995, ZN => n18004);
   U2352 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n18466, B1 => 
                           REGISTERS_10_21_port, B2 => n18467, ZN => n18002);
   U2353 : AOI22_X1 port map( A1 => REGISTERS_11_21_port, A2 => n18383, B1 => 
                           REGISTERS_15_21_port, B2 => n18458, ZN => n18001);
   U2354 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n18457, B1 => 
                           REGISTERS_14_21_port, B2 => n18456, ZN => n18000);
   U2355 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n18519, B1 => 
                           REGISTERS_9_21_port, B2 => n18459, ZN => n17999);
   U2356 : NAND4_X1 port map( A1 => n18002, A2 => n18001, A3 => n18000, A4 => 
                           n17999, ZN => n18003);
   U2357 : AOI22_X1 port map( A1 => n18339, A2 => n18004, B1 => n18363, B2 => 
                           n18003, ZN => n18005);
   U2358 : OAI21_X1 port map( B1 => n18531, B2 => n18006, A => n18005, ZN => 
                           N406);
   U2359 : AOI22_X1 port map( A1 => REGISTERS_22_20_port, A2 => n18441, B1 => 
                           REGISTERS_26_20_port, B2 => n18440, ZN => n18010);
   U2360 : AOI22_X1 port map( A1 => REGISTERS_23_20_port, A2 => n18442, B1 => 
                           REGISTERS_31_20_port, B2 => n18322, ZN => n18009);
   U2361 : AOI22_X1 port map( A1 => REGISTERS_19_20_port, A2 => n18205, B1 => 
                           REGISTERS_18_20_port, B2 => n18295, ZN => n18008);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n18368, B1 => 
                           REGISTERS_28_20_port, B2 => n18272, ZN => n18007);
   U2363 : NAND4_X1 port map( A1 => n18010, A2 => n18009, A3 => n18008, A4 => 
                           n18007, ZN => n18016);
   U2364 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n18448, B1 => 
                           REGISTERS_25_20_port, B2 => n18342, ZN => n18014);
   U2365 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n18495, B1 => 
                           REGISTERS_29_20_port, B2 => n18481, ZN => n18013);
   U2366 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n18396, B1 => 
                           REGISTERS_17_20_port, B2 => n18347, ZN => n18012);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_21_20_port, A2 => n18415, B1 => 
                           REGISTERS_30_20_port, B2 => n18483, ZN => n18011);
   U2368 : NAND4_X1 port map( A1 => n18014, A2 => n18013, A3 => n18012, A4 => 
                           n18011, ZN => n18015);
   U2369 : NOR2_X1 port map( A1 => n18016, A2 => n18015, ZN => n18028);
   U2370 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n18519, B1 => 
                           REGISTERS_3_20_port, B2 => n18383, ZN => n18020);
   U2371 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n18518, B1 => 
                           REGISTERS_7_20_port, B2 => n18504, ZN => n18019);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n18459, B1 => 
                           REGISTERS_2_20_port, B2 => n18467, ZN => n18018);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_6_20_port, A2 => n18465, B1 => 
                           REGISTERS_4_20_port, B2 => n18466, ZN => n18017);
   U2374 : NAND4_X1 port map( A1 => n18020, A2 => n18019, A3 => n18018, A4 => 
                           n18017, ZN => n18026);
   U2375 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n18519, B1 => 
                           REGISTERS_11_20_port, B2 => n18383, ZN => n18024);
   U2376 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n18427, B1 => 
                           REGISTERS_12_20_port, B2 => n18466, ZN => n18023);
   U2377 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n18457, B1 => 
                           REGISTERS_15_20_port, B2 => n18520, ZN => n18022);
   U2378 : AOI22_X1 port map( A1 => REGISTERS_10_20_port, A2 => n18467, B1 => 
                           REGISTERS_14_20_port, B2 => n18456, ZN => n18021);
   U2379 : NAND4_X1 port map( A1 => n18024, A2 => n18023, A3 => n18022, A4 => 
                           n18021, ZN => n18025);
   U2380 : AOI22_X1 port map( A1 => n18339, A2 => n18026, B1 => n18526, B2 => 
                           n18025, ZN => n18027);
   U2381 : OAI21_X1 port map( B1 => n18531, B2 => n18028, A => n18027, ZN => 
                           N405);
   U2382 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n18484, B1 => 
                           REGISTERS_17_19_port, B2 => n18347, ZN => n18032);
   U2383 : AOI22_X1 port map( A1 => REGISTERS_31_19_port, A2 => n18322, B1 => 
                           REGISTERS_29_19_port, B2 => n18481, ZN => n18031);
   U2384 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n18448, B1 => 
                           REGISTERS_28_19_port, B2 => n18272, ZN => n18030);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n18342, B1 => 
                           REGISTERS_19_19_port, B2 => n18491, ZN => n18029);
   U2386 : NAND4_X1 port map( A1 => n18032, A2 => n18031, A3 => n18030, A4 => 
                           n18029, ZN => n18038);
   U2387 : AOI22_X1 port map( A1 => REGISTERS_18_19_port, A2 => n18493, B1 => 
                           REGISTERS_27_19_port, B2 => n18368, ZN => n18036);
   U2388 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n18442, B1 => 
                           REGISTERS_20_19_port, B2 => n18495, ZN => n18035);
   U2389 : AOI22_X1 port map( A1 => REGISTERS_30_19_port, A2 => n18483, B1 => 
                           REGISTERS_26_19_port, B2 => n18440, ZN => n18034);
   U2390 : AOI22_X1 port map( A1 => REGISTERS_22_19_port, A2 => n18441, B1 => 
                           REGISTERS_16_19_port, B2 => n18494, ZN => n18033);
   U2391 : NAND4_X1 port map( A1 => n18036, A2 => n18035, A3 => n18034, A4 => 
                           n18033, ZN => n18037);
   U2392 : NOR2_X1 port map( A1 => n18038, A2 => n18037, ZN => n18050);
   U2393 : CLKBUF_X1 port map( A => n18528, Z => n18365);
   U2394 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n18519, B1 => 
                           REGISTERS_1_19_port, B2 => n18459, ZN => n18042);
   U2395 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n18506, B1 => 
                           REGISTERS_7_19_port, B2 => n18458, ZN => n18041);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_2_19_port, A2 => n18467, B1 => 
                           REGISTERS_6_19_port, B2 => n18456, ZN => n18040);
   U2397 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n18518, B1 => 
                           REGISTERS_3_19_port, B2 => n18383, ZN => n18039);
   U2398 : NAND4_X1 port map( A1 => n18042, A2 => n18041, A3 => n18040, A4 => 
                           n18039, ZN => n18048);
   U2399 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n18513, B1 => 
                           REGISTERS_8_19_port, B2 => n18503, ZN => n18046);
   U2400 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n18518, B1 => 
                           REGISTERS_10_19_port, B2 => n18516, ZN => n18045);
   U2401 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n18504, B1 => 
                           REGISTERS_9_19_port, B2 => n18459, ZN => n18044);
   U2402 : AOI22_X1 port map( A1 => REGISTERS_14_19_port, A2 => n18465, B1 => 
                           REGISTERS_12_19_port, B2 => n18506, ZN => n18043);
   U2403 : NAND4_X1 port map( A1 => n18046, A2 => n18045, A3 => n18044, A4 => 
                           n18043, ZN => n18047);
   U2404 : AOI22_X1 port map( A1 => n18365, A2 => n18048, B1 => n18363, B2 => 
                           n18047, ZN => n18049);
   U2405 : OAI21_X1 port map( B1 => n18531, B2 => n18050, A => n18049, ZN => 
                           N404);
   U2406 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n18489, B1 => 
                           REGISTERS_16_18_port, B2 => n18396, ZN => n18054);
   U2407 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n18347, B1 => 
                           REGISTERS_22_18_port, B2 => n18441, ZN => n18053);
   U2408 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n18368, B1 => 
                           REGISTERS_28_18_port, B2 => n18482, ZN => n18052);
   U2409 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n18420, B1 => 
                           REGISTERS_25_18_port, B2 => n18342, ZN => n18051);
   U2410 : NAND4_X1 port map( A1 => n18054, A2 => n18053, A3 => n18052, A4 => 
                           n18051, ZN => n18060);
   U2411 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n18492, B1 => 
                           REGISTERS_26_18_port, B2 => n18440, ZN => n18058);
   U2412 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n18484, B1 => 
                           REGISTERS_19_18_port, B2 => n18491, ZN => n18057);
   U2413 : AOI22_X1 port map( A1 => REGISTERS_30_18_port, A2 => n18483, B1 => 
                           REGISTERS_18_18_port, B2 => n18295, ZN => n18056);
   U2414 : AOI22_X1 port map( A1 => REGISTERS_31_18_port, A2 => n18479, B1 => 
                           REGISTERS_20_18_port, B2 => n18495, ZN => n18055);
   U2415 : NAND4_X1 port map( A1 => n18058, A2 => n18057, A3 => n18056, A4 => 
                           n18055, ZN => n18059);
   U2416 : NOR2_X1 port map( A1 => n18060, A2 => n18059, ZN => n18072);
   U2417 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n18464, B1 => 
                           REGISTERS_2_18_port, B2 => n18508, ZN => n18064);
   U2418 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n18515, B1 => 
                           REGISTERS_3_18_port, B2 => n18507, ZN => n18063);
   U2419 : AOI22_X1 port map( A1 => REGISTERS_6_18_port, A2 => n18465, B1 => 
                           REGISTERS_4_18_port, B2 => n18506, ZN => n18062);
   U2420 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n18504, B1 => 
                           REGISTERS_5_18_port, B2 => n18518, ZN => n18061);
   U2421 : NAND4_X1 port map( A1 => n18064, A2 => n18063, A3 => n18062, A4 => 
                           n18061, ZN => n18070);
   U2422 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n18514, B1 => 
                           REGISTERS_8_18_port, B2 => n18464, ZN => n18068);
   U2423 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n18505, B1 => 
                           REGISTERS_11_18_port, B2 => n18383, ZN => n18067);
   U2424 : AOI22_X1 port map( A1 => REGISTERS_10_18_port, A2 => n18508, B1 => 
                           REGISTERS_14_18_port, B2 => n18456, ZN => n18066);
   U2425 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n18427, B1 => 
                           REGISTERS_15_18_port, B2 => n18520, ZN => n18065);
   U2426 : NAND4_X1 port map( A1 => n18068, A2 => n18067, A3 => n18066, A4 => 
                           n18065, ZN => n18069);
   U2427 : AOI22_X1 port map( A1 => n18365, A2 => n18070, B1 => n18363, B2 => 
                           n18069, ZN => n18071);
   U2428 : OAI21_X1 port map( B1 => n18531, B2 => n18072, A => n18071, ZN => 
                           N403);
   U2429 : AOI22_X1 port map( A1 => REGISTERS_26_17_port, A2 => n18490, B1 => 
                           REGISTERS_20_17_port, B2 => n18495, ZN => n18076);
   U2430 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n18396, B1 => 
                           REGISTERS_25_17_port, B2 => n18342, ZN => n18075);
   U2431 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n18415, B1 => 
                           REGISTERS_22_17_port, B2 => n18478, ZN => n18074);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_30_17_port, A2 => n18483, B1 => 
                           REGISTERS_23_17_port, B2 => n18442, ZN => n18073);
   U2433 : NAND4_X1 port map( A1 => n18076, A2 => n18075, A3 => n18074, A4 => 
                           n18073, ZN => n18082);
   U2434 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n18420, B1 => 
                           REGISTERS_19_17_port, B2 => n18491, ZN => n18080);
   U2435 : AOI22_X1 port map( A1 => REGISTERS_27_17_port, A2 => n18368, B1 => 
                           REGISTERS_17_17_port, B2 => n18347, ZN => n18079);
   U2436 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n18272, B1 => 
                           REGISTERS_24_17_port, B2 => n18492, ZN => n18078);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_18_17_port, A2 => n18295, B1 => 
                           REGISTERS_31_17_port, B2 => n18322, ZN => n18077);
   U2438 : NAND4_X1 port map( A1 => n18080, A2 => n18079, A3 => n18078, A4 => 
                           n18077, ZN => n18081);
   U2439 : NOR2_X1 port map( A1 => n18082, A2 => n18081, ZN => n18094);
   U2440 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n18466, B1 => 
                           REGISTERS_2_17_port, B2 => n18516, ZN => n18086);
   U2441 : AOI22_X1 port map( A1 => REGISTERS_6_17_port, A2 => n18465, B1 => 
                           REGISTERS_3_17_port, B2 => n18383, ZN => n18085);
   U2442 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n18464, B1 => 
                           REGISTERS_1_17_port, B2 => n18459, ZN => n18084);
   U2443 : AOI22_X1 port map( A1 => REGISTERS_5_17_port, A2 => n18457, B1 => 
                           REGISTERS_7_17_port, B2 => n18458, ZN => n18083);
   U2444 : NAND4_X1 port map( A1 => n18086, A2 => n18085, A3 => n18084, A4 => 
                           n18083, ZN => n18092);
   U2445 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n18504, B1 => 
                           REGISTERS_8_17_port, B2 => n18464, ZN => n18090);
   U2446 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n18506, B1 => 
                           REGISTERS_14_17_port, B2 => n18456, ZN => n18089);
   U2447 : AOI22_X1 port map( A1 => REGISTERS_9_17_port, A2 => n18515, B1 => 
                           REGISTERS_10_17_port, B2 => n18467, ZN => n18088);
   U2448 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n18507, B1 => 
                           REGISTERS_13_17_port, B2 => n18518, ZN => n18087);
   U2449 : NAND4_X1 port map( A1 => n18090, A2 => n18089, A3 => n18088, A4 => 
                           n18087, ZN => n18091);
   U2450 : AOI22_X1 port map( A1 => n18365, A2 => n18092, B1 => n18363, B2 => 
                           n18091, ZN => n18093);
   U2451 : OAI21_X1 port map( B1 => n18531, B2 => n18094, A => n18093, ZN => 
                           N402);
   U2452 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n18420, B1 => 
                           REGISTERS_22_16_port, B2 => n18478, ZN => n18098);
   U2453 : AOI22_X1 port map( A1 => REGISTERS_18_16_port, A2 => n18493, B1 => 
                           REGISTERS_19_16_port, B2 => n18491, ZN => n18097);
   U2454 : AOI22_X1 port map( A1 => REGISTERS_27_16_port, A2 => n18368, B1 => 
                           REGISTERS_17_16_port, B2 => n18347, ZN => n18096);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n18495, B1 => 
                           REGISTERS_28_16_port, B2 => n18482, ZN => n18095);
   U2456 : NAND4_X1 port map( A1 => n18098, A2 => n18097, A3 => n18096, A4 => 
                           n18095, ZN => n18104);
   U2457 : AOI22_X1 port map( A1 => REGISTERS_23_16_port, A2 => n18489, B1 => 
                           REGISTERS_26_16_port, B2 => n18440, ZN => n18102);
   U2458 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n18492, B1 => 
                           REGISTERS_25_16_port, B2 => n18496, ZN => n18101);
   U2459 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n18494, B1 => 
                           REGISTERS_31_16_port, B2 => n18322, ZN => n18100);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_21_16_port, A2 => n18415, B1 => 
                           REGISTERS_30_16_port, B2 => n18483, ZN => n18099);
   U2461 : NAND4_X1 port map( A1 => n18102, A2 => n18101, A3 => n18100, A4 => 
                           n18099, ZN => n18103);
   U2462 : NOR2_X1 port map( A1 => n18104, A2 => n18103, ZN => n18116);
   U2463 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n18505, B1 => 
                           REGISTERS_2_16_port, B2 => n18467, ZN => n18108);
   U2464 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n18519, B1 => 
                           REGISTERS_7_16_port, B2 => n18520, ZN => n18107);
   U2465 : AOI22_X1 port map( A1 => REGISTERS_6_16_port, A2 => n18456, B1 => 
                           REGISTERS_4_16_port, B2 => n18514, ZN => n18106);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n18427, B1 => 
                           REGISTERS_3_16_port, B2 => n18383, ZN => n18105);
   U2467 : NAND4_X1 port map( A1 => n18108, A2 => n18107, A3 => n18106, A4 => 
                           n18105, ZN => n18114);
   U2468 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n18513, B1 => 
                           REGISTERS_14_16_port, B2 => n18517, ZN => n18112);
   U2469 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n18516, B1 => 
                           REGISTERS_13_16_port, B2 => n18518, ZN => n18111);
   U2470 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n18504, B1 => 
                           REGISTERS_8_16_port, B2 => n18503, ZN => n18110);
   U2471 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n18506, B1 => 
                           REGISTERS_9_16_port, B2 => n18459, ZN => n18109);
   U2472 : NAND4_X1 port map( A1 => n18112, A2 => n18111, A3 => n18110, A4 => 
                           n18109, ZN => n18113);
   U2473 : AOI22_X1 port map( A1 => n18365, A2 => n18114, B1 => n18363, B2 => 
                           n18113, ZN => n18115);
   U2474 : OAI21_X1 port map( B1 => n18531, B2 => n18116, A => n18115, ZN => 
                           N401);
   U2475 : AOI22_X1 port map( A1 => REGISTERS_18_15_port, A2 => n18493, B1 => 
                           REGISTERS_26_15_port, B2 => n18440, ZN => n18120);
   U2476 : AOI22_X1 port map( A1 => REGISTERS_23_15_port, A2 => n18489, B1 => 
                           REGISTERS_20_15_port, B2 => n18495, ZN => n18119);
   U2477 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n18415, B1 => 
                           REGISTERS_17_15_port, B2 => n18347, ZN => n18118);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n18448, B1 => 
                           REGISTERS_16_15_port, B2 => n18494, ZN => n18117);
   U2479 : NAND4_X1 port map( A1 => n18120, A2 => n18119, A3 => n18118, A4 => 
                           n18117, ZN => n18126);
   U2480 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n18205, B1 => 
                           REGISTERS_29_15_port, B2 => n18420, ZN => n18124);
   U2481 : AOI22_X1 port map( A1 => REGISTERS_30_15_port, A2 => n18449, B1 => 
                           REGISTERS_25_15_port, B2 => n18496, ZN => n18123);
   U2482 : AOI22_X1 port map( A1 => REGISTERS_22_15_port, A2 => n18478, B1 => 
                           REGISTERS_28_15_port, B2 => n18482, ZN => n18122);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n18479, B1 => 
                           REGISTERS_27_15_port, B2 => n18368, ZN => n18121);
   U2484 : NAND4_X1 port map( A1 => n18124, A2 => n18123, A3 => n18122, A4 => 
                           n18121, ZN => n18125);
   U2485 : NOR2_X1 port map( A1 => n18126, A2 => n18125, ZN => n18138);
   U2486 : AOI22_X1 port map( A1 => REGISTERS_6_15_port, A2 => n18456, B1 => 
                           REGISTERS_3_15_port, B2 => n18383, ZN => n18130);
   U2487 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n18506, B1 => 
                           REGISTERS_7_15_port, B2 => n18458, ZN => n18129);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_2_15_port, A2 => n18508, B1 => 
                           REGISTERS_0_15_port, B2 => n18464, ZN => n18128);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n18518, B1 => 
                           REGISTERS_1_15_port, B2 => n18459, ZN => n18127);
   U2490 : NAND4_X1 port map( A1 => n18130, A2 => n18129, A3 => n18128, A4 => 
                           n18127, ZN => n18136);
   U2491 : AOI22_X1 port map( A1 => REGISTERS_11_15_port, A2 => n18383, B1 => 
                           REGISTERS_10_15_port, B2 => n18467, ZN => n18134);
   U2492 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n18515, B1 => 
                           REGISTERS_14_15_port, B2 => n18517, ZN => n18133);
   U2493 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n18504, B1 => 
                           REGISTERS_12_15_port, B2 => n18514, ZN => n18132);
   U2494 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n18505, B1 => 
                           REGISTERS_8_15_port, B2 => n18503, ZN => n18131);
   U2495 : NAND4_X1 port map( A1 => n18134, A2 => n18133, A3 => n18132, A4 => 
                           n18131, ZN => n18135);
   U2496 : AOI22_X1 port map( A1 => n18365, A2 => n18136, B1 => n18363, B2 => 
                           n18135, ZN => n18137);
   U2497 : OAI21_X1 port map( B1 => n18476, B2 => n18138, A => n18137, ZN => 
                           N400);
   U2498 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n18481, B1 => 
                           REGISTERS_17_14_port, B2 => n18480, ZN => n18142);
   U2499 : AOI22_X1 port map( A1 => REGISTERS_22_14_port, A2 => n18478, B1 => 
                           REGISTERS_25_14_port, B2 => n18496, ZN => n18141);
   U2500 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n18448, B1 => 
                           REGISTERS_19_14_port, B2 => n18491, ZN => n18140);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_27_14_port, A2 => n18368, B1 => 
                           REGISTERS_20_14_port, B2 => n18495, ZN => n18139);
   U2502 : NAND4_X1 port map( A1 => n18142, A2 => n18141, A3 => n18140, A4 => 
                           n18139, ZN => n18148);
   U2503 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n18482, B1 => 
                           REGISTERS_23_14_port, B2 => n18442, ZN => n18146);
   U2504 : AOI22_X1 port map( A1 => REGISTERS_30_14_port, A2 => n18449, B1 => 
                           REGISTERS_16_14_port, B2 => n18494, ZN => n18145);
   U2505 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n18415, B1 => 
                           REGISTERS_26_14_port, B2 => n18440, ZN => n18144);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_18_14_port, A2 => n18493, B1 => 
                           REGISTERS_31_14_port, B2 => n18479, ZN => n18143);
   U2507 : NAND4_X1 port map( A1 => n18146, A2 => n18145, A3 => n18144, A4 => 
                           n18143, ZN => n18147);
   U2508 : NOR2_X1 port map( A1 => n18148, A2 => n18147, ZN => n18160);
   U2509 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n18504, B1 => 
                           REGISTERS_1_14_port, B2 => n18459, ZN => n18152);
   U2510 : AOI22_X1 port map( A1 => REGISTERS_6_14_port, A2 => n18465, B1 => 
                           REGISTERS_4_14_port, B2 => n18466, ZN => n18151);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_2_14_port, A2 => n18467, B1 => 
                           REGISTERS_0_14_port, B2 => n18464, ZN => n18150);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_3_14_port, A2 => n18513, B1 => 
                           REGISTERS_5_14_port, B2 => n18518, ZN => n18149);
   U2513 : NAND4_X1 port map( A1 => n18152, A2 => n18151, A3 => n18150, A4 => 
                           n18149, ZN => n18158);
   U2514 : AOI22_X1 port map( A1 => REGISTERS_9_14_port, A2 => n18515, B1 => 
                           REGISTERS_13_14_port, B2 => n18518, ZN => n18156);
   U2515 : AOI22_X1 port map( A1 => REGISTERS_15_14_port, A2 => n18504, B1 => 
                           REGISTERS_14_14_port, B2 => n18517, ZN => n18155);
   U2516 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n18507, B1 => 
                           REGISTERS_10_14_port, B2 => n18467, ZN => n18154);
   U2517 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n18506, B1 => 
                           REGISTERS_8_14_port, B2 => n18503, ZN => n18153);
   U2518 : NAND4_X1 port map( A1 => n18156, A2 => n18155, A3 => n18154, A4 => 
                           n18153, ZN => n18157);
   U2519 : AOI22_X1 port map( A1 => n18365, A2 => n18158, B1 => n18363, B2 => 
                           n18157, ZN => n18159);
   U2520 : OAI21_X1 port map( B1 => n18531, B2 => n18160, A => n18159, ZN => 
                           N399);
   U2521 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n18494, B1 => 
                           REGISTERS_18_13_port, B2 => n18493, ZN => n18164);
   U2522 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n18482, B1 => 
                           REGISTERS_31_13_port, B2 => n18479, ZN => n18163);
   U2523 : AOI22_X1 port map( A1 => REGISTERS_26_13_port, A2 => n18490, B1 => 
                           REGISTERS_24_13_port, B2 => n18492, ZN => n18162);
   U2524 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n18481, B1 => 
                           REGISTERS_17_13_port, B2 => n18480, ZN => n18161);
   U2525 : NAND4_X1 port map( A1 => n18164, A2 => n18163, A3 => n18162, A4 => 
                           n18161, ZN => n18170);
   U2526 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n18496, B1 => 
                           REGISTERS_27_13_port, B2 => n18368, ZN => n18168);
   U2527 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n18442, B1 => 
                           REGISTERS_20_13_port, B2 => n18495, ZN => n18167);
   U2528 : AOI22_X1 port map( A1 => REGISTERS_22_13_port, A2 => n18478, B1 => 
                           REGISTERS_19_13_port, B2 => n18491, ZN => n18166);
   U2529 : AOI22_X1 port map( A1 => REGISTERS_30_13_port, A2 => n18449, B1 => 
                           REGISTERS_21_13_port, B2 => n18415, ZN => n18165);
   U2530 : NAND4_X1 port map( A1 => n18168, A2 => n18167, A3 => n18166, A4 => 
                           n18165, ZN => n18169);
   U2531 : NOR2_X1 port map( A1 => n18170, A2 => n18169, ZN => n18182);
   U2532 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n18464, B1 => 
                           REGISTERS_5_13_port, B2 => n18518, ZN => n18174);
   U2533 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n18427, B1 => 
                           REGISTERS_6_13_port, B2 => n18517, ZN => n18173);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_2_13_port, A2 => n18508, B1 => 
                           REGISTERS_3_13_port, B2 => n18383, ZN => n18172);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n18504, B1 => 
                           REGISTERS_4_13_port, B2 => n18506, ZN => n18171);
   U2536 : NAND4_X1 port map( A1 => n18174, A2 => n18173, A3 => n18172, A4 => 
                           n18171, ZN => n18180);
   U2537 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n18504, B1 => 
                           REGISTERS_11_13_port, B2 => n18383, ZN => n18178);
   U2538 : AOI22_X1 port map( A1 => REGISTERS_10_13_port, A2 => n18516, B1 => 
                           REGISTERS_12_13_port, B2 => n18466, ZN => n18177);
   U2539 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n18427, B1 => 
                           REGISTERS_8_13_port, B2 => n18464, ZN => n18176);
   U2540 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n18457, B1 => 
                           REGISTERS_14_13_port, B2 => n18517, ZN => n18175);
   U2541 : NAND4_X1 port map( A1 => n18178, A2 => n18177, A3 => n18176, A4 => 
                           n18175, ZN => n18179);
   U2542 : AOI22_X1 port map( A1 => n18365, A2 => n18180, B1 => n18363, B2 => 
                           n18179, ZN => n18181);
   U2543 : OAI21_X1 port map( B1 => n18476, B2 => n18182, A => n18181, ZN => 
                           N398);
   U2544 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n18415, B1 => 
                           REGISTERS_26_12_port, B2 => n18490, ZN => n18186);
   U2545 : AOI22_X1 port map( A1 => REGISTERS_31_12_port, A2 => n18322, B1 => 
                           REGISTERS_30_12_port, B2 => n18449, ZN => n18185);
   U2546 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n18448, B1 => 
                           REGISTERS_22_12_port, B2 => n18478, ZN => n18184);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n18496, B1 => 
                           REGISTERS_17_12_port, B2 => n18480, ZN => n18183);
   U2548 : NAND4_X1 port map( A1 => n18186, A2 => n18185, A3 => n18184, A4 => 
                           n18183, ZN => n18192);
   U2549 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n18495, B1 => 
                           REGISTERS_19_12_port, B2 => n18491, ZN => n18190);
   U2550 : AOI22_X1 port map( A1 => REGISTERS_27_12_port, A2 => n18368, B1 => 
                           REGISTERS_23_12_port, B2 => n18489, ZN => n18189);
   U2551 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n18482, B1 => 
                           REGISTERS_18_12_port, B2 => n18493, ZN => n18188);
   U2552 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n18481, B1 => 
                           REGISTERS_16_12_port, B2 => n18494, ZN => n18187);
   U2553 : NAND4_X1 port map( A1 => n18190, A2 => n18189, A3 => n18188, A4 => 
                           n18187, ZN => n18191);
   U2554 : NOR2_X1 port map( A1 => n18192, A2 => n18191, ZN => n18204);
   U2555 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n18504, B1 => 
                           REGISTERS_6_12_port, B2 => n18517, ZN => n18196);
   U2556 : AOI22_X1 port map( A1 => REGISTERS_3_12_port, A2 => n18507, B1 => 
                           REGISTERS_5_12_port, B2 => n18518, ZN => n18195);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n18506, B1 => 
                           REGISTERS_1_12_port, B2 => n18515, ZN => n18194);
   U2558 : AOI22_X1 port map( A1 => REGISTERS_2_12_port, A2 => n18516, B1 => 
                           REGISTERS_0_12_port, B2 => n18503, ZN => n18193);
   U2559 : NAND4_X1 port map( A1 => n18196, A2 => n18195, A3 => n18194, A4 => 
                           n18193, ZN => n18202);
   U2560 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n18504, B1 => 
                           REGISTERS_13_12_port, B2 => n18505, ZN => n18200);
   U2561 : AOI22_X1 port map( A1 => REGISTERS_14_12_port, A2 => n18517, B1 => 
                           REGISTERS_11_12_port, B2 => n18513, ZN => n18199);
   U2562 : AOI22_X1 port map( A1 => REGISTERS_10_12_port, A2 => n18467, B1 => 
                           REGISTERS_8_12_port, B2 => n18464, ZN => n18198);
   U2563 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n18506, B1 => 
                           REGISTERS_9_12_port, B2 => n18515, ZN => n18197);
   U2564 : NAND4_X1 port map( A1 => n18200, A2 => n18199, A3 => n18198, A4 => 
                           n18197, ZN => n18201);
   U2565 : AOI22_X1 port map( A1 => n18365, A2 => n18202, B1 => n18363, B2 => 
                           n18201, ZN => n18203);
   U2566 : OAI21_X1 port map( B1 => n18531, B2 => n18204, A => n18203, ZN => 
                           N397);
   U2567 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n18448, B1 => 
                           REGISTERS_30_11_port, B2 => n18449, ZN => n18209);
   U2568 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n18496, B1 => 
                           REGISTERS_20_11_port, B2 => n18495, ZN => n18208);
   U2569 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n18205, B1 => 
                           REGISTERS_27_11_port, B2 => n18368, ZN => n18207);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_18_11_port, A2 => n18493, B1 => 
                           REGISTERS_16_11_port, B2 => n18396, ZN => n18206);
   U2571 : NAND4_X1 port map( A1 => n18209, A2 => n18208, A3 => n18207, A4 => 
                           n18206, ZN => n18215);
   U2572 : AOI22_X1 port map( A1 => REGISTERS_26_11_port, A2 => n18440, B1 => 
                           REGISTERS_31_11_port, B2 => n18479, ZN => n18213);
   U2573 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n18481, B1 => 
                           REGISTERS_22_11_port, B2 => n18478, ZN => n18212);
   U2574 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n18482, B1 => 
                           REGISTERS_21_11_port, B2 => n18415, ZN => n18211);
   U2575 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n18442, B1 => 
                           REGISTERS_17_11_port, B2 => n18480, ZN => n18210);
   U2576 : NAND4_X1 port map( A1 => n18213, A2 => n18212, A3 => n18211, A4 => 
                           n18210, ZN => n18214);
   U2577 : NOR2_X1 port map( A1 => n18215, A2 => n18214, ZN => n18227);
   U2578 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n18519, B1 => 
                           REGISTERS_1_11_port, B2 => n18515, ZN => n18219);
   U2579 : AOI22_X1 port map( A1 => REGISTERS_2_11_port, A2 => n18508, B1 => 
                           REGISTERS_4_11_port, B2 => n18514, ZN => n18218);
   U2580 : AOI22_X1 port map( A1 => REGISTERS_6_11_port, A2 => n18465, B1 => 
                           REGISTERS_7_11_port, B2 => n18520, ZN => n18217);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n18457, B1 => 
                           REGISTERS_3_11_port, B2 => n18383, ZN => n18216);
   U2582 : NAND4_X1 port map( A1 => n18219, A2 => n18218, A3 => n18217, A4 => 
                           n18216, ZN => n18225);
   U2583 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n18506, B1 => 
                           REGISTERS_9_11_port, B2 => n18515, ZN => n18223);
   U2584 : AOI22_X1 port map( A1 => REGISTERS_11_11_port, A2 => n18383, B1 => 
                           REGISTERS_13_11_port, B2 => n18518, ZN => n18222);
   U2585 : AOI22_X1 port map( A1 => REGISTERS_14_11_port, A2 => n18517, B1 => 
                           REGISTERS_10_11_port, B2 => n18467, ZN => n18221);
   U2586 : AOI22_X1 port map( A1 => REGISTERS_15_11_port, A2 => n18504, B1 => 
                           REGISTERS_8_11_port, B2 => n18503, ZN => n18220);
   U2587 : NAND4_X1 port map( A1 => n18223, A2 => n18222, A3 => n18221, A4 => 
                           n18220, ZN => n18224);
   U2588 : AOI22_X1 port map( A1 => n18365, A2 => n18225, B1 => n18363, B2 => 
                           n18224, ZN => n18226);
   U2589 : OAI21_X1 port map( B1 => n18531, B2 => n18227, A => n18226, ZN => 
                           N396);
   U2590 : AOI22_X1 port map( A1 => REGISTERS_25_10_port, A2 => n18496, B1 => 
                           REGISTERS_21_10_port, B2 => n18415, ZN => n18231);
   U2591 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n18272, B1 => 
                           REGISTERS_29_10_port, B2 => n18481, ZN => n18230);
   U2592 : AOI22_X1 port map( A1 => REGISTERS_31_10_port, A2 => n18479, B1 => 
                           REGISTERS_23_10_port, B2 => n18489, ZN => n18229);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_18_10_port, A2 => n18493, B1 => 
                           REGISTERS_30_10_port, B2 => n18449, ZN => n18228);
   U2594 : NAND4_X1 port map( A1 => n18231, A2 => n18230, A3 => n18229, A4 => 
                           n18228, ZN => n18237);
   U2595 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n18480, B1 => 
                           REGISTERS_22_10_port, B2 => n18478, ZN => n18235);
   U2596 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n18494, B1 => 
                           REGISTERS_26_10_port, B2 => n18490, ZN => n18234);
   U2597 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n18491, B1 => 
                           REGISTERS_27_10_port, B2 => n18477, ZN => n18233);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n18495, B1 => 
                           REGISTERS_24_10_port, B2 => n18492, ZN => n18232);
   U2599 : NAND4_X1 port map( A1 => n18235, A2 => n18234, A3 => n18233, A4 => 
                           n18232, ZN => n18236);
   U2600 : NOR2_X1 port map( A1 => n18237, A2 => n18236, ZN => n18249);
   U2601 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n18518, B1 => 
                           REGISTERS_6_10_port, B2 => n18517, ZN => n18241);
   U2602 : AOI22_X1 port map( A1 => REGISTERS_3_10_port, A2 => n18513, B1 => 
                           REGISTERS_1_10_port, B2 => n18515, ZN => n18240);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n18506, B1 => 
                           REGISTERS_0_10_port, B2 => n18464, ZN => n18239);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n18504, B1 => 
                           REGISTERS_2_10_port, B2 => n18467, ZN => n18238);
   U2605 : NAND4_X1 port map( A1 => n18241, A2 => n18240, A3 => n18239, A4 => 
                           n18238, ZN => n18247);
   U2606 : AOI22_X1 port map( A1 => REGISTERS_14_10_port, A2 => n18456, B1 => 
                           REGISTERS_10_10_port, B2 => n18467, ZN => n18245);
   U2607 : AOI22_X1 port map( A1 => REGISTERS_15_10_port, A2 => n18504, B1 => 
                           REGISTERS_12_10_port, B2 => n18514, ZN => n18244);
   U2608 : AOI22_X1 port map( A1 => REGISTERS_13_10_port, A2 => n18505, B1 => 
                           REGISTERS_11_10_port, B2 => n18383, ZN => n18243);
   U2609 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n18503, B1 => 
                           REGISTERS_9_10_port, B2 => n18515, ZN => n18242);
   U2610 : NAND4_X1 port map( A1 => n18245, A2 => n18244, A3 => n18243, A4 => 
                           n18242, ZN => n18246);
   U2611 : AOI22_X1 port map( A1 => n18365, A2 => n18247, B1 => n18363, B2 => 
                           n18246, ZN => n18248);
   U2612 : OAI21_X1 port map( B1 => n18531, B2 => n18249, A => n18248, ZN => 
                           N395);
   U2613 : AOI22_X1 port map( A1 => REGISTERS_26_9_port, A2 => n18490, B1 => 
                           REGISTERS_29_9_port, B2 => n18420, ZN => n18253);
   U2614 : AOI22_X1 port map( A1 => REGISTERS_30_9_port, A2 => n18449, B1 => 
                           REGISTERS_22_9_port, B2 => n18441, ZN => n18252);
   U2615 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n18442, B1 => 
                           REGISTERS_24_9_port, B2 => n18492, ZN => n18251);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n18495, B1 => 
                           REGISTERS_25_9_port, B2 => n18496, ZN => n18250);
   U2617 : NAND4_X1 port map( A1 => n18253, A2 => n18252, A3 => n18251, A4 => 
                           n18250, ZN => n18259);
   U2618 : AOI22_X1 port map( A1 => REGISTERS_19_9_port, A2 => n18491, B1 => 
                           REGISTERS_18_9_port, B2 => n18493, ZN => n18257);
   U2619 : AOI22_X1 port map( A1 => REGISTERS_31_9_port, A2 => n18479, B1 => 
                           REGISTERS_27_9_port, B2 => n18368, ZN => n18256);
   U2620 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n18480, B1 => 
                           REGISTERS_28_9_port, B2 => n18482, ZN => n18255);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n18494, B1 => 
                           REGISTERS_21_9_port, B2 => n18484, ZN => n18254);
   U2622 : NAND4_X1 port map( A1 => n18257, A2 => n18256, A3 => n18255, A4 => 
                           n18254, ZN => n18258);
   U2623 : NOR2_X1 port map( A1 => n18259, A2 => n18258, ZN => n18271);
   U2624 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n18504, B1 => 
                           REGISTERS_6_9_port, B2 => n18456, ZN => n18263);
   U2625 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n18507, B1 => 
                           REGISTERS_4_9_port, B2 => n18466, ZN => n18262);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n18464, B1 => 
                           REGISTERS_5_9_port, B2 => n18518, ZN => n18261);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n18427, B1 => 
                           REGISTERS_2_9_port, B2 => n18467, ZN => n18260);
   U2628 : NAND4_X1 port map( A1 => n18263, A2 => n18262, A3 => n18261, A4 => 
                           n18260, ZN => n18269);
   U2629 : AOI22_X1 port map( A1 => REGISTERS_14_9_port, A2 => n18465, B1 => 
                           REGISTERS_12_9_port, B2 => n18514, ZN => n18267);
   U2630 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n18457, B1 => 
                           REGISTERS_8_9_port, B2 => n18519, ZN => n18266);
   U2631 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n18427, B1 => 
                           REGISTERS_15_9_port, B2 => n18458, ZN => n18265);
   U2632 : AOI22_X1 port map( A1 => REGISTERS_11_9_port, A2 => n18383, B1 => 
                           REGISTERS_10_9_port, B2 => n18467, ZN => n18264);
   U2633 : NAND4_X1 port map( A1 => n18267, A2 => n18266, A3 => n18265, A4 => 
                           n18264, ZN => n18268);
   U2634 : AOI22_X1 port map( A1 => n18365, A2 => n18269, B1 => n18363, B2 => 
                           n18268, ZN => n18270);
   U2635 : OAI21_X1 port map( B1 => n18476, B2 => n18271, A => n18270, ZN => 
                           N394);
   U2636 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n18415, B1 => 
                           REGISTERS_31_8_port, B2 => n18479, ZN => n18276);
   U2637 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n18342, B1 => 
                           REGISTERS_29_8_port, B2 => n18420, ZN => n18275);
   U2638 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n18272, B1 => 
                           REGISTERS_24_8_port, B2 => n18448, ZN => n18274);
   U2639 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n18442, B1 => 
                           REGISTERS_26_8_port, B2 => n18490, ZN => n18273);
   U2640 : NAND4_X1 port map( A1 => n18276, A2 => n18275, A3 => n18274, A4 => 
                           n18273, ZN => n18282);
   U2641 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n18491, B1 => 
                           REGISTERS_22_8_port, B2 => n18441, ZN => n18280);
   U2642 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n18480, B1 => 
                           REGISTERS_18_8_port, B2 => n18493, ZN => n18279);
   U2643 : AOI22_X1 port map( A1 => REGISTERS_30_8_port, A2 => n18449, B1 => 
                           REGISTERS_20_8_port, B2 => n18443, ZN => n18278);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n18477, B1 => 
                           REGISTERS_16_8_port, B2 => n18396, ZN => n18277);
   U2645 : NAND4_X1 port map( A1 => n18280, A2 => n18279, A3 => n18278, A4 => 
                           n18277, ZN => n18281);
   U2646 : NOR2_X1 port map( A1 => n18282, A2 => n18281, ZN => n18294);
   U2647 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n18506, B1 => 
                           REGISTERS_6_8_port, B2 => n18517, ZN => n18286);
   U2648 : AOI22_X1 port map( A1 => REGISTERS_1_8_port, A2 => n18427, B1 => 
                           REGISTERS_2_8_port, B2 => n18508, ZN => n18285);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n18458, B1 => 
                           REGISTERS_5_8_port, B2 => n18505, ZN => n18284);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_3_8_port, A2 => n18513, B1 => 
                           REGISTERS_0_8_port, B2 => n18519, ZN => n18283);
   U2651 : NAND4_X1 port map( A1 => n18286, A2 => n18285, A3 => n18284, A4 => 
                           n18283, ZN => n18292);
   U2652 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n18520, B1 => 
                           REGISTERS_8_8_port, B2 => n18464, ZN => n18290);
   U2653 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n18506, B1 => 
                           REGISTERS_13_8_port, B2 => n18505, ZN => n18289);
   U2654 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n18383, B1 => 
                           REGISTERS_9_8_port, B2 => n18515, ZN => n18288);
   U2655 : AOI22_X1 port map( A1 => REGISTERS_14_8_port, A2 => n18465, B1 => 
                           REGISTERS_10_8_port, B2 => n18508, ZN => n18287);
   U2656 : NAND4_X1 port map( A1 => n18290, A2 => n18289, A3 => n18288, A4 => 
                           n18287, ZN => n18291);
   U2657 : AOI22_X1 port map( A1 => n18365, A2 => n18292, B1 => n18363, B2 => 
                           n18291, ZN => n18293);
   U2658 : OAI21_X1 port map( B1 => n18531, B2 => n18294, A => n18293, ZN => 
                           N393);
   U2659 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n18478, B1 => 
                           REGISTERS_27_7_port, B2 => n18477, ZN => n18299);
   U2660 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n18481, B1 => 
                           REGISTERS_26_7_port, B2 => n18490, ZN => n18298);
   U2661 : AOI22_X1 port map( A1 => REGISTERS_18_7_port, A2 => n18295, B1 => 
                           REGISTERS_23_7_port, B2 => n18489, ZN => n18297);
   U2662 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n18480, B1 => 
                           REGISTERS_21_7_port, B2 => n18484, ZN => n18296);
   U2663 : NAND4_X1 port map( A1 => n18299, A2 => n18298, A3 => n18297, A4 => 
                           n18296, ZN => n18305);
   U2664 : AOI22_X1 port map( A1 => REGISTERS_30_7_port, A2 => n18449, B1 => 
                           REGISTERS_25_7_port, B2 => n18496, ZN => n18303);
   U2665 : AOI22_X1 port map( A1 => REGISTERS_19_7_port, A2 => n18491, B1 => 
                           REGISTERS_20_7_port, B2 => n18443, ZN => n18302);
   U2666 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n18494, B1 => 
                           REGISTERS_31_7_port, B2 => n18479, ZN => n18301);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n18482, B1 => 
                           REGISTERS_24_7_port, B2 => n18448, ZN => n18300);
   U2668 : NAND4_X1 port map( A1 => n18303, A2 => n18302, A3 => n18301, A4 => 
                           n18300, ZN => n18304);
   U2669 : NOR2_X1 port map( A1 => n18305, A2 => n18304, ZN => n18317);
   U2670 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n18506, B1 => 
                           REGISTERS_6_7_port, B2 => n18465, ZN => n18309);
   U2671 : AOI22_X1 port map( A1 => REGISTERS_2_7_port, A2 => n18516, B1 => 
                           REGISTERS_1_7_port, B2 => n18515, ZN => n18308);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n18503, B1 => 
                           REGISTERS_7_7_port, B2 => n18458, ZN => n18307);
   U2673 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n18507, B1 => 
                           REGISTERS_5_7_port, B2 => n18505, ZN => n18306);
   U2674 : NAND4_X1 port map( A1 => n18309, A2 => n18308, A3 => n18307, A4 => 
                           n18306, ZN => n18315);
   U2675 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n18519, B1 => 
                           REGISTERS_13_7_port, B2 => n18505, ZN => n18313);
   U2676 : AOI22_X1 port map( A1 => REGISTERS_15_7_port, A2 => n18504, B1 => 
                           REGISTERS_9_7_port, B2 => n18427, ZN => n18312);
   U2677 : AOI22_X1 port map( A1 => REGISTERS_10_7_port, A2 => n18467, B1 => 
                           REGISTERS_12_7_port, B2 => n18514, ZN => n18311);
   U2678 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n18383, B1 => 
                           REGISTERS_14_7_port, B2 => n18517, ZN => n18310);
   U2679 : NAND4_X1 port map( A1 => n18313, A2 => n18312, A3 => n18311, A4 => 
                           n18310, ZN => n18314);
   U2680 : AOI22_X1 port map( A1 => n18365, A2 => n18315, B1 => n18363, B2 => 
                           n18314, ZN => n18316);
   U2681 : OAI21_X1 port map( B1 => n18476, B2 => n18317, A => n18316, ZN => 
                           N392);
   U2682 : AOI22_X1 port map( A1 => REGISTERS_19_6_port, A2 => n18491, B1 => 
                           REGISTERS_25_6_port, B2 => n18496, ZN => n18321);
   U2683 : AOI22_X1 port map( A1 => REGISTERS_22_6_port, A2 => n18478, B1 => 
                           REGISTERS_26_6_port, B2 => n18490, ZN => n18320);
   U2684 : AOI22_X1 port map( A1 => REGISTERS_30_6_port, A2 => n18449, B1 => 
                           REGISTERS_18_6_port, B2 => n18493, ZN => n18319);
   U2685 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n18448, B1 => 
                           REGISTERS_27_6_port, B2 => n18477, ZN => n18318);
   U2686 : NAND4_X1 port map( A1 => n18321, A2 => n18320, A3 => n18319, A4 => 
                           n18318, ZN => n18328);
   U2687 : AOI22_X1 port map( A1 => REGISTERS_23_6_port, A2 => n18442, B1 => 
                           REGISTERS_28_6_port, B2 => n18482, ZN => n18326);
   U2688 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n18481, B1 => 
                           REGISTERS_16_6_port, B2 => n18396, ZN => n18325);
   U2689 : AOI22_X1 port map( A1 => REGISTERS_31_6_port, A2 => n18322, B1 => 
                           REGISTERS_20_6_port, B2 => n18443, ZN => n18324);
   U2690 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n18480, B1 => 
                           REGISTERS_21_6_port, B2 => n18484, ZN => n18323);
   U2691 : NAND4_X1 port map( A1 => n18326, A2 => n18325, A3 => n18324, A4 => 
                           n18323, ZN => n18327);
   U2692 : NOR2_X1 port map( A1 => n18328, A2 => n18327, ZN => n18341);
   U2693 : AOI22_X1 port map( A1 => REGISTERS_7_6_port, A2 => n18458, B1 => 
                           REGISTERS_3_6_port, B2 => n18513, ZN => n18332);
   U2694 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n18427, B1 => 
                           REGISTERS_5_6_port, B2 => n18505, ZN => n18331);
   U2695 : AOI22_X1 port map( A1 => REGISTERS_6_6_port, A2 => n18465, B1 => 
                           REGISTERS_4_6_port, B2 => n18466, ZN => n18330);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n18503, B1 => 
                           REGISTERS_2_6_port, B2 => n18508, ZN => n18329);
   U2697 : NAND4_X1 port map( A1 => n18332, A2 => n18331, A3 => n18330, A4 => 
                           n18329, ZN => n18338);
   U2698 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n18427, B1 => 
                           REGISTERS_14_6_port, B2 => n18517, ZN => n18336);
   U2699 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n18506, B1 => 
                           REGISTERS_8_6_port, B2 => n18519, ZN => n18335);
   U2700 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n18518, B1 => 
                           REGISTERS_15_6_port, B2 => n18458, ZN => n18334);
   U2701 : AOI22_X1 port map( A1 => REGISTERS_10_6_port, A2 => n18508, B1 => 
                           REGISTERS_11_6_port, B2 => n18513, ZN => n18333);
   U2702 : NAND4_X1 port map( A1 => n18336, A2 => n18335, A3 => n18334, A4 => 
                           n18333, ZN => n18337);
   U2703 : AOI22_X1 port map( A1 => n18339, A2 => n18338, B1 => n18363, B2 => 
                           n18337, ZN => n18340);
   U2704 : OAI21_X1 port map( B1 => n18531, B2 => n18341, A => n18340, ZN => 
                           N391);
   U2705 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n18415, B1 => 
                           REGISTERS_30_5_port, B2 => n18449, ZN => n18346);
   U2706 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n18342, B1 => 
                           REGISTERS_24_5_port, B2 => n18448, ZN => n18345);
   U2707 : AOI22_X1 port map( A1 => REGISTERS_26_5_port, A2 => n18440, B1 => 
                           REGISTERS_29_5_port, B2 => n18420, ZN => n18344);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n18494, B1 => 
                           REGISTERS_27_5_port, B2 => n18477, ZN => n18343);
   U2709 : NAND4_X1 port map( A1 => n18346, A2 => n18345, A3 => n18344, A4 => 
                           n18343, ZN => n18353);
   U2710 : AOI22_X1 port map( A1 => REGISTERS_17_5_port, A2 => n18347, B1 => 
                           REGISTERS_22_5_port, B2 => n18441, ZN => n18351);
   U2711 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n18442, B1 => 
                           REGISTERS_28_5_port, B2 => n18482, ZN => n18350);
   U2712 : AOI22_X1 port map( A1 => REGISTERS_31_5_port, A2 => n18479, B1 => 
                           REGISTERS_18_5_port, B2 => n18493, ZN => n18349);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n18495, B1 => 
                           REGISTERS_19_5_port, B2 => n18491, ZN => n18348);
   U2714 : NAND4_X1 port map( A1 => n18351, A2 => n18350, A3 => n18349, A4 => 
                           n18348, ZN => n18352);
   U2715 : NOR2_X1 port map( A1 => n18353, A2 => n18352, ZN => n18367);
   U2716 : AOI22_X1 port map( A1 => REGISTERS_6_5_port, A2 => n18465, B1 => 
                           REGISTERS_7_5_port, B2 => n18458, ZN => n18357);
   U2717 : AOI22_X1 port map( A1 => REGISTERS_5_5_port, A2 => n18505, B1 => 
                           REGISTERS_4_5_port, B2 => n18466, ZN => n18356);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_2_5_port, A2 => n18516, B1 => 
                           REGISTERS_3_5_port, B2 => n18513, ZN => n18355);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n18459, B1 => 
                           REGISTERS_0_5_port, B2 => n18503, ZN => n18354);
   U2720 : NAND4_X1 port map( A1 => n18357, A2 => n18356, A3 => n18355, A4 => 
                           n18354, ZN => n18364);
   U2721 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n18519, B1 => 
                           REGISTERS_12_5_port, B2 => n18514, ZN => n18361);
   U2722 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n18427, B1 => 
                           REGISTERS_14_5_port, B2 => n18465, ZN => n18360);
   U2723 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n18513, B1 => 
                           REGISTERS_15_5_port, B2 => n18458, ZN => n18359);
   U2724 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n18457, B1 => 
                           REGISTERS_10_5_port, B2 => n18508, ZN => n18358);
   U2725 : NAND4_X1 port map( A1 => n18361, A2 => n18360, A3 => n18359, A4 => 
                           n18358, ZN => n18362);
   U2726 : AOI22_X1 port map( A1 => n18365, A2 => n18364, B1 => n18363, B2 => 
                           n18362, ZN => n18366);
   U2727 : OAI21_X1 port map( B1 => n18476, B2 => n18367, A => n18366, ZN => 
                           N390);
   U2728 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n18368, B1 => 
                           REGISTERS_21_4_port, B2 => n18484, ZN => n18372);
   U2729 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n18481, B1 => 
                           REGISTERS_17_4_port, B2 => n18480, ZN => n18371);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_26_4_port, A2 => n18490, B1 => 
                           REGISTERS_20_4_port, B2 => n18443, ZN => n18370);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n18496, B1 => 
                           REGISTERS_24_4_port, B2 => n18448, ZN => n18369);
   U2732 : NAND4_X1 port map( A1 => n18372, A2 => n18371, A3 => n18370, A4 => 
                           n18369, ZN => n18378);
   U2733 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n18482, B1 => 
                           REGISTERS_16_4_port, B2 => n18396, ZN => n18376);
   U2734 : AOI22_X1 port map( A1 => REGISTERS_22_4_port, A2 => n18441, B1 => 
                           REGISTERS_18_4_port, B2 => n18493, ZN => n18375);
   U2735 : AOI22_X1 port map( A1 => REGISTERS_19_4_port, A2 => n18491, B1 => 
                           REGISTERS_23_4_port, B2 => n18489, ZN => n18374);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_30_4_port, A2 => n18449, B1 => 
                           REGISTERS_31_4_port, B2 => n18479, ZN => n18373);
   U2737 : NAND4_X1 port map( A1 => n18376, A2 => n18375, A3 => n18374, A4 => 
                           n18373, ZN => n18377);
   U2738 : NOR2_X1 port map( A1 => n18378, A2 => n18377, ZN => n18391);
   U2739 : AOI22_X1 port map( A1 => REGISTERS_1_4_port, A2 => n18459, B1 => 
                           REGISTERS_4_4_port, B2 => n18466, ZN => n18382);
   U2740 : AOI22_X1 port map( A1 => REGISTERS_3_4_port, A2 => n18507, B1 => 
                           REGISTERS_6_4_port, B2 => n18456, ZN => n18381);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n18519, B1 => 
                           REGISTERS_5_4_port, B2 => n18505, ZN => n18380);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_2_4_port, A2 => n18467, B1 => 
                           REGISTERS_7_4_port, B2 => n18458, ZN => n18379);
   U2743 : NAND4_X1 port map( A1 => n18382, A2 => n18381, A3 => n18380, A4 => 
                           n18379, ZN => n18389);
   U2744 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n18459, B1 => 
                           REGISTERS_8_4_port, B2 => n18519, ZN => n18387);
   U2745 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n18520, B1 => 
                           REGISTERS_12_4_port, B2 => n18514, ZN => n18386);
   U2746 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n18383, B1 => 
                           REGISTERS_14_4_port, B2 => n18456, ZN => n18385);
   U2747 : AOI22_X1 port map( A1 => REGISTERS_13_4_port, A2 => n18505, B1 => 
                           REGISTERS_10_4_port, B2 => n18508, ZN => n18384);
   U2748 : NAND4_X1 port map( A1 => n18387, A2 => n18386, A3 => n18385, A4 => 
                           n18384, ZN => n18388);
   U2749 : AOI22_X1 port map( A1 => n18528, A2 => n18389, B1 => n18526, B2 => 
                           n18388, ZN => n18390);
   U2750 : OAI21_X1 port map( B1 => n18531, B2 => n18391, A => n18390, ZN => 
                           N389);
   U2751 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n18482, B1 => 
                           REGISTERS_30_3_port, B2 => n18449, ZN => n18395);
   U2752 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n18491, B1 => 
                           REGISTERS_24_3_port, B2 => n18448, ZN => n18394);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_22_3_port, A2 => n18478, B1 => 
                           REGISTERS_20_3_port, B2 => n18443, ZN => n18393);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_23_3_port, A2 => n18442, B1 => 
                           REGISTERS_25_3_port, B2 => n18496, ZN => n18392);
   U2755 : NAND4_X1 port map( A1 => n18395, A2 => n18394, A3 => n18393, A4 => 
                           n18392, ZN => n18402);
   U2756 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n18481, B1 => 
                           REGISTERS_16_3_port, B2 => n18396, ZN => n18400);
   U2757 : AOI22_X1 port map( A1 => REGISTERS_31_3_port, A2 => n18479, B1 => 
                           REGISTERS_27_3_port, B2 => n18477, ZN => n18399);
   U2758 : AOI22_X1 port map( A1 => REGISTERS_18_3_port, A2 => n18493, B1 => 
                           REGISTERS_21_3_port, B2 => n18484, ZN => n18398);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n18480, B1 => 
                           REGISTERS_26_3_port, B2 => n18490, ZN => n18397);
   U2760 : NAND4_X1 port map( A1 => n18400, A2 => n18399, A3 => n18398, A4 => 
                           n18397, ZN => n18401);
   U2761 : NOR2_X1 port map( A1 => n18402, A2 => n18401, ZN => n18414);
   U2762 : AOI22_X1 port map( A1 => REGISTERS_6_3_port, A2 => n18456, B1 => 
                           REGISTERS_4_3_port, B2 => n18466, ZN => n18406);
   U2763 : AOI22_X1 port map( A1 => REGISTERS_2_3_port, A2 => n18508, B1 => 
                           REGISTERS_3_3_port, B2 => n18513, ZN => n18405);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n18519, B1 => 
                           REGISTERS_5_3_port, B2 => n18505, ZN => n18404);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_7_3_port, A2 => n18504, B1 => 
                           REGISTERS_1_3_port, B2 => n18515, ZN => n18403);
   U2766 : NAND4_X1 port map( A1 => n18406, A2 => n18405, A3 => n18404, A4 => 
                           n18403, ZN => n18412);
   U2767 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n18427, B1 => 
                           REGISTERS_12_3_port, B2 => n18514, ZN => n18410);
   U2768 : AOI22_X1 port map( A1 => REGISTERS_14_3_port, A2 => n18456, B1 => 
                           REGISTERS_8_3_port, B2 => n18503, ZN => n18409);
   U2769 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n18513, B1 => 
                           REGISTERS_10_3_port, B2 => n18508, ZN => n18408);
   U2770 : AOI22_X1 port map( A1 => REGISTERS_15_3_port, A2 => n18458, B1 => 
                           REGISTERS_13_3_port, B2 => n18505, ZN => n18407);
   U2771 : NAND4_X1 port map( A1 => n18410, A2 => n18409, A3 => n18408, A4 => 
                           n18407, ZN => n18411);
   U2772 : AOI22_X1 port map( A1 => n18528, A2 => n18412, B1 => n18526, B2 => 
                           n18411, ZN => n18413);
   U2773 : OAI21_X1 port map( B1 => n18476, B2 => n18414, A => n18413, ZN => 
                           N388);
   U2774 : AOI22_X1 port map( A1 => REGISTERS_30_2_port, A2 => n18449, B1 => 
                           REGISTERS_31_2_port, B2 => n18479, ZN => n18419);
   U2775 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n18442, B1 => 
                           REGISTERS_28_2_port, B2 => n18482, ZN => n18418);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_18_2_port, A2 => n18493, B1 => 
                           REGISTERS_19_2_port, B2 => n18491, ZN => n18417);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n18415, B1 => 
                           REGISTERS_26_2_port, B2 => n18490, ZN => n18416);
   U2778 : NAND4_X1 port map( A1 => n18419, A2 => n18418, A3 => n18417, A4 => 
                           n18416, ZN => n18426);
   U2779 : AOI22_X1 port map( A1 => REGISTERS_22_2_port, A2 => n18478, B1 => 
                           REGISTERS_27_2_port, B2 => n18477, ZN => n18424);
   U2780 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n18494, B1 => 
                           REGISTERS_24_2_port, B2 => n18448, ZN => n18423);
   U2781 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n18480, B1 => 
                           REGISTERS_25_2_port, B2 => n18496, ZN => n18422);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n18495, B1 => 
                           REGISTERS_29_2_port, B2 => n18420, ZN => n18421);
   U2783 : NAND4_X1 port map( A1 => n18424, A2 => n18423, A3 => n18422, A4 => 
                           n18421, ZN => n18425);
   U2784 : NOR2_X1 port map( A1 => n18426, A2 => n18425, ZN => n18439);
   U2785 : AOI22_X1 port map( A1 => REGISTERS_6_2_port, A2 => n18517, B1 => 
                           REGISTERS_3_2_port, B2 => n18513, ZN => n18431);
   U2786 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n18505, B1 => 
                           REGISTERS_4_2_port, B2 => n18466, ZN => n18430);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n18520, B1 => 
                           REGISTERS_2_2_port, B2 => n18508, ZN => n18429);
   U2788 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n18427, B1 => 
                           REGISTERS_0_2_port, B2 => n18464, ZN => n18428);
   U2789 : NAND4_X1 port map( A1 => n18431, A2 => n18430, A3 => n18429, A4 => 
                           n18428, ZN => n18437);
   U2790 : AOI22_X1 port map( A1 => REGISTERS_10_2_port, A2 => n18516, B1 => 
                           REGISTERS_8_2_port, B2 => n18464, ZN => n18435);
   U2791 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n18504, B1 => 
                           REGISTERS_12_2_port, B2 => n18466, ZN => n18434);
   U2792 : AOI22_X1 port map( A1 => REGISTERS_13_2_port, A2 => n18457, B1 => 
                           REGISTERS_14_2_port, B2 => n18465, ZN => n18433);
   U2793 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n18515, B1 => 
                           REGISTERS_11_2_port, B2 => n18513, ZN => n18432);
   U2794 : NAND4_X1 port map( A1 => n18435, A2 => n18434, A3 => n18433, A4 => 
                           n18432, ZN => n18436);
   U2795 : AOI22_X1 port map( A1 => n18528, A2 => n18437, B1 => n18526, B2 => 
                           n18436, ZN => n18438);
   U2796 : OAI21_X1 port map( B1 => n18531, B2 => n18439, A => n18438, ZN => 
                           N387);
   U2797 : AOI22_X1 port map( A1 => REGISTERS_26_1_port, A2 => n18440, B1 => 
                           REGISTERS_21_1_port, B2 => n18484, ZN => n18447);
   U2798 : AOI22_X1 port map( A1 => REGISTERS_23_1_port, A2 => n18442, B1 => 
                           REGISTERS_22_1_port, B2 => n18441, ZN => n18446);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n18481, B1 => 
                           REGISTERS_28_1_port, B2 => n18482, ZN => n18445);
   U2800 : AOI22_X1 port map( A1 => REGISTERS_18_1_port, A2 => n18493, B1 => 
                           REGISTERS_20_1_port, B2 => n18443, ZN => n18444);
   U2801 : NAND4_X1 port map( A1 => n18447, A2 => n18446, A3 => n18445, A4 => 
                           n18444, ZN => n18455);
   U2802 : AOI22_X1 port map( A1 => REGISTERS_17_1_port, A2 => n18480, B1 => 
                           REGISTERS_27_1_port, B2 => n18477, ZN => n18453);
   U2803 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n18494, B1 => 
                           REGISTERS_31_1_port, B2 => n18479, ZN => n18452);
   U2804 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n18496, B1 => 
                           REGISTERS_19_1_port, B2 => n18491, ZN => n18451);
   U2805 : AOI22_X1 port map( A1 => REGISTERS_30_1_port, A2 => n18449, B1 => 
                           REGISTERS_24_1_port, B2 => n18448, ZN => n18450);
   U2806 : NAND4_X1 port map( A1 => n18453, A2 => n18452, A3 => n18451, A4 => 
                           n18450, ZN => n18454);
   U2807 : NOR2_X1 port map( A1 => n18455, A2 => n18454, ZN => n18475);
   U2808 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n18506, B1 => 
                           REGISTERS_0_1_port, B2 => n18503, ZN => n18463);
   U2809 : AOI22_X1 port map( A1 => REGISTERS_6_1_port, A2 => n18456, B1 => 
                           REGISTERS_3_1_port, B2 => n18507, ZN => n18462);
   U2810 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n18458, B1 => 
                           REGISTERS_5_1_port, B2 => n18457, ZN => n18461);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n18459, B1 => 
                           REGISTERS_2_1_port, B2 => n18516, ZN => n18460);
   U2812 : NAND4_X1 port map( A1 => n18463, A2 => n18462, A3 => n18461, A4 => 
                           n18460, ZN => n18473);
   U2813 : AOI22_X1 port map( A1 => REGISTERS_15_1_port, A2 => n18520, B1 => 
                           REGISTERS_8_1_port, B2 => n18464, ZN => n18471);
   U2814 : AOI22_X1 port map( A1 => REGISTERS_14_1_port, A2 => n18465, B1 => 
                           REGISTERS_9_1_port, B2 => n18515, ZN => n18470);
   U2815 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n18518, B1 => 
                           REGISTERS_11_1_port, B2 => n18507, ZN => n18469);
   U2816 : AOI22_X1 port map( A1 => REGISTERS_10_1_port, A2 => n18467, B1 => 
                           REGISTERS_12_1_port, B2 => n18466, ZN => n18468);
   U2817 : NAND4_X1 port map( A1 => n18471, A2 => n18470, A3 => n18469, A4 => 
                           n18468, ZN => n18472);
   U2818 : AOI22_X1 port map( A1 => n18528, A2 => n18473, B1 => n18526, B2 => 
                           n18472, ZN => n18474);
   U2819 : OAI21_X1 port map( B1 => n18476, B2 => n18475, A => n18474, ZN => 
                           N386);
   U2820 : AOI22_X1 port map( A1 => REGISTERS_22_0_port, A2 => n18478, B1 => 
                           REGISTERS_27_0_port, B2 => n18477, ZN => n18488);
   U2821 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n18480, B1 => 
                           REGISTERS_31_0_port, B2 => n18479, ZN => n18487);
   U2822 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n18482, B1 => 
                           REGISTERS_29_0_port, B2 => n18481, ZN => n18486);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_21_0_port, A2 => n18484, B1 => 
                           REGISTERS_30_0_port, B2 => n18483, ZN => n18485);
   U2824 : NAND4_X1 port map( A1 => n18488, A2 => n18487, A3 => n18486, A4 => 
                           n18485, ZN => n18502);
   U2825 : AOI22_X1 port map( A1 => REGISTERS_26_0_port, A2 => n18490, B1 => 
                           REGISTERS_23_0_port, B2 => n18489, ZN => n18500);
   U2826 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n18492, B1 => 
                           REGISTERS_19_0_port, B2 => n18491, ZN => n18499);
   U2827 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n18494, B1 => 
                           REGISTERS_18_0_port, B2 => n18493, ZN => n18498);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_25_0_port, A2 => n18496, B1 => 
                           REGISTERS_20_0_port, B2 => n18495, ZN => n18497);
   U2829 : NAND4_X1 port map( A1 => n18500, A2 => n18499, A3 => n18498, A4 => 
                           n18497, ZN => n18501);
   U2830 : NOR2_X1 port map( A1 => n18502, A2 => n18501, ZN => n18530);
   U2831 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n18504, B1 => 
                           REGISTERS_0_0_port, B2 => n18503, ZN => n18512);
   U2832 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n18505, B1 => 
                           REGISTERS_1_0_port, B2 => n18515, ZN => n18511);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n18506, B1 => 
                           REGISTERS_6_0_port, B2 => n18517, ZN => n18510);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_2_0_port, A2 => n18508, B1 => 
                           REGISTERS_3_0_port, B2 => n18507, ZN => n18509);
   U2835 : NAND4_X1 port map( A1 => n18512, A2 => n18511, A3 => n18510, A4 => 
                           n18509, ZN => n18527);
   U2836 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n18514, B1 => 
                           REGISTERS_11_0_port, B2 => n18513, ZN => n18524);
   U2837 : AOI22_X1 port map( A1 => REGISTERS_10_0_port, A2 => n18516, B1 => 
                           REGISTERS_9_0_port, B2 => n18515, ZN => n18523);
   U2838 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n18518, B1 => 
                           REGISTERS_14_0_port, B2 => n18517, ZN => n18522);
   U2839 : AOI22_X1 port map( A1 => REGISTERS_15_0_port, A2 => n18520, B1 => 
                           REGISTERS_8_0_port, B2 => n18519, ZN => n18521);
   U2840 : NAND4_X1 port map( A1 => n18524, A2 => n18523, A3 => n18522, A4 => 
                           n18521, ZN => n18525);
   U2841 : AOI22_X1 port map( A1 => n18528, A2 => n18527, B1 => n18526, B2 => 
                           n18525, ZN => n18529);
   U2842 : OAI21_X1 port map( B1 => n18531, B2 => n18530, A => n18529, ZN => 
                           N385);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ENABLE_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, curr_instruction_to_cu_i_31_port, 
      curr_instruction_to_cu_i_30_port, curr_instruction_to_cu_i_28_port, 
      curr_instruction_to_cu_i_27_port, curr_instruction_to_cu_i_26_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_18_port, curr_instruction_to_cu_i_17_port, 
      curr_instruction_to_cu_i_16_port, curr_instruction_to_cu_i_15_port, 
      curr_instruction_to_cu_i_14_port, curr_instruction_to_cu_i_13_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_5_port, curr_instruction_to_cu_i_4_port, 
      curr_instruction_to_cu_i_3_port, curr_instruction_to_cu_i_2_port, 
      curr_instruction_to_cu_i_1_port, curr_instruction_to_cu_i_0_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n131, cu_i_n127, 
      cu_i_n126, cu_i_n125, cu_i_n124, cu_i_n123, cu_i_n210, cu_i_n209, 
      cu_i_n145, cu_i_n26, cu_i_n25, cu_i_n23, cu_i_cw1_i_4_port, 
      cu_i_cw1_i_7_port, cu_i_cw1_i_8_port, cu_i_cw3_6_port, cu_i_cw2_5_port, 
      cu_i_cw2_6_port, cu_i_cw2_7_port, cu_i_cw2_8_port, cu_i_cw1_0_port, 
      cu_i_cw1_1_port, cu_i_cw1_2_port, cu_i_cw1_3_port, cu_i_cw1_4_port, 
      cu_i_cw1_5_port, cu_i_cw1_6_port, cu_i_cw1_7_port, cu_i_cw1_8_port, 
      cu_i_cw1_10_port, cu_i_cw1_11_port, cu_i_cw1_12_port, cu_i_N279, 
      cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, cu_i_N273, 
      cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, cu_i_cmd_alu_op_type_0_port, 
      cu_i_cmd_alu_op_type_1_port, cu_i_cmd_alu_op_type_2_port, 
      cu_i_cmd_alu_op_type_3_port, cu_i_cmd_word_1_port, cu_i_cmd_word_3_port, 
      cu_i_cmd_word_4_port, cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, 
      cu_i_cmd_word_8_port, cu_i_next_stall, cu_i_next_val_counter_mul_0_port, 
      cu_i_next_val_counter_mul_1_port, cu_i_next_val_counter_mul_2_port, 
      cu_i_next_val_counter_mul_3_port, datapath_i_data_from_alu_i_0_port, 
      datapath_i_data_from_alu_i_1_port, datapath_i_data_from_alu_i_2_port, 
      datapath_i_data_from_alu_i_3_port, datapath_i_data_from_alu_i_4_port, 
      datapath_i_data_from_alu_i_5_port, datapath_i_data_from_alu_i_6_port, 
      datapath_i_data_from_alu_i_7_port, datapath_i_data_from_alu_i_8_port, 
      datapath_i_data_from_alu_i_9_port, datapath_i_data_from_alu_i_10_port, 
      datapath_i_data_from_alu_i_11_port, datapath_i_data_from_alu_i_12_port, 
      datapath_i_data_from_alu_i_13_port, datapath_i_data_from_alu_i_14_port, 
      datapath_i_data_from_alu_i_15_port, datapath_i_data_from_alu_i_16_port, 
      datapath_i_data_from_alu_i_17_port, datapath_i_data_from_alu_i_18_port, 
      datapath_i_data_from_alu_i_19_port, datapath_i_data_from_alu_i_20_port, 
      datapath_i_data_from_alu_i_21_port, datapath_i_data_from_alu_i_22_port, 
      datapath_i_data_from_alu_i_23_port, datapath_i_data_from_alu_i_24_port, 
      datapath_i_data_from_alu_i_25_port, datapath_i_data_from_alu_i_26_port, 
      datapath_i_data_from_alu_i_27_port, datapath_i_data_from_alu_i_28_port, 
      datapath_i_data_from_alu_i_29_port, datapath_i_data_from_alu_i_30_port, 
      datapath_i_data_from_alu_i_31_port, datapath_i_data_from_memory_i_0_port,
      datapath_i_data_from_memory_i_1_port, 
      datapath_i_data_from_memory_i_2_port, 
      datapath_i_data_from_memory_i_3_port, 
      datapath_i_data_from_memory_i_4_port, 
      datapath_i_data_from_memory_i_5_port, 
      datapath_i_data_from_memory_i_6_port, 
      datapath_i_data_from_memory_i_7_port, 
      datapath_i_data_from_memory_i_8_port, 
      datapath_i_data_from_memory_i_9_port, 
      datapath_i_data_from_memory_i_10_port, 
      datapath_i_data_from_memory_i_11_port, 
      datapath_i_data_from_memory_i_12_port, 
      datapath_i_data_from_memory_i_13_port, 
      datapath_i_data_from_memory_i_14_port, 
      datapath_i_data_from_memory_i_15_port, 
      datapath_i_data_from_memory_i_16_port, 
      datapath_i_data_from_memory_i_17_port, 
      datapath_i_data_from_memory_i_18_port, 
      datapath_i_data_from_memory_i_19_port, 
      datapath_i_data_from_memory_i_20_port, 
      datapath_i_data_from_memory_i_21_port, 
      datapath_i_data_from_memory_i_22_port, 
      datapath_i_data_from_memory_i_23_port, 
      datapath_i_data_from_memory_i_24_port, 
      datapath_i_data_from_memory_i_25_port, 
      datapath_i_data_from_memory_i_26_port, 
      datapath_i_data_from_memory_i_27_port, 
      datapath_i_data_from_memory_i_28_port, 
      datapath_i_data_from_memory_i_29_port, 
      datapath_i_data_from_memory_i_30_port, 
      datapath_i_data_from_memory_i_31_port, datapath_i_value_to_mem_i_0_port, 
      datapath_i_value_to_mem_i_1_port, datapath_i_value_to_mem_i_2_port, 
      datapath_i_value_to_mem_i_3_port, datapath_i_value_to_mem_i_4_port, 
      datapath_i_value_to_mem_i_5_port, datapath_i_value_to_mem_i_6_port, 
      datapath_i_value_to_mem_i_7_port, datapath_i_value_to_mem_i_8_port, 
      datapath_i_value_to_mem_i_9_port, datapath_i_value_to_mem_i_10_port, 
      datapath_i_value_to_mem_i_11_port, datapath_i_value_to_mem_i_12_port, 
      datapath_i_value_to_mem_i_13_port, datapath_i_value_to_mem_i_14_port, 
      datapath_i_value_to_mem_i_15_port, datapath_i_value_to_mem_i_16_port, 
      datapath_i_value_to_mem_i_17_port, datapath_i_value_to_mem_i_18_port, 
      datapath_i_value_to_mem_i_19_port, datapath_i_value_to_mem_i_20_port, 
      datapath_i_value_to_mem_i_21_port, datapath_i_value_to_mem_i_22_port, 
      datapath_i_value_to_mem_i_23_port, datapath_i_value_to_mem_i_24_port, 
      datapath_i_value_to_mem_i_25_port, datapath_i_value_to_mem_i_26_port, 
      datapath_i_value_to_mem_i_27_port, datapath_i_value_to_mem_i_28_port, 
      datapath_i_value_to_mem_i_29_port, datapath_i_value_to_mem_i_30_port, 
      datapath_i_value_to_mem_i_31_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, datapath_i_val_immediate_i_0_port, 
      datapath_i_val_immediate_i_1_port, datapath_i_val_immediate_i_2_port, 
      datapath_i_val_immediate_i_3_port, datapath_i_val_immediate_i_4_port, 
      datapath_i_val_immediate_i_5_port, datapath_i_val_immediate_i_6_port, 
      datapath_i_val_immediate_i_7_port, datapath_i_val_immediate_i_8_port, 
      datapath_i_val_immediate_i_9_port, datapath_i_val_immediate_i_10_port, 
      datapath_i_val_immediate_i_11_port, datapath_i_val_immediate_i_12_port, 
      datapath_i_val_immediate_i_13_port, datapath_i_val_immediate_i_14_port, 
      datapath_i_val_immediate_i_15_port, datapath_i_val_immediate_i_16_port, 
      datapath_i_val_immediate_i_17_port, datapath_i_val_immediate_i_18_port, 
      datapath_i_val_immediate_i_19_port, datapath_i_val_immediate_i_20_port, 
      datapath_i_val_immediate_i_21_port, datapath_i_val_immediate_i_22_port, 
      datapath_i_val_immediate_i_23_port, datapath_i_val_immediate_i_24_port, 
      datapath_i_val_immediate_i_25_port, datapath_i_val_b_i_0_port, 
      datapath_i_val_b_i_1_port, datapath_i_val_b_i_2_port, 
      datapath_i_val_b_i_3_port, datapath_i_val_b_i_4_port, 
      datapath_i_val_b_i_5_port, datapath_i_val_b_i_6_port, 
      datapath_i_val_b_i_7_port, datapath_i_val_b_i_8_port, 
      datapath_i_val_b_i_9_port, datapath_i_val_b_i_10_port, 
      datapath_i_val_b_i_11_port, datapath_i_val_b_i_12_port, 
      datapath_i_val_b_i_13_port, datapath_i_val_b_i_14_port, 
      datapath_i_val_b_i_15_port, datapath_i_val_b_i_16_port, 
      datapath_i_val_b_i_17_port, datapath_i_val_b_i_18_port, 
      datapath_i_val_b_i_19_port, datapath_i_val_b_i_20_port, 
      datapath_i_val_b_i_21_port, datapath_i_val_b_i_22_port, 
      datapath_i_val_b_i_23_port, datapath_i_val_b_i_24_port, 
      datapath_i_val_b_i_25_port, datapath_i_val_b_i_26_port, 
      datapath_i_val_b_i_27_port, datapath_i_val_b_i_28_port, 
      datapath_i_val_b_i_29_port, datapath_i_val_b_i_30_port, 
      datapath_i_val_b_i_31_port, datapath_i_val_a_i_0_port, 
      datapath_i_val_a_i_1_port, datapath_i_val_a_i_2_port, 
      datapath_i_val_a_i_3_port, datapath_i_val_a_i_4_port, 
      datapath_i_val_a_i_5_port, datapath_i_val_a_i_6_port, 
      datapath_i_val_a_i_7_port, datapath_i_val_a_i_8_port, 
      datapath_i_val_a_i_9_port, datapath_i_val_a_i_10_port, 
      datapath_i_val_a_i_11_port, datapath_i_val_a_i_12_port, 
      datapath_i_val_a_i_13_port, datapath_i_val_a_i_14_port, 
      datapath_i_val_a_i_15_port, datapath_i_val_a_i_16_port, 
      datapath_i_val_a_i_17_port, datapath_i_val_a_i_18_port, 
      datapath_i_val_a_i_19_port, datapath_i_val_a_i_20_port, 
      datapath_i_val_a_i_21_port, datapath_i_val_a_i_22_port, 
      datapath_i_val_a_i_23_port, datapath_i_val_a_i_24_port, 
      datapath_i_val_a_i_25_port, datapath_i_val_a_i_26_port, 
      datapath_i_val_a_i_27_port, datapath_i_val_a_i_28_port, 
      datapath_i_val_a_i_29_port, datapath_i_val_a_i_30_port, 
      datapath_i_val_a_i_31_port, datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_5_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_7_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_9_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_11_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_13_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_15_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_17_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_19_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_21_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_23_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_25_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_27_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_29_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, 
      datapath_i_new_pc_value_mem_stage_i_31_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_n69, 
      datapath_i_fetch_stage_dp_n68, datapath_i_fetch_stage_dp_n67, 
      datapath_i_fetch_stage_dp_n66, datapath_i_fetch_stage_dp_n65, 
      datapath_i_fetch_stage_dp_n64, datapath_i_fetch_stage_dp_n63, 
      datapath_i_fetch_stage_dp_n62, datapath_i_fetch_stage_dp_n61, 
      datapath_i_fetch_stage_dp_n60, datapath_i_fetch_stage_dp_n59, 
      datapath_i_fetch_stage_dp_n58, datapath_i_fetch_stage_dp_n57, 
      datapath_i_fetch_stage_dp_n56, datapath_i_fetch_stage_dp_n55, 
      datapath_i_fetch_stage_dp_n54, datapath_i_fetch_stage_dp_n53, 
      datapath_i_fetch_stage_dp_n52, datapath_i_fetch_stage_dp_n51, 
      datapath_i_fetch_stage_dp_n50, datapath_i_fetch_stage_dp_n49, 
      datapath_i_fetch_stage_dp_n48, datapath_i_fetch_stage_dp_n47, 
      datapath_i_fetch_stage_dp_n46, datapath_i_fetch_stage_dp_n45, 
      datapath_i_fetch_stage_dp_n44, datapath_i_fetch_stage_dp_n43, 
      datapath_i_fetch_stage_dp_n42, datapath_i_fetch_stage_dp_n41, 
      datapath_i_fetch_stage_dp_n40, datapath_i_fetch_stage_dp_n39, 
      datapath_i_fetch_stage_dp_n38, datapath_i_fetch_stage_dp_n37, 
      datapath_i_fetch_stage_dp_n36, datapath_i_fetch_stage_dp_n35, 
      datapath_i_fetch_stage_dp_n34, datapath_i_fetch_stage_dp_n33, 
      datapath_i_fetch_stage_dp_n32, datapath_i_fetch_stage_dp_n31, 
      datapath_i_fetch_stage_dp_n30, datapath_i_fetch_stage_dp_n29, 
      datapath_i_fetch_stage_dp_n28, datapath_i_fetch_stage_dp_n27, 
      datapath_i_fetch_stage_dp_n26, datapath_i_fetch_stage_dp_n25, 
      datapath_i_fetch_stage_dp_n24, datapath_i_fetch_stage_dp_n23, 
      datapath_i_fetch_stage_dp_n22, datapath_i_fetch_stage_dp_n21, 
      datapath_i_fetch_stage_dp_n20, datapath_i_fetch_stage_dp_n19, 
      datapath_i_fetch_stage_dp_n18, datapath_i_fetch_stage_dp_n17, 
      datapath_i_fetch_stage_dp_n16, datapath_i_fetch_stage_dp_n15, 
      datapath_i_fetch_stage_dp_n14, datapath_i_fetch_stage_dp_n13, 
      datapath_i_fetch_stage_dp_n12, datapath_i_fetch_stage_dp_n11, 
      datapath_i_fetch_stage_dp_n10, datapath_i_fetch_stage_dp_n9, 
      datapath_i_fetch_stage_dp_n4, datapath_i_fetch_stage_dp_n3, 
      datapath_i_fetch_stage_dp_n2, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port, datapath_i_fetch_stage_dp_N6, 
      datapath_i_fetch_stage_dp_N5, datapath_i_decode_stage_dp_n78, 
      datapath_i_decode_stage_dp_n43, datapath_i_decode_stage_dp_n42, 
      datapath_i_decode_stage_dp_n41, datapath_i_decode_stage_dp_n40, 
      datapath_i_decode_stage_dp_n39, datapath_i_decode_stage_dp_n38, 
      datapath_i_decode_stage_dp_n37, datapath_i_decode_stage_dp_n36, 
      datapath_i_decode_stage_dp_n35, datapath_i_decode_stage_dp_n34, 
      datapath_i_decode_stage_dp_n33, datapath_i_decode_stage_dp_n32, 
      datapath_i_decode_stage_dp_n31, datapath_i_decode_stage_dp_n30, 
      datapath_i_decode_stage_dp_n29, datapath_i_decode_stage_dp_n28, 
      datapath_i_decode_stage_dp_n27, datapath_i_decode_stage_dp_n26, 
      datapath_i_decode_stage_dp_n25, datapath_i_decode_stage_dp_n24, 
      datapath_i_decode_stage_dp_n23, datapath_i_decode_stage_dp_n22, 
      datapath_i_decode_stage_dp_n21, datapath_i_decode_stage_dp_n20, 
      datapath_i_decode_stage_dp_n19, datapath_i_decode_stage_dp_n18, 
      datapath_i_decode_stage_dp_n17, datapath_i_decode_stage_dp_n16, 
      datapath_i_decode_stage_dp_n15, datapath_i_decode_stage_dp_n14, 
      datapath_i_decode_stage_dp_n13, datapath_i_decode_stage_dp_n12, 
      datapath_i_decode_stage_dp_pc_delay3_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_1_port, 
      datapath_i_decode_stage_dp_pc_delay2_2_port, 
      datapath_i_decode_stage_dp_pc_delay2_3_port, 
      datapath_i_decode_stage_dp_pc_delay2_4_port, 
      datapath_i_decode_stage_dp_pc_delay2_5_port, 
      datapath_i_decode_stage_dp_pc_delay2_6_port, 
      datapath_i_decode_stage_dp_pc_delay2_7_port, 
      datapath_i_decode_stage_dp_pc_delay2_8_port, 
      datapath_i_decode_stage_dp_pc_delay2_9_port, 
      datapath_i_decode_stage_dp_pc_delay2_10_port, 
      datapath_i_decode_stage_dp_pc_delay2_11_port, 
      datapath_i_decode_stage_dp_pc_delay2_12_port, 
      datapath_i_decode_stage_dp_pc_delay2_13_port, 
      datapath_i_decode_stage_dp_pc_delay2_14_port, 
      datapath_i_decode_stage_dp_pc_delay2_15_port, 
      datapath_i_decode_stage_dp_pc_delay2_16_port, 
      datapath_i_decode_stage_dp_pc_delay2_17_port, 
      datapath_i_decode_stage_dp_pc_delay2_18_port, 
      datapath_i_decode_stage_dp_pc_delay2_19_port, 
      datapath_i_decode_stage_dp_pc_delay2_20_port, 
      datapath_i_decode_stage_dp_pc_delay2_21_port, 
      datapath_i_decode_stage_dp_pc_delay2_22_port, 
      datapath_i_decode_stage_dp_pc_delay2_23_port, 
      datapath_i_decode_stage_dp_pc_delay2_24_port, 
      datapath_i_decode_stage_dp_pc_delay2_25_port, 
      datapath_i_decode_stage_dp_pc_delay2_26_port, 
      datapath_i_decode_stage_dp_pc_delay2_27_port, 
      datapath_i_decode_stage_dp_pc_delay2_28_port, 
      datapath_i_decode_stage_dp_pc_delay2_29_port, 
      datapath_i_decode_stage_dp_pc_delay2_30_port, 
      datapath_i_decode_stage_dp_pc_delay2_31_port, 
      datapath_i_decode_stage_dp_pc_delay2_32_port, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_0_port, 
      datapath_i_decode_stage_dp_address_rf_write_1_port, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_decode_stage_dp_address_rf_write_3_port, 
      datapath_i_decode_stage_dp_address_rf_write_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_out_0_port, 
      datapath_i_execute_stage_dp_alu_out_1_port, 
      datapath_i_execute_stage_dp_alu_out_2_port, 
      datapath_i_execute_stage_dp_alu_out_3_port, 
      datapath_i_execute_stage_dp_alu_out_4_port, 
      datapath_i_execute_stage_dp_alu_out_5_port, 
      datapath_i_execute_stage_dp_alu_out_6_port, 
      datapath_i_execute_stage_dp_alu_out_7_port, 
      datapath_i_execute_stage_dp_alu_out_8_port, 
      datapath_i_execute_stage_dp_alu_out_9_port, 
      datapath_i_execute_stage_dp_alu_out_10_port, 
      datapath_i_execute_stage_dp_alu_out_11_port, 
      datapath_i_execute_stage_dp_alu_out_12_port, 
      datapath_i_execute_stage_dp_alu_out_13_port, 
      datapath_i_execute_stage_dp_alu_out_14_port, 
      datapath_i_execute_stage_dp_alu_out_15_port, 
      datapath_i_execute_stage_dp_alu_out_16_port, 
      datapath_i_execute_stage_dp_alu_out_17_port, 
      datapath_i_execute_stage_dp_alu_out_18_port, 
      datapath_i_execute_stage_dp_alu_out_19_port, 
      datapath_i_execute_stage_dp_alu_out_20_port, 
      datapath_i_execute_stage_dp_alu_out_21_port, 
      datapath_i_execute_stage_dp_alu_out_22_port, 
      datapath_i_execute_stage_dp_alu_out_23_port, 
      datapath_i_execute_stage_dp_alu_out_24_port, 
      datapath_i_execute_stage_dp_alu_out_25_port, 
      datapath_i_execute_stage_dp_alu_out_26_port, 
      datapath_i_execute_stage_dp_alu_out_27_port, 
      datapath_i_execute_stage_dp_alu_out_28_port, 
      datapath_i_execute_stage_dp_alu_out_29_port, 
      datapath_i_execute_stage_dp_alu_out_30_port, 
      datapath_i_execute_stage_dp_alu_out_31_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, 
      datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
      datapath_i_memory_stage_dp_n2, datapath_i_memory_stage_dp_data_ir_0_port,
      datapath_i_memory_stage_dp_data_ir_1_port, 
      datapath_i_memory_stage_dp_data_ir_2_port, 
      datapath_i_memory_stage_dp_data_ir_3_port, 
      datapath_i_memory_stage_dp_data_ir_4_port, 
      datapath_i_memory_stage_dp_data_ir_5_port, 
      datapath_i_memory_stage_dp_data_ir_6_port, 
      datapath_i_memory_stage_dp_data_ir_7_port, 
      datapath_i_memory_stage_dp_data_ir_8_port, 
      datapath_i_memory_stage_dp_data_ir_9_port, 
      datapath_i_memory_stage_dp_data_ir_10_port, 
      datapath_i_memory_stage_dp_data_ir_11_port, 
      datapath_i_memory_stage_dp_data_ir_12_port, 
      datapath_i_memory_stage_dp_data_ir_13_port, 
      datapath_i_memory_stage_dp_data_ir_14_port, 
      datapath_i_memory_stage_dp_data_ir_15_port, 
      datapath_i_memory_stage_dp_data_ir_16_port, 
      datapath_i_memory_stage_dp_data_ir_17_port, 
      datapath_i_memory_stage_dp_data_ir_18_port, 
      datapath_i_memory_stage_dp_data_ir_19_port, 
      datapath_i_memory_stage_dp_data_ir_20_port, 
      datapath_i_memory_stage_dp_data_ir_21_port, 
      datapath_i_memory_stage_dp_data_ir_22_port, 
      datapath_i_memory_stage_dp_data_ir_23_port, 
      datapath_i_memory_stage_dp_data_ir_24_port, 
      datapath_i_memory_stage_dp_data_ir_25_port, 
      datapath_i_memory_stage_dp_data_ir_26_port, 
      datapath_i_memory_stage_dp_data_ir_27_port, 
      datapath_i_memory_stage_dp_data_ir_28_port, 
      datapath_i_memory_stage_dp_data_ir_29_port, 
      datapath_i_memory_stage_dp_data_ir_30_port, 
      datapath_i_memory_stage_dp_data_ir_31_port, n309, n311, n691, n697, n699,
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n737, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n756, 
      n758, n759, n760, n761, n762, n763, n764, n1152, n2319, n4276, n4277, 
      n4278, n4279, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, 
      n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, 
      n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, 
      n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, 
      n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, 
      n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, 
      n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, 
      n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, 
      n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, 
      n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
      n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, 
      n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, 
      n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
      n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, 
      n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, 
      n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, 
      n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, 
      n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
      n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, 
      n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, 
      n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
      n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
      n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, 
      n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, 
      n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, 
      n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, 
      n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, 
      n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, 
      n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, 
      n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, 
      n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, 
      n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, 
      n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, 
      n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, 
      n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, 
      n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, 
      n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, 
      n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, 
      n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, 
      n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, 
      DRAM_ENABLE_port, n4679, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, 
      n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, 
      n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, 
      n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, 
      n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, 
      n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, 
      n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, 
      n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, 
      n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, 
      n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, 
      n_1797, n_1798 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   DRAM_ENABLE <= DRAM_ENABLE_port;
   
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_next_val_counter_mul_3_port);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_next_val_counter_mul_0_port);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => cu_i_n145, Q => 
                           cu_i_next_stall);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           ADD_WR(3) => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           ADD_WR(2) => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ADD_WR(1) => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ADD_WR(0) => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n12, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n43, OUT1(31) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
                           OUT1(30) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
                           OUT1(29) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
                           OUT1(28) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
                           OUT1(27) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
                           OUT1(26) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
                           OUT1(25) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
                           OUT1(24) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
                           OUT1(23) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
                           OUT1(22) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
                           OUT1(21) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
                           OUT1(20) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
                           OUT1(19) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
                           OUT1(18) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
                           OUT1(17) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
                           OUT1(16) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
                           OUT1(15) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
                           OUT1(14) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
                           OUT1(13) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
                           OUT1(12) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
                           OUT1(11) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
                           OUT1(10) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
                           OUT1(9) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
                           OUT1(8) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
                           OUT1(7) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
                           OUT1(6) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
                           OUT1(5) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
                           OUT1(4) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
                           OUT1(3) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
                           OUT1(2) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
                           OUT1(1) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
                           OUT1(0) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
                           OUT2(31) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
                           OUT2(30) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
                           OUT2(29) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
                           OUT2(28) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
                           OUT2(27) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
                           OUT2(26) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
                           OUT2(25) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
                           OUT2(24) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
                           OUT2(23) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
                           OUT2(22) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
                           OUT2(21) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
                           OUT2(20) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
                           OUT2(19) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
                           OUT2(18) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
                           OUT2(17) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
                           OUT2(16) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
                           OUT2(15) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
                           OUT2(14) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
                           OUT2(13) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
                           OUT2(12) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
                           OUT2(11) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
                           OUT2(10) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
                           OUT2(9) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
                           OUT2(8) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
                           OUT2(7) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
                           OUT2(6) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
                           OUT2(5) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
                           OUT2(4) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
                           OUT2(3) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
                           OUT2(2) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
                           OUT2(1) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
                           OUT2(0) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
                           RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_1413, mul_exeception => 
                           n_1414, FUNC(0) => n4281, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_1415, 
                           OUTALU(31) => 
                           datapath_i_execute_stage_dp_alu_out_31_port, 
                           OUTALU(30) => 
                           datapath_i_execute_stage_dp_alu_out_30_port, 
                           OUTALU(29) => 
                           datapath_i_execute_stage_dp_alu_out_29_port, 
                           OUTALU(28) => 
                           datapath_i_execute_stage_dp_alu_out_28_port, 
                           OUTALU(27) => 
                           datapath_i_execute_stage_dp_alu_out_27_port, 
                           OUTALU(26) => 
                           datapath_i_execute_stage_dp_alu_out_26_port, 
                           OUTALU(25) => 
                           datapath_i_execute_stage_dp_alu_out_25_port, 
                           OUTALU(24) => 
                           datapath_i_execute_stage_dp_alu_out_24_port, 
                           OUTALU(23) => 
                           datapath_i_execute_stage_dp_alu_out_23_port, 
                           OUTALU(22) => 
                           datapath_i_execute_stage_dp_alu_out_22_port, 
                           OUTALU(21) => 
                           datapath_i_execute_stage_dp_alu_out_21_port, 
                           OUTALU(20) => 
                           datapath_i_execute_stage_dp_alu_out_20_port, 
                           OUTALU(19) => 
                           datapath_i_execute_stage_dp_alu_out_19_port, 
                           OUTALU(18) => 
                           datapath_i_execute_stage_dp_alu_out_18_port, 
                           OUTALU(17) => 
                           datapath_i_execute_stage_dp_alu_out_17_port, 
                           OUTALU(16) => 
                           datapath_i_execute_stage_dp_alu_out_16_port, 
                           OUTALU(15) => 
                           datapath_i_execute_stage_dp_alu_out_15_port, 
                           OUTALU(14) => 
                           datapath_i_execute_stage_dp_alu_out_14_port, 
                           OUTALU(13) => 
                           datapath_i_execute_stage_dp_alu_out_13_port, 
                           OUTALU(12) => 
                           datapath_i_execute_stage_dp_alu_out_12_port, 
                           OUTALU(11) => 
                           datapath_i_execute_stage_dp_alu_out_11_port, 
                           OUTALU(10) => 
                           datapath_i_execute_stage_dp_alu_out_10_port, 
                           OUTALU(9) => 
                           datapath_i_execute_stage_dp_alu_out_9_port, 
                           OUTALU(8) => 
                           datapath_i_execute_stage_dp_alu_out_8_port, 
                           OUTALU(7) => 
                           datapath_i_execute_stage_dp_alu_out_7_port, 
                           OUTALU(6) => 
                           datapath_i_execute_stage_dp_alu_out_6_port, 
                           OUTALU(5) => 
                           datapath_i_execute_stage_dp_alu_out_5_port, 
                           OUTALU(4) => 
                           datapath_i_execute_stage_dp_alu_out_4_port, 
                           OUTALU(3) => 
                           datapath_i_execute_stage_dp_alu_out_3_port, 
                           OUTALU(2) => 
                           datapath_i_execute_stage_dp_alu_out_2_port, 
                           OUTALU(1) => 
                           datapath_i_execute_stage_dp_alu_out_1_port, 
                           OUTALU(0) => 
                           datapath_i_execute_stage_dp_alu_out_0_port, rst_BAR 
                           => RST);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n309, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n4677, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n4677, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n4677, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n4677, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n4677, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n309, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n4677, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n4677, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n4677, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n309, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n309, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n4677, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n4677, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n309, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n309, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n4677, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n4677, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n4677, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n4677, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n4677, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n4677, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n309, Z =>
                           DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n309, Z =>
                           DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n4677, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n4677, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n4677, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n309, Z =>
                           DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n4677, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n4677, Z 
                           => DRAM_ADDRESS_2_port);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_9_port, EN => n4679, Z => 
                           DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_31_port, EN => n4679, Z =>
                           DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_30_port, EN => n4679, Z =>
                           DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_29_port, EN => n4679, Z =>
                           DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_28_port, EN => n4679, Z =>
                           DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_27_port, EN => n4679, Z =>
                           DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_26_port, EN => n4679, Z =>
                           DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_25_port, EN => n4679, Z =>
                           DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_24_port, EN => n4679, Z =>
                           DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_23_port, EN => n4679, Z =>
                           DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_22_port, EN => n4679, Z =>
                           DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_21_port, EN => n4679, Z =>
                           DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_20_port, EN => n4679, Z =>
                           DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_19_port, EN => n4679, Z =>
                           DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_18_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_17_port, EN => n4679, Z =>
                           DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_16_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_15_port, EN => n4679, Z =>
                           DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_14_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_13_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_12_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_11_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_10_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_8_port, EN => n4679, Z => 
                           DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_7_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_6_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_5_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_4_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_3_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_2_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_1_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_0_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(0));
   cu_i_e_reg_D_I_0_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_0_port, QN => 
                           n_1416);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n4675, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n4676, D => datapath_i_n18, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n4675, D => datapath_i_n17, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n4676, D => datapath_i_n16, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n4675, D => datapath_i_n15, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n4676, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n4676, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n4674, D => datapath_i_n18, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n4674, D => datapath_i_n17, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n4674, D => datapath_i_n16, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n4674, D => datapath_i_n15, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n4674, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_16_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_17_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_18_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_19_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n4674, D => 
                           curr_instruction_to_cu_i_20_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n4674, D => datapath_i_n13, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n4674, D => datapath_i_n12, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n4674, D => datapath_i_n11, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n4674, D => datapath_i_n10, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n4674, D => datapath_i_n9, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   cu_i_wb_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n4282, CK => CLK, RN => RST
                           , Q => cu_i_cw3_6_port, QN => n_1417);
   cu_i_wb_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n131, CK => CLK, RN =>
                           RST, Q => n_1418, QN => n699);
   cu_i_m_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_8_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_8_port, QN => n_1419);
   cu_i_m_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_7_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_7_port, QN => n_1420);
   cu_i_m_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n127, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_6_port, QN => n_1421);
   cu_i_m_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n126, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_5_port, QN => n4673);
   cu_i_m_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_4_port, CK => CLK
                           , RN => RST, Q => n_1422, QN => n756);
   cu_i_e_reg_D_I_13_Q_reg : DFFR_X1 port map( D => n4676, CK => CLK, RN => RST
                           , Q => n_1423, QN => n2319);
   cu_i_e_reg_D_I_12_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_12_port, QN => n_1424)
                           ;
   cu_i_e_reg_D_I_11_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_11_port, QN => n_1425)
                           ;
   cu_i_e_reg_D_I_10_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_10_port, QN => n_1426)
                           ;
   cu_i_e_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_8_port, QN => n_1427);
   cu_i_e_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_7_port, QN => n_1428);
   cu_i_e_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n311, CK => CLK, RN => RST, 
                           Q => cu_i_cw1_6_port, QN => n_1429);
   cu_i_e_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_1_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_5_port, QN => n_1430);
   cu_i_e_reg_D_I_4_Q_reg : DFFR_X1 port map( D => n1152, CK => CLK, RN => RST,
                           Q => cu_i_cw1_4_port, QN => n_1431);
   cu_i_e_reg_D_I_3_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_3_port, QN => 
                           n_1432);
   cu_i_e_reg_D_I_2_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_2_port, QN => 
                           n_1433);
   cu_i_e_reg_D_I_1_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_1_port, QN => 
                           n_1434);
   datapath_i_memory_stage_dp_delay_regg_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_31_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_31_port, QN 
                           => n_1435);
   datapath_i_memory_stage_dp_delay_regg_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_30_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_30_port, QN 
                           => n_1436);
   datapath_i_memory_stage_dp_delay_regg_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_29_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_29_port, QN 
                           => n_1437);
   datapath_i_memory_stage_dp_delay_regg_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_28_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_28_port, QN 
                           => n_1438);
   datapath_i_memory_stage_dp_delay_regg_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_27_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_27_port, QN 
                           => n_1439);
   datapath_i_memory_stage_dp_delay_regg_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_26_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_26_port, QN 
                           => n_1440);
   datapath_i_memory_stage_dp_delay_regg_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_25_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_25_port, QN 
                           => n_1441);
   datapath_i_memory_stage_dp_delay_regg_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_24_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_24_port, QN 
                           => n_1442);
   datapath_i_memory_stage_dp_delay_regg_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_23_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_23_port, QN 
                           => n_1443);
   datapath_i_memory_stage_dp_delay_regg_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_22_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_22_port, QN 
                           => n_1444);
   datapath_i_memory_stage_dp_delay_regg_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_21_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_21_port, QN 
                           => n_1445);
   datapath_i_memory_stage_dp_delay_regg_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_20_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_20_port, QN 
                           => n_1446);
   datapath_i_memory_stage_dp_delay_regg_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_19_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_19_port, QN 
                           => n_1447);
   datapath_i_memory_stage_dp_delay_regg_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_18_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_18_port, QN 
                           => n_1448);
   datapath_i_memory_stage_dp_delay_regg_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_17_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_17_port, QN 
                           => n_1449);
   datapath_i_memory_stage_dp_delay_regg_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_16_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_16_port, QN 
                           => n_1450);
   datapath_i_memory_stage_dp_delay_regg_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_15_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_15_port, QN 
                           => n_1451);
   datapath_i_memory_stage_dp_delay_regg_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_14_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_14_port, QN 
                           => n_1452);
   datapath_i_memory_stage_dp_delay_regg_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_13_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_13_port, QN 
                           => n_1453);
   datapath_i_memory_stage_dp_delay_regg_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_12_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_12_port, QN 
                           => n_1454);
   datapath_i_memory_stage_dp_delay_regg_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_11_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_11_port, QN 
                           => n_1455);
   datapath_i_memory_stage_dp_delay_regg_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_10_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_10_port, QN 
                           => n_1456);
   datapath_i_memory_stage_dp_delay_regg_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_9_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_9_port, QN => 
                           n_1457);
   datapath_i_memory_stage_dp_delay_regg_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_8_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_8_port, QN => 
                           n_1458);
   datapath_i_memory_stage_dp_delay_regg_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_7_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_7_port, QN => 
                           n_1459);
   datapath_i_memory_stage_dp_delay_regg_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_6_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_6_port, QN => 
                           n_1460);
   datapath_i_memory_stage_dp_delay_regg_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_5_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_5_port, QN => 
                           n_1461);
   datapath_i_memory_stage_dp_delay_regg_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_4_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_4_port, QN => 
                           n_1462);
   datapath_i_memory_stage_dp_delay_regg_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_3_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_3_port, QN => 
                           n_1463);
   datapath_i_memory_stage_dp_delay_regg_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_2_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_2_port, QN => 
                           n_1464);
   datapath_i_memory_stage_dp_delay_regg_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_1_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_1_port, QN => 
                           n_1465);
   datapath_i_memory_stage_dp_delay_regg_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_0_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_0_port, QN => 
                           n_1466);
   datapath_i_memory_stage_dp_lmd_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_31_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_31_port, QN => n_1467)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_30_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_30_port, QN => n_1468)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_29_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_29_port, QN => n_1469)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_28_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_28_port, QN => n_1470)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_27_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_27_port, QN => n_1471)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_26_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_26_port, QN => n_1472)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_25_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_25_port, QN => n_1473)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_24_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_24_port, QN => n_1474)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_23_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_23_port, QN => n_1475)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_22_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_22_port, QN => n_1476)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_21_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_21_port, QN => n_1477)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_20_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_20_port, QN => n_1478)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_19_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_19_port, QN => n_1479)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_18_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_18_port, QN => n_1480)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_17_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_17_port, QN => n_1481)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_16_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_16_port, QN => n_1482)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_15_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_15_port, QN => n_1483)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_14_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_14_port, QN => n_1484)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_13_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_13_port, QN => n_1485)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_12_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_12_port, QN => n_1486)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_11_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_11_port, QN => n_1487)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_10_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_10_port, QN => n_1488)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_9_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_9_port, QN => n_1489);
   datapath_i_memory_stage_dp_lmd_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_8_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_8_port, QN => n_1490);
   datapath_i_memory_stage_dp_lmd_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_7_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_7_port, QN => n_1491);
   datapath_i_memory_stage_dp_lmd_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_6_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_6_port, QN => n_1492);
   datapath_i_memory_stage_dp_lmd_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_5_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_5_port, QN => n_1493);
   datapath_i_memory_stage_dp_lmd_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_4_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_4_port, QN => n_1494);
   datapath_i_memory_stage_dp_lmd_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_3_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_3_port, QN => n_1495);
   datapath_i_memory_stage_dp_lmd_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_2_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_2_port, QN => n_1496);
   datapath_i_memory_stage_dp_lmd_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_1_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_1_port, QN => n_1497);
   datapath_i_memory_stage_dp_lmd_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_0_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_0_port, QN => n_1498);
   datapath_i_execute_stage_dp_reg_del_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_31_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_31_port, QN => n_1499);
   datapath_i_execute_stage_dp_reg_del_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_30_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_30_port, QN => n_1500);
   datapath_i_execute_stage_dp_reg_del_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_29_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_29_port, QN => n_1501);
   datapath_i_execute_stage_dp_reg_del_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_28_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_28_port, QN => n_1502);
   datapath_i_execute_stage_dp_reg_del_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_27_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_27_port, QN => n_1503);
   datapath_i_execute_stage_dp_reg_del_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_26_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_26_port, QN => n_1504);
   datapath_i_execute_stage_dp_reg_del_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_25_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_25_port, QN => n_1505);
   datapath_i_execute_stage_dp_reg_del_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_24_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_24_port, QN => n_1506);
   datapath_i_execute_stage_dp_reg_del_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_23_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_23_port, QN => n_1507);
   datapath_i_execute_stage_dp_reg_del_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_22_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_22_port, QN => n_1508);
   datapath_i_execute_stage_dp_reg_del_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_21_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_21_port, QN => n_1509);
   datapath_i_execute_stage_dp_reg_del_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_20_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_20_port, QN => n_1510);
   datapath_i_execute_stage_dp_reg_del_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_19_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_19_port, QN => n_1511);
   datapath_i_execute_stage_dp_reg_del_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_18_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_18_port, QN => n_1512);
   datapath_i_execute_stage_dp_reg_del_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_17_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_17_port, QN => n_1513);
   datapath_i_execute_stage_dp_reg_del_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_16_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_16_port, QN => n_1514);
   datapath_i_execute_stage_dp_reg_del_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_15_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_15_port, QN => n_1515);
   datapath_i_execute_stage_dp_reg_del_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_14_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_14_port, QN => n_1516);
   datapath_i_execute_stage_dp_reg_del_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_13_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_13_port, QN => n_1517);
   datapath_i_execute_stage_dp_reg_del_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_12_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_12_port, QN => n_1518);
   datapath_i_execute_stage_dp_reg_del_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_11_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_11_port, QN => n_1519);
   datapath_i_execute_stage_dp_reg_del_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_10_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_10_port, QN => n_1520);
   datapath_i_execute_stage_dp_reg_del_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_9_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_9_port, QN => n_1521);
   datapath_i_execute_stage_dp_reg_del_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_8_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_8_port, QN => n_1522);
   datapath_i_execute_stage_dp_reg_del_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_7_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_7_port, QN => n_1523);
   datapath_i_execute_stage_dp_reg_del_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_6_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_6_port, QN => n_1524);
   datapath_i_execute_stage_dp_reg_del_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_5_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_5_port, QN => n_1525);
   datapath_i_execute_stage_dp_reg_del_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_4_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_4_port, QN => n_1526);
   datapath_i_execute_stage_dp_reg_del_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_3_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_3_port, QN => n_1527);
   datapath_i_execute_stage_dp_reg_del_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_2_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_2_port, QN => n_1528);
   datapath_i_execute_stage_dp_reg_del_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_1_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_1_port, QN => n_1529);
   datapath_i_execute_stage_dp_reg_del_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_0_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_0_port, QN => n_1530);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_31_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_31_port, QN => n_1531);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_30_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_30_port, QN => n_1532);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_29_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_29_port, QN => n_1533);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_28_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_28_port, QN => n_1534);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_27_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_27_port, QN => n_1535);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_26_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_26_port, QN => n_1536);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_25_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_25_port, QN => n_1537);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_24_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_24_port, QN => n_1538);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_23_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_23_port, QN => n_1539);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_22_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_22_port, QN => n_1540);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_21_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_21_port, QN => n_1541);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_20_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_20_port, QN => n_1542);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_19_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_19_port, QN => n_1543);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_18_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_18_port, QN => n_1544);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_17_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_17_port, QN => n_1545);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_16_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_16_port, QN => n_1546);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_15_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_15_port, QN => n_1547);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_14_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_14_port, QN => n_1548);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_13_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_13_port, QN => n_1549);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_12_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_12_port, QN => n_1550);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_11_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_11_port, QN => n_1551);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_10_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_10_port, QN => n_1552);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_9_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_9_port, QN => n_1553);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_8_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_8_port, QN => n_1554);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_7_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_7_port, QN => n_1555);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_6_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_6_port, QN => n_1556);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_5_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_5_port, QN => n_1557);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_4_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_4_port, QN => n_1558);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_3_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_3_port, QN => n_1559);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_2_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_2_port, QN => n_1560);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_1_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_1_port, QN => n_1561);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_0_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_0_port, QN => n_1562);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_32_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_32_port, CK 
                           => CLK, RN => RST, Q => n_1563, QN => n703);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_31_port, CK 
                           => CLK, RN => RST, Q => n_1564, QN => n727);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_30_port, CK 
                           => CLK, RN => RST, Q => n_1565, QN => n726);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_29_port, CK 
                           => CLK, RN => RST, Q => n_1566, QN => n725);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_28_port, CK 
                           => CLK, RN => RST, Q => n_1567, QN => n724);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_27_port, CK 
                           => CLK, RN => RST, Q => n_1568, QN => n691);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_26_port, CK 
                           => CLK, RN => RST, Q => n_1569, QN => n723);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_25_port, CK 
                           => CLK, RN => RST, Q => n_1570, QN => n722);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_24_port, CK 
                           => CLK, RN => RST, Q => n_1571, QN => n721);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_23_port, CK 
                           => CLK, RN => RST, Q => n_1572, QN => n720);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_22_port, CK 
                           => CLK, RN => RST, Q => n_1573, QN => n719);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_21_port, CK 
                           => CLK, RN => RST, Q => n_1574, QN => n718);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_20_port, CK 
                           => CLK, RN => RST, Q => n_1575, QN => n717);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_19_port, CK 
                           => CLK, RN => RST, Q => n_1576, QN => n716);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_18_port, CK 
                           => CLK, RN => RST, Q => n_1577, QN => n715);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_17_port, CK 
                           => CLK, RN => RST, Q => n_1578, QN => n714);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_16_port, CK 
                           => CLK, RN => RST, Q => n_1579, QN => n713);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_15_port, CK 
                           => CLK, RN => RST, Q => n_1580, QN => n712);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_14_port, CK 
                           => CLK, RN => RST, Q => n_1581, QN => n711);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_13_port, CK 
                           => CLK, RN => RST, Q => n_1582, QN => n710);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_12_port, CK 
                           => CLK, RN => RST, Q => n_1583, QN => n709);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_11_port, CK 
                           => CLK, RN => RST, Q => n_1584, QN => n708);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_10_port, CK 
                           => CLK, RN => RST, Q => n_1585, QN => n707);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_9_port, CK 
                           => CLK, RN => RST, Q => n_1586, QN => n706);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_8_port, CK 
                           => CLK, RN => RST, Q => n_1587, QN => n705);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_7_port, CK 
                           => CLK, RN => RST, Q => n_1588, QN => n732);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_6_port, CK 
                           => CLK, RN => RST, Q => n_1589, QN => n731);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_5_port, CK 
                           => CLK, RN => RST, Q => n_1590, QN => n730);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_4_port, CK 
                           => CLK, RN => RST, Q => n_1591, QN => n729);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_3_port, CK 
                           => CLK, RN => RST, Q => n_1592, QN => n728);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_2_port, CK 
                           => CLK, RN => RST, Q => n_1593, QN => n734);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_1_port, CK 
                           => CLK, RN => RST, Q => n_1594, QN => n733);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_31_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_32_port, QN => 
                           n_1595);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_30_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_31_port, QN => 
                           n_1596);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_29_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_30_port, QN => 
                           n_1597);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_28_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_29_port, QN => 
                           n_1598);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_27_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_28_port, QN => 
                           n_1599);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_26_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_27_port, QN => 
                           n_1600);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_25_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_26_port, QN => 
                           n_1601);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_24_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_25_port, QN => 
                           n_1602);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_23_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_24_port, QN => 
                           n_1603);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_22_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_23_port, QN => 
                           n_1604);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_21_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_22_port, QN => 
                           n_1605);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_20_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_21_port, QN => 
                           n_1606);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_19_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_20_port, QN => 
                           n_1607);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_18_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_19_port, QN => 
                           n_1608);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_17_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_18_port, QN => 
                           n_1609);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_16_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_17_port, QN => 
                           n_1610);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_15_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_16_port, QN => 
                           n_1611);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_14_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_15_port, QN => 
                           n_1612);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_13_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_14_port, QN => 
                           n_1613);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_12_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_13_port, QN => 
                           n_1614);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_11_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_12_port, QN => 
                           n_1615);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_10_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_11_port, QN => 
                           n_1616);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_9_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_10_port, QN => 
                           n_1617);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_8_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_9_port, QN => 
                           n_1618);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_7_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_8_port, QN => 
                           n_1619);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_6_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_7_port, QN => 
                           n_1620);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_5_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_6_port, QN => 
                           n_1621);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_4_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_5_port, QN => 
                           n_1622);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_3_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_4_port, QN => 
                           n_1623);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_2_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_3_port, QN => 
                           n_1624);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_1_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_2_port, QN => 
                           n_1625);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_0_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_1_port, QN => 
                           n_1626);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n4674, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_0_port, QN => 
                           n_1627);
   datapath_i_decode_stage_dp_reg_immediate_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_25_port, QN 
                           => n_1628);
   datapath_i_decode_stage_dp_reg_immediate_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_24_port, QN 
                           => n_1629);
   datapath_i_decode_stage_dp_reg_immediate_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_23_port, QN 
                           => n_1630);
   datapath_i_decode_stage_dp_reg_immediate_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_22_port, QN 
                           => n_1631);
   datapath_i_decode_stage_dp_reg_immediate_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_21_port, QN 
                           => n_1632);
   datapath_i_decode_stage_dp_reg_immediate_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_20_port, QN 
                           => n_1633);
   datapath_i_decode_stage_dp_reg_immediate_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_19_port, QN 
                           => n_1634);
   datapath_i_decode_stage_dp_reg_immediate_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_18_port, QN 
                           => n_1635);
   datapath_i_decode_stage_dp_reg_immediate_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_17_port, QN 
                           => n_1636);
   datapath_i_decode_stage_dp_reg_immediate_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_16_port, QN 
                           => n_1637);
   datapath_i_decode_stage_dp_reg_immediate_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_15_port, QN 
                           => n_1638);
   datapath_i_decode_stage_dp_reg_immediate_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_14_port, QN 
                           => n_1639);
   datapath_i_decode_stage_dp_reg_immediate_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_13_port, QN 
                           => n_1640);
   datapath_i_decode_stage_dp_reg_immediate_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_12_port, QN 
                           => n_1641);
   datapath_i_decode_stage_dp_reg_immediate_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_11_port, QN 
                           => n_1642);
   datapath_i_decode_stage_dp_reg_immediate_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_10_port, QN 
                           => n_1643);
   datapath_i_decode_stage_dp_reg_immediate_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_9_port, QN 
                           => n_1644);
   datapath_i_decode_stage_dp_reg_immediate_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_8_port, QN 
                           => n_1645);
   datapath_i_decode_stage_dp_reg_immediate_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_7_port, QN 
                           => n_1646);
   datapath_i_decode_stage_dp_reg_immediate_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_6_port, QN 
                           => n_1647);
   datapath_i_decode_stage_dp_reg_immediate_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_5_port, QN 
                           => n_1648);
   datapath_i_decode_stage_dp_reg_immediate_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_4_port, QN 
                           => n_1649);
   datapath_i_decode_stage_dp_reg_immediate_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_3_port, QN 
                           => n_1650);
   datapath_i_decode_stage_dp_reg_immediate_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_2_port, QN 
                           => n_1651);
   datapath_i_decode_stage_dp_reg_immediate_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_1_port, QN 
                           => n_1652);
   datapath_i_decode_stage_dp_reg_immediate_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_0_port, QN 
                           => n_1653);
   datapath_i_decode_stage_dp_reg_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_31_port, 
                           QN => n764);
   datapath_i_decode_stage_dp_reg_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_30_port, 
                           QN => n763);
   datapath_i_decode_stage_dp_reg_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_29_port, 
                           QN => n762);
   datapath_i_decode_stage_dp_reg_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_28_port, 
                           QN => n761);
   datapath_i_decode_stage_dp_reg_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_27_port, 
                           QN => n760);
   datapath_i_decode_stage_dp_reg_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_26_port, 
                           QN => n759);
   datapath_i_decode_stage_dp_reg_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_25_port, 
                           QN => n758);
   datapath_i_decode_stage_dp_reg_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_24_port, 
                           QN => n_1654);
   datapath_i_decode_stage_dp_reg_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_23_port, 
                           QN => n_1655);
   datapath_i_decode_stage_dp_reg_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_22_port, 
                           QN => n_1656);
   datapath_i_decode_stage_dp_reg_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_21_port, 
                           QN => n_1657);
   datapath_i_decode_stage_dp_reg_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_20_port, 
                           QN => n_1658);
   datapath_i_decode_stage_dp_reg_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_19_port, 
                           QN => n_1659);
   datapath_i_decode_stage_dp_reg_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_18_port, 
                           QN => n_1660);
   datapath_i_decode_stage_dp_reg_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_17_port, 
                           QN => n_1661);
   datapath_i_decode_stage_dp_reg_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_16_port, 
                           QN => n_1662);
   datapath_i_decode_stage_dp_reg_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_15_port, 
                           QN => n_1663);
   datapath_i_decode_stage_dp_reg_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_14_port, 
                           QN => n_1664);
   datapath_i_decode_stage_dp_reg_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_13_port, 
                           QN => n_1665);
   datapath_i_decode_stage_dp_reg_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_12_port, 
                           QN => n_1666);
   datapath_i_decode_stage_dp_reg_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_11_port, 
                           QN => n_1667);
   datapath_i_decode_stage_dp_reg_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_10_port, 
                           QN => n_1668);
   datapath_i_decode_stage_dp_reg_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_9_port, QN 
                           => n_1669);
   datapath_i_decode_stage_dp_reg_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_8_port, QN 
                           => n_1670);
   datapath_i_decode_stage_dp_reg_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_7_port, QN 
                           => n_1671);
   datapath_i_decode_stage_dp_reg_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_6_port, QN 
                           => n_1672);
   datapath_i_decode_stage_dp_reg_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_5_port, QN 
                           => n_1673);
   datapath_i_decode_stage_dp_reg_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_4_port, QN 
                           => n_1674);
   datapath_i_decode_stage_dp_reg_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_3_port, QN 
                           => n_1675);
   datapath_i_decode_stage_dp_reg_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_2_port, QN 
                           => n_1676);
   datapath_i_decode_stage_dp_reg_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_1_port, QN 
                           => n_1677);
   datapath_i_decode_stage_dp_reg_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_0_port, QN 
                           => n_1678);
   datapath_i_decode_stage_dp_reg_a_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_31_port, 
                           QN => n_1679);
   datapath_i_decode_stage_dp_reg_a_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_30_port, 
                           QN => n_1680);
   datapath_i_decode_stage_dp_reg_a_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_29_port, 
                           QN => n_1681);
   datapath_i_decode_stage_dp_reg_a_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_28_port, 
                           QN => n_1682);
   datapath_i_decode_stage_dp_reg_a_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_27_port, 
                           QN => n_1683);
   datapath_i_decode_stage_dp_reg_a_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_26_port, 
                           QN => n_1684);
   datapath_i_decode_stage_dp_reg_a_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_25_port, 
                           QN => n_1685);
   datapath_i_decode_stage_dp_reg_a_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_24_port, 
                           QN => n_1686);
   datapath_i_decode_stage_dp_reg_a_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_23_port, 
                           QN => n_1687);
   datapath_i_decode_stage_dp_reg_a_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_22_port, 
                           QN => n_1688);
   datapath_i_decode_stage_dp_reg_a_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_21_port, 
                           QN => n_1689);
   datapath_i_decode_stage_dp_reg_a_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_20_port, 
                           QN => n_1690);
   datapath_i_decode_stage_dp_reg_a_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_19_port, 
                           QN => n_1691);
   datapath_i_decode_stage_dp_reg_a_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_18_port, 
                           QN => n_1692);
   datapath_i_decode_stage_dp_reg_a_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_17_port, 
                           QN => n_1693);
   datapath_i_decode_stage_dp_reg_a_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_16_port, 
                           QN => n_1694);
   datapath_i_decode_stage_dp_reg_a_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_15_port, 
                           QN => n_1695);
   datapath_i_decode_stage_dp_reg_a_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_14_port, 
                           QN => n_1696);
   datapath_i_decode_stage_dp_reg_a_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_13_port, 
                           QN => n_1697);
   datapath_i_decode_stage_dp_reg_a_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_12_port, 
                           QN => n_1698);
   datapath_i_decode_stage_dp_reg_a_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_11_port, 
                           QN => n_1699);
   datapath_i_decode_stage_dp_reg_a_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_10_port, 
                           QN => n_1700);
   datapath_i_decode_stage_dp_reg_a_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_9_port, QN 
                           => n_1701);
   datapath_i_decode_stage_dp_reg_a_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_8_port, QN 
                           => n_1702);
   datapath_i_decode_stage_dp_reg_a_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_7_port, QN 
                           => n_1703);
   datapath_i_decode_stage_dp_reg_a_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_6_port, QN 
                           => n_1704);
   datapath_i_decode_stage_dp_reg_a_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_5_port, QN 
                           => n_1705);
   datapath_i_decode_stage_dp_reg_a_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_4_port, QN 
                           => n_1706);
   datapath_i_decode_stage_dp_reg_a_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_3_port, QN 
                           => n_1707);
   datapath_i_decode_stage_dp_reg_a_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_2_port, QN 
                           => n_1708);
   datapath_i_decode_stage_dp_reg_a_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_1_port, QN 
                           => n_1709);
   datapath_i_decode_stage_dp_reg_a_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_0_port, QN 
                           => n_1710);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           QN => n_1711);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           QN => n_1712);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           QN => n_1713);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           QN => n_1714);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           QN => n_1715);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_4_port, QN 
                           => n_1716);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_3_port, QN 
                           => n_1717);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_2_port, QN 
                           => n_1718);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_1_port, QN 
                           => n_1719);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_0_port, QN 
                           => n_1720);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => n4279, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_4_port, QN 
                           => n_1721);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => n4278, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_3_port, QN 
                           => n_1722);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n78, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_2_port, QN 
                           => n_1723);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => n4277, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_1_port, QN 
                           => n_1724);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n4276, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_0_port, QN 
                           => n_1725);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n69, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_31_port, QN => 
                           n4669);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n68, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_30_port, QN => 
                           n_1726);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n67, CK => CLK, RN => 
                           RST, Q => n4655, QN => n737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n66, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_28_port, QN => 
                           n4664);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n65, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_27_port, QN => 
                           n4658);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n64, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_26_port, QN => 
                           n4656);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n63, CK => CLK, RN => 
                           RST, Q => datapath_i_n9, QN => n_1727);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n62, CK => CLK, RN => 
                           RST, Q => datapath_i_n10, QN => n_1728);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n61, CK => CLK, RN => 
                           RST, Q => datapath_i_n11, QN => n_1729);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n60, CK => CLK, RN => 
                           RST, Q => datapath_i_n12, QN => n_1730);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n59, CK => CLK, RN => 
                           RST, Q => datapath_i_n13, QN => n_1731);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n58, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_20_port, QN => 
                           n_1732);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n57, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_19_port, QN => 
                           n_1733);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n56, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_18_port, QN => 
                           n697);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n55, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_17_port, QN => 
                           n_1734);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n54, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_16_port, QN => 
                           n_1735);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n53, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_15_port, QN => 
                           n_1736);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n52, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_14_port, QN => 
                           n_1737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n51, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_13_port, QN => 
                           n740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n50, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_12_port, QN => 
                           n_1738);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n49, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_11_port, QN => 
                           n_1739);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n48, CK => CLK, RN => 
                           RST, Q => datapath_i_n14, QN => n_1740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n47, CK => CLK, RN => 
                           RST, Q => datapath_i_n15, QN => n_1741);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n46, CK => CLK, RN => 
                           RST, Q => datapath_i_n16, QN => n_1742);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n45, CK => CLK, RN => 
                           RST, Q => datapath_i_n17, QN => n_1743);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n44, CK => CLK, RN => 
                           RST, Q => datapath_i_n18, QN => n_1744);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n43, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_5_port, QN => 
                           n4672);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n42, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_4_port, QN => 
                           n4670);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n41, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_3_port, QN => 
                           n4660);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n40, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_2_port, QN => 
                           n4661);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n39, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_1_port, QN => 
                           n_1745);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n38, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_0_port, QN => 
                           n4666);
   datapath_i_fetch_stage_dp_new_program_counter_D_I_31_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n2, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_31_port, QN => n_1746
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_30_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n3, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_30_port, QN => n_1747
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_29_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n4, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_29_port, QN => n_1748
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_28_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n9, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_28_port, QN => n_1749
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_27_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n10, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_27_port, QN => n_1750
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_26_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n11, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_26_port, QN => n_1751
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_25_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n12, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_25_port, QN => n_1752
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_24_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n13, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_24_port, QN => n_1753
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_23_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n14, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_23_port, QN => n_1754
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_22_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n15, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_22_port, QN => n_1755
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_21_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n16, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_21_port, QN => n_1756
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_20_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n17, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_20_port, QN => n_1757
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_19_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n18, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_19_port, QN => n_1758
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_18_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n19, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_18_port, QN => n_1759
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_17_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n20, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_17_port, QN => n_1760
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_16_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n21, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_16_port, QN => n_1761
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_15_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n22, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_15_port, QN => n_1762
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_14_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n23, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_14_port, QN => n_1763
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_13_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n24, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_13_port, QN => n_1764
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_12_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n25, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_12_port, QN => n_1765
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_11_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n26, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_11_port, QN => n_1766
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_10_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n27, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_10_port, QN => n_1767
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_9_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n28, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_9_port, QN => n_1768)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_8_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n29, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_8_port, QN => n_1769)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_7_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n30, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_7_port, QN => n_1770)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_6_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n31, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_6_port, QN => n_1771)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_5_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n32, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_5_port, QN => n_1772)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_4_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n33, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_4_port, QN => n_1773)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_3_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n34, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_3_port, QN => n_1774)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_2_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n35, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_2_port, QN => n_1775)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_1_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n36, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_1_port, QN => n_1776)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n37, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_0_port, QN => n_1777)
                           ;
   datapath_i_fetch_stage_dp_program_counter_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_31_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_31_port, QN => 
                           n_1778);
   datapath_i_fetch_stage_dp_program_counter_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_30_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_30_port, QN => 
                           n_1779);
   datapath_i_fetch_stage_dp_program_counter_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_29_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_29_port, QN => 
                           n753);
   datapath_i_fetch_stage_dp_program_counter_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_28_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_28_port, QN => 
                           n_1780);
   datapath_i_fetch_stage_dp_program_counter_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_27_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_27_port, QN => 
                           n751);
   datapath_i_fetch_stage_dp_program_counter_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_26_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_26_port, QN => 
                           n_1781);
   datapath_i_fetch_stage_dp_program_counter_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_25_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_25_port, QN => 
                           n750);
   datapath_i_fetch_stage_dp_program_counter_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_24_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_24_port, QN => 
                           n_1782);
   datapath_i_fetch_stage_dp_program_counter_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_23_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_23_port, QN => 
                           n749);
   datapath_i_fetch_stage_dp_program_counter_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_22_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_22_port, QN => 
                           n_1783);
   datapath_i_fetch_stage_dp_program_counter_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_21_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_21_port, QN => 
                           n748);
   datapath_i_fetch_stage_dp_program_counter_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_20_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_20_port, QN => 
                           n_1784);
   datapath_i_fetch_stage_dp_program_counter_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_19_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_19_port, QN => 
                           n747);
   datapath_i_fetch_stage_dp_program_counter_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_18_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_18_port, QN => 
                           n_1785);
   datapath_i_fetch_stage_dp_program_counter_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_17_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_17_port, QN => 
                           n746);
   datapath_i_fetch_stage_dp_program_counter_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_16_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_16_port, QN => 
                           n_1786);
   datapath_i_fetch_stage_dp_program_counter_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_15_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_15_port, QN => 
                           n745);
   datapath_i_fetch_stage_dp_program_counter_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_14_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_14_port, QN => 
                           n_1787);
   datapath_i_fetch_stage_dp_program_counter_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_13_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_13_port, QN => 
                           n752);
   datapath_i_fetch_stage_dp_program_counter_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_12_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_12_port, QN => 
                           n_1788);
   datapath_i_fetch_stage_dp_program_counter_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_11_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_11_port, QN => 
                           n744);
   datapath_i_fetch_stage_dp_program_counter_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_10_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_10_port, QN => 
                           n_1789);
   datapath_i_fetch_stage_dp_program_counter_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_9_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_9_port, QN => n743
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_8_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_8_port, QN => 
                           n_1790);
   datapath_i_fetch_stage_dp_program_counter_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_7_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_7_port, QN => n742
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_6_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_6_port, QN => 
                           n_1791);
   datapath_i_fetch_stage_dp_program_counter_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_5_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_5_port, QN => n741
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_4_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_1792);
   datapath_i_fetch_stage_dp_program_counter_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_3_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_1793);
   datapath_i_fetch_stage_dp_program_counter_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_2_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_2_port, QN => 
                           n_1794);
   datapath_i_fetch_stage_dp_program_counter_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N6, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N40_port, QN => 
                           n_1795);
   datapath_i_fetch_stage_dp_program_counter_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N5, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N39_port, QN => 
                           n_1796);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   datapath_i_execute_stage_dp_condition_delay_reg_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
                           CK => CLK, RN => RST, Q => n4657, QN => n4662);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_0_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, QN => 
                           n_1797);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_counter_mul_reg_1_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_1_port, CK => CLK, RN => 
                           RST, Q => n4665, QN => cu_i_n26);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_counter_mul_reg_2_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_2_port, CK => CLK, RN => 
                           RST, Q => n4671, QN => cu_i_n25);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_counter_mul_reg_3_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_3_port, CK => CLK, RN => 
                           RST, Q => n4667, QN => cu_i_n124);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_next_val_counter_mul_1_port);
   cu_i_counter_mul_reg_0_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_0_port, CK => CLK, RN => 
                           RST, Q => n4659, QN => cu_i_n125);
   U3963 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(0), ZN => 
                           datapath_i_memory_stage_dp_data_ir_0_port);
   U3964 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(10), ZN => 
                           datapath_i_memory_stage_dp_data_ir_10_port);
   U3965 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(11), ZN => 
                           datapath_i_memory_stage_dp_data_ir_11_port);
   U3966 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(12), ZN => 
                           datapath_i_memory_stage_dp_data_ir_12_port);
   U3967 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(13), ZN => 
                           datapath_i_memory_stage_dp_data_ir_13_port);
   U3968 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(14), ZN => 
                           datapath_i_memory_stage_dp_data_ir_14_port);
   U3969 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(15), ZN => 
                           datapath_i_memory_stage_dp_data_ir_15_port);
   U3970 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(16), ZN => 
                           datapath_i_memory_stage_dp_data_ir_16_port);
   U3971 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(17), ZN => 
                           datapath_i_memory_stage_dp_data_ir_17_port);
   U3972 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(18), ZN => 
                           datapath_i_memory_stage_dp_data_ir_18_port);
   U3973 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(19), ZN => 
                           datapath_i_memory_stage_dp_data_ir_19_port);
   U3974 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(1), ZN => 
                           datapath_i_memory_stage_dp_data_ir_1_port);
   U3975 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(20), ZN => 
                           datapath_i_memory_stage_dp_data_ir_20_port);
   U3976 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(21), ZN => 
                           datapath_i_memory_stage_dp_data_ir_21_port);
   U3977 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(22), ZN => 
                           datapath_i_memory_stage_dp_data_ir_22_port);
   U3978 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(23), ZN => 
                           datapath_i_memory_stage_dp_data_ir_23_port);
   U3979 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(24), ZN => 
                           datapath_i_memory_stage_dp_data_ir_24_port);
   U3980 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(25), ZN => 
                           datapath_i_memory_stage_dp_data_ir_25_port);
   U3981 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(26), ZN => 
                           datapath_i_memory_stage_dp_data_ir_26_port);
   U3982 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(27), ZN => 
                           datapath_i_memory_stage_dp_data_ir_27_port);
   U3983 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(28), ZN => 
                           datapath_i_memory_stage_dp_data_ir_28_port);
   U3984 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(29), ZN => 
                           datapath_i_memory_stage_dp_data_ir_29_port);
   U3985 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(2), ZN => 
                           datapath_i_memory_stage_dp_data_ir_2_port);
   U3986 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(30), ZN => 
                           datapath_i_memory_stage_dp_data_ir_30_port);
   U3987 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(31), ZN => 
                           datapath_i_memory_stage_dp_data_ir_31_port);
   U3988 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(3), ZN => 
                           datapath_i_memory_stage_dp_data_ir_3_port);
   U3989 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(4), ZN => 
                           datapath_i_memory_stage_dp_data_ir_4_port);
   U3990 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(5), ZN => 
                           datapath_i_memory_stage_dp_data_ir_5_port);
   U3991 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(6), ZN => 
                           datapath_i_memory_stage_dp_data_ir_6_port);
   U3992 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(7), ZN => 
                           datapath_i_memory_stage_dp_data_ir_7_port);
   U3993 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(8), ZN => 
                           datapath_i_memory_stage_dp_data_ir_8_port);
   U3994 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(9), ZN => 
                           datapath_i_memory_stage_dp_data_ir_9_port);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_next_val_counter_mul_2_port);
   cu_i_curr_state_reg_1_inst : DFFR_X1 port map( D => cu_i_n209, CK => CLK, RN
                           => RST, Q => n_1798, QN => cu_i_n123);
   cu_i_curr_state_reg_0_inst : DFFS_X1 port map( D => cu_i_n210, CK => CLK, SN
                           => RST, Q => n4668, QN => cu_i_n23);
   cu_i_stall_reg : DFFR_X2 port map( D => cu_i_next_stall, CK => CLK, RN => 
                           RST, Q => n704, QN => n4663);
   U3995 : NAND2_X1 port map( A1 => n4283, A2 => n4667, ZN => n4413);
   U3996 : NOR4_X1 port map( A1 => n4395, A2 => n4670, A3 => n4410, A4 => n4660
                           , ZN => n4374);
   U3997 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           n4669, A3 => n4656, A4 => n4418, ZN => 
                           cu_i_cmd_word_4_port);
   U3998 : AOI21_X1 port map( B1 => n4545, B2 => n4544, A => cu_i_cw3_6_port, 
                           ZN => n4546);
   U3999 : AND2_X1 port map( A1 => n4568, A2 => n4546, ZN => n4583);
   U4000 : OAI21_X1 port map( B1 => n4413, B2 => n4414, A => n699, ZN => 
                           write_rf_i);
   U4001 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_0_port, B1
                           => cu_i_cw1_0_port, B2 => n4663, ZN => n4377);
   U4002 : NAND2_X1 port map( A1 => cu_i_n25, A2 => cu_i_n26, ZN => n4283);
   U4003 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U4004 : NOR2_X1 port map( A1 => n4377, A2 => n4364, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U4005 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           curr_instruction_to_cu_i_27_port, A3 => 
                           curr_instruction_to_cu_i_30_port, A4 => n4362, ZN =>
                           n4426);
   U4006 : NOR2_X1 port map( A1 => cu_i_n123, A2 => n4668, ZN => n4363);
   U4007 : CLKBUF_X1 port map( A => n4654, Z => n4643);
   U4008 : CLKBUF_X1 port map( A => n4533, Z => n4348);
   U4009 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n4662, ZN => n4533);
   U4010 : CLKBUF_X1 port map( A => n4490, Z => n4539);
   U4011 : AOI21_X1 port map( B1 => n4292, B2 => n4374, A => n4390, ZN => n4542
                           );
   U4012 : INV_X1 port map( A => n704, ZN => n4436);
   U4013 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n4363, A3 => n4664, ZN => n4418);
   U4014 : OAI22_X1 port map( A1 => n4663, A2 => cu_i_cmd_word_4_port, B1 => 
                           cu_i_cw2_8_port, B2 => n704, ZN => n309);
   U4015 : INV_X1 port map( A => n309, ZN => DRAM_ENABLE_port);
   U4016 : INV_X1 port map( A => cu_i_cmd_word_4_port, ZN => n4540);
   U4017 : NOR2_X1 port map( A1 => n4655, A2 => n4540, ZN => 
                           cu_i_cmd_word_3_port);
   U4018 : OAI22_X1 port map( A1 => n4663, A2 => cu_i_cmd_word_3_port, B1 => 
                           cu_i_cw2_7_port, B2 => n704, ZN => n4375);
   U4019 : NAND2_X1 port map( A1 => DRAM_ENABLE_port, A2 => n4375, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U4020 : CLKBUF_X1 port map( A => datapath_i_memory_stage_dp_n2, Z => n4679);
   U4021 : INV_X1 port map( A => DRAM_ENABLE_port, ZN => n4677);
   U4022 : NAND4_X1 port map( A1 => cu_i_n26, A2 => cu_i_n25, A3 => n4659, A4 
                           => n4667, ZN => cu_i_n145);
   U4023 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           curr_instruction_to_cu_i_31_port, ZN => n4360);
   U4024 : NAND3_X1 port map( A1 => n4363, A2 => n737, A3 => n4360, ZN => n4291
                           );
   U4025 : OR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n4658
                           , A3 => n4291, ZN => n4586);
   U4026 : INV_X1 port map( A => n4586, ZN => n4674);
   U4027 : NAND2_X1 port map( A1 => cu_i_n145, A2 => n4413, ZN => n4292);
   U4028 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_1_port, A2 => 
                           curr_instruction_to_cu_i_5_port, ZN => n4395);
   U4029 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => 
                           curr_instruction_to_cu_i_0_port, ZN => n4410);
   U4030 : NOR3_X1 port map( A1 => n4655, A2 => 
                           curr_instruction_to_cu_i_31_port, A3 => 
                           curr_instruction_to_cu_i_26_port, ZN => n4359);
   U4031 : INV_X1 port map( A => n4359, ZN => n4362);
   U4032 : NAND2_X1 port map( A1 => n4363, A2 => n4426, ZN => n4390);
   U4033 : INV_X1 port map( A => n4542, ZN => n4541);
   U4034 : AOI221_X1 port map( B1 => n4541, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n4542, C2 =>
                           curr_instruction_to_cu_i_11_port, A => n4674, ZN => 
                           n4284);
   U4035 : INV_X1 port map( A => n4284, ZN => n4276);
   U4036 : AOI221_X1 port map( B1 => n4541, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n4542, C2 =>
                           curr_instruction_to_cu_i_12_port, A => n4674, ZN => 
                           n4285);
   U4037 : INV_X1 port map( A => n4285, ZN => n4277);
   U4038 : AOI221_X1 port map( B1 => n4541, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n4542, C2 =>
                           curr_instruction_to_cu_i_14_port, A => n4674, ZN => 
                           n4286);
   U4039 : INV_X1 port map( A => n4286, ZN => n4278);
   U4040 : INV_X1 port map( A => n4662, ZN => n4531);
   U4041 : NOR2_X1 port map( A1 => n4657, A2 => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, ZN => 
                           n4530);
   U4042 : CLKBUF_X1 port map( A => n4530, Z => n4524);
   U4043 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_2_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_2_port, ZN => 
                           n4287);
   U4044 : OAI21_X1 port map( B1 => n728, B2 => n4348, A => n4287, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U4045 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_3_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_3_port, ZN => 
                           n4288);
   U4046 : OAI21_X1 port map( B1 => n729, B2 => n4348, A => n4288, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U4047 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_5_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_5_port, ZN => 
                           n4289);
   U4048 : OAI21_X1 port map( B1 => n731, B2 => n4533, A => n4289, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_5_port);
   U4049 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_4_port, ZN => 
                           n4290);
   U4050 : OAI21_X1 port map( B1 => n730, B2 => n4348, A => n4290, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U4051 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n4658, ZN => n4368);
   U4052 : OR2_X1 port map( A1 => n4291, A2 => n4368, ZN => n4587);
   U4053 : NAND2_X1 port map( A1 => n4586, A2 => n4587, ZN => n1152);
   U4054 : NAND2_X1 port map( A1 => n4374, A2 => n4426, ZN => n4367);
   U4055 : OAI21_X1 port map( B1 => n4292, B2 => n4367, A => n4363, ZN => n4293
                           );
   U4056 : NAND2_X1 port map( A1 => cu_i_n123, A2 => n4668, ZN => n4430);
   U4057 : AOI21_X1 port map( B1 => n4293, B2 => n4430, A => n704, ZN => 
                           IRAM_ENABLE_port);
   U4058 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_5_port, ZN
                           => n4294);
   U4059 : NAND3_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port,
                           A2 => datapath_i_new_pc_value_mem_stage_i_2_port, A3
                           => datapath_i_new_pc_value_mem_stage_i_3_port, ZN =>
                           n4445);
   U4060 : INV_X1 port map( A => n1152, ZN => n4431);
   U4061 : OAI221_X1 port map( B1 => n4663, B2 => n4431, C1 => n704, C2 => n756
                           , A => n4662, ZN => n4442);
   U4062 : INV_X1 port map( A => n4442, ZN => n4490);
   U4063 : NOR2_X1 port map( A1 => n4294, A2 => n4445, ZN => n4452);
   U4064 : AOI211_X1 port map( C1 => n4294, C2 => n4445, A => n4490, B => n4452
                           , ZN => n4296);
   U4065 : NAND2_X1 port map( A1 => IRAM_ENABLE_port, A2 => IRAM_ADDRESS_2_port
                           , ZN => n4439);
   U4066 : INV_X1 port map( A => n4439, ZN => n4441);
   U4067 : AND2_X1 port map( A1 => n4441, A2 => IRAM_ADDRESS_3_port, ZN => 
                           n4448);
   U4068 : NAND2_X1 port map( A1 => n4448, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n4447);
   U4069 : NOR2_X1 port map( A1 => n741, A2 => n4447, ZN => n4454);
   U4070 : AOI211_X1 port map( C1 => n741, C2 => n4447, A => n4454, B => n4442,
                           ZN => n4295);
   U4071 : OR2_X1 port map( A1 => n4296, A2 => n4295, ZN => 
                           datapath_i_fetch_stage_dp_n32);
   U4072 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_7_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_7_port, ZN => 
                           n4297);
   U4073 : OAI21_X1 port map( B1 => n705, B2 => n4533, A => n4297, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_7_port);
   U4074 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_6_port, ZN => 
                           n4298);
   U4075 : OAI21_X1 port map( B1 => n732, B2 => n4348, A => n4298, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U4076 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_7_port, ZN
                           => n4299);
   U4077 : NAND2_X1 port map( A1 => n4452, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, ZN => 
                           n4451);
   U4078 : NOR2_X1 port map( A1 => n4299, A2 => n4451, ZN => n4458);
   U4079 : AOI211_X1 port map( C1 => n4299, C2 => n4451, A => n4490, B => n4458
                           , ZN => n4301);
   U4080 : NAND2_X1 port map( A1 => n4454, A2 => IRAM_ADDRESS_6_port, ZN => 
                           n4453);
   U4081 : NOR2_X1 port map( A1 => n742, A2 => n4453, ZN => n4460);
   U4082 : INV_X1 port map( A => n4539, ZN => n4536);
   U4083 : AOI211_X1 port map( C1 => n742, C2 => n4453, A => n4460, B => n4536,
                           ZN => n4300);
   U4084 : OR2_X1 port map( A1 => n4301, A2 => n4300, ZN => 
                           datapath_i_fetch_stage_dp_n30);
   U4085 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_9_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_9_port, ZN => 
                           n4302);
   U4086 : OAI21_X1 port map( B1 => n707, B2 => n4533, A => n4302, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_9_port);
   U4087 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_8_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_8_port, ZN => 
                           n4303);
   U4088 : OAI21_X1 port map( B1 => n706, B2 => n4348, A => n4303, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U4089 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_9_port, ZN
                           => n4304);
   U4090 : NAND2_X1 port map( A1 => n4458, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, ZN => 
                           n4457);
   U4091 : NOR2_X1 port map( A1 => n4304, A2 => n4457, ZN => n4464);
   U4092 : AOI211_X1 port map( C1 => n4304, C2 => n4457, A => n4539, B => n4464
                           , ZN => n4306);
   U4093 : NAND2_X1 port map( A1 => n4460, A2 => IRAM_ADDRESS_8_port, ZN => 
                           n4459);
   U4094 : NOR2_X1 port map( A1 => n743, A2 => n4459, ZN => n4466);
   U4095 : AOI211_X1 port map( C1 => n743, C2 => n4459, A => n4466, B => n4536,
                           ZN => n4305);
   U4096 : OR2_X1 port map( A1 => n4306, A2 => n4305, ZN => 
                           datapath_i_fetch_stage_dp_n28);
   U4097 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_11_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_11_port, ZN => 
                           n4307);
   U4098 : OAI21_X1 port map( B1 => n709, B2 => n4348, A => n4307, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_11_port);
   U4099 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_10_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_10_port, ZN => 
                           n4308);
   U4100 : OAI21_X1 port map( B1 => n708, B2 => n4348, A => n4308, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U4101 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_11_port, 
                           ZN => n4309);
   U4102 : NAND2_X1 port map( A1 => n4464, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, ZN => 
                           n4463);
   U4103 : NOR2_X1 port map( A1 => n4309, A2 => n4463, ZN => n4470);
   U4104 : AOI211_X1 port map( C1 => n4309, C2 => n4463, A => n4539, B => n4470
                           , ZN => n4311);
   U4105 : NAND2_X1 port map( A1 => n4466, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n4465);
   U4106 : NOR2_X1 port map( A1 => n744, A2 => n4465, ZN => n4472);
   U4107 : AOI211_X1 port map( C1 => n744, C2 => n4465, A => n4472, B => n4442,
                           ZN => n4310);
   U4108 : OR2_X1 port map( A1 => n4311, A2 => n4310, ZN => 
                           datapath_i_fetch_stage_dp_n26);
   U4109 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_13_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_13_port, ZN => 
                           n4312);
   U4110 : OAI21_X1 port map( B1 => n711, B2 => n4533, A => n4312, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_13_port);
   U4111 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_12_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_12_port, ZN => 
                           n4313);
   U4112 : OAI21_X1 port map( B1 => n710, B2 => n4348, A => n4313, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U4113 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_13_port, 
                           ZN => n4314);
   U4114 : NAND2_X1 port map( A1 => n4470, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, ZN => 
                           n4469);
   U4115 : NOR2_X1 port map( A1 => n4314, A2 => n4469, ZN => n4476);
   U4116 : AOI211_X1 port map( C1 => n4314, C2 => n4469, A => n4539, B => n4476
                           , ZN => n4316);
   U4117 : NAND2_X1 port map( A1 => n4472, A2 => IRAM_ADDRESS_12_port, ZN => 
                           n4471);
   U4118 : NOR2_X1 port map( A1 => n752, A2 => n4471, ZN => n4478);
   U4119 : AOI211_X1 port map( C1 => n752, C2 => n4471, A => n4478, B => n4442,
                           ZN => n4315);
   U4120 : OR2_X1 port map( A1 => n4316, A2 => n4315, ZN => 
                           datapath_i_fetch_stage_dp_n24);
   U4121 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_15_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_15_port, ZN => 
                           n4317);
   U4122 : OAI21_X1 port map( B1 => n713, B2 => n4348, A => n4317, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_15_port);
   U4123 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_14_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_14_port, ZN => 
                           n4318);
   U4124 : OAI21_X1 port map( B1 => n712, B2 => n4348, A => n4318, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U4125 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_15_port, 
                           ZN => n4319);
   U4126 : NAND2_X1 port map( A1 => n4476, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, ZN => 
                           n4475);
   U4127 : NOR2_X1 port map( A1 => n4319, A2 => n4475, ZN => n4482);
   U4128 : AOI211_X1 port map( C1 => n4319, C2 => n4475, A => n4490, B => n4482
                           , ZN => n4321);
   U4129 : NAND2_X1 port map( A1 => n4478, A2 => IRAM_ADDRESS_14_port, ZN => 
                           n4477);
   U4130 : NOR2_X1 port map( A1 => n745, A2 => n4477, ZN => n4484);
   U4131 : AOI211_X1 port map( C1 => n745, C2 => n4477, A => n4484, B => n4442,
                           ZN => n4320);
   U4132 : OR2_X1 port map( A1 => n4321, A2 => n4320, ZN => 
                           datapath_i_fetch_stage_dp_n22);
   U4133 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_17_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_17_port, ZN => 
                           n4322);
   U4134 : OAI21_X1 port map( B1 => n715, B2 => n4533, A => n4322, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_17_port);
   U4135 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_16_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_16_port, ZN => 
                           n4323);
   U4136 : OAI21_X1 port map( B1 => n714, B2 => n4348, A => n4323, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U4137 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_17_port, 
                           ZN => n4324);
   U4138 : NAND2_X1 port map( A1 => n4482, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, ZN => 
                           n4481);
   U4139 : NOR2_X1 port map( A1 => n4324, A2 => n4481, ZN => n4488);
   U4140 : AOI211_X1 port map( C1 => n4324, C2 => n4481, A => n4490, B => n4488
                           , ZN => n4326);
   U4141 : NAND2_X1 port map( A1 => n4484, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n4483);
   U4142 : NOR2_X1 port map( A1 => n746, A2 => n4483, ZN => n4491);
   U4143 : AOI211_X1 port map( C1 => n746, C2 => n4483, A => n4491, B => n4536,
                           ZN => n4325);
   U4144 : OR2_X1 port map( A1 => n4326, A2 => n4325, ZN => 
                           datapath_i_fetch_stage_dp_n20);
   U4145 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_19_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_19_port, ZN => 
                           n4327);
   U4146 : OAI21_X1 port map( B1 => n717, B2 => n4348, A => n4327, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_19_port);
   U4147 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_18_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_18_port, ZN => 
                           n4328);
   U4148 : OAI21_X1 port map( B1 => n716, B2 => n4348, A => n4328, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U4149 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_19_port, 
                           ZN => n4329);
   U4150 : NAND2_X1 port map( A1 => n4488, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, ZN => 
                           n4487);
   U4151 : NOR2_X1 port map( A1 => n4329, A2 => n4487, ZN => n4495);
   U4152 : AOI211_X1 port map( C1 => n4329, C2 => n4487, A => n4490, B => n4495
                           , ZN => n4331);
   U4153 : NAND2_X1 port map( A1 => n4491, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n4489);
   U4154 : NOR2_X1 port map( A1 => n747, A2 => n4489, ZN => n4497);
   U4155 : AOI211_X1 port map( C1 => n747, C2 => n4489, A => n4497, B => n4536,
                           ZN => n4330);
   U4156 : OR2_X1 port map( A1 => n4331, A2 => n4330, ZN => 
                           datapath_i_fetch_stage_dp_n18);
   U4157 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_21_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_21_port, ZN => 
                           n4332);
   U4158 : OAI21_X1 port map( B1 => n719, B2 => n4533, A => n4332, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_21_port);
   U4159 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_20_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_20_port, ZN => 
                           n4333);
   U4160 : OAI21_X1 port map( B1 => n718, B2 => n4348, A => n4333, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U4161 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_21_port, 
                           ZN => n4334);
   U4162 : NAND2_X1 port map( A1 => n4495, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, ZN => 
                           n4494);
   U4163 : NOR2_X1 port map( A1 => n4334, A2 => n4494, ZN => n4501);
   U4164 : AOI211_X1 port map( C1 => n4334, C2 => n4494, A => n4490, B => n4501
                           , ZN => n4336);
   U4165 : NAND2_X1 port map( A1 => n4497, A2 => IRAM_ADDRESS_20_port, ZN => 
                           n4496);
   U4166 : NOR2_X1 port map( A1 => n748, A2 => n4496, ZN => n4503);
   U4167 : AOI211_X1 port map( C1 => n748, C2 => n4496, A => n4503, B => n4536,
                           ZN => n4335);
   U4168 : OR2_X1 port map( A1 => n4336, A2 => n4335, ZN => 
                           datapath_i_fetch_stage_dp_n16);
   U4169 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_23_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_23_port, ZN => 
                           n4337);
   U4170 : OAI21_X1 port map( B1 => n721, B2 => n4348, A => n4337, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_23_port);
   U4171 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_22_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_22_port, ZN => 
                           n4338);
   U4172 : OAI21_X1 port map( B1 => n720, B2 => n4348, A => n4338, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U4173 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_23_port, 
                           ZN => n4339);
   U4174 : NAND2_X1 port map( A1 => n4501, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, ZN => 
                           n4500);
   U4175 : NOR2_X1 port map( A1 => n4339, A2 => n4500, ZN => n4507);
   U4176 : AOI211_X1 port map( C1 => n4339, C2 => n4500, A => n4490, B => n4507
                           , ZN => n4341);
   U4177 : NAND2_X1 port map( A1 => n4503, A2 => IRAM_ADDRESS_22_port, ZN => 
                           n4502);
   U4178 : NOR2_X1 port map( A1 => n749, A2 => n4502, ZN => n4509);
   U4179 : AOI211_X1 port map( C1 => n749, C2 => n4502, A => n4509, B => n4536,
                           ZN => n4340);
   U4180 : OR2_X1 port map( A1 => n4341, A2 => n4340, ZN => 
                           datapath_i_fetch_stage_dp_n14);
   U4181 : AOI22_X1 port map( A1 => n4657, A2 => 
                           datapath_i_alu_output_val_i_25_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_25_port, ZN => 
                           n4342);
   U4182 : OAI21_X1 port map( B1 => n723, B2 => n4533, A => n4342, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_25_port);
   U4183 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_24_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_24_port, ZN => 
                           n4343);
   U4184 : OAI21_X1 port map( B1 => n722, B2 => n4533, A => n4343, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U4185 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_25_port, 
                           ZN => n4344);
   U4186 : NAND2_X1 port map( A1 => n4507, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, ZN => 
                           n4506);
   U4187 : NOR2_X1 port map( A1 => n4344, A2 => n4506, ZN => n4513);
   U4188 : AOI211_X1 port map( C1 => n4344, C2 => n4506, A => n4539, B => n4513
                           , ZN => n4346);
   U4189 : NAND2_X1 port map( A1 => n4509, A2 => IRAM_ADDRESS_24_port, ZN => 
                           n4508);
   U4190 : NOR2_X1 port map( A1 => n750, A2 => n4508, ZN => n4515);
   U4191 : AOI211_X1 port map( C1 => n750, C2 => n4508, A => n4515, B => n4442,
                           ZN => n4345);
   U4192 : OR2_X1 port map( A1 => n4346, A2 => n4345, ZN => 
                           datapath_i_fetch_stage_dp_n12);
   U4193 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_27_port, B1 => n4530, B2
                           => datapath_i_new_pc_value_decode_27_port, ZN => 
                           n4347);
   U4194 : OAI21_X1 port map( B1 => n724, B2 => n4348, A => n4347, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_27_port);
   U4195 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_26_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_26_port, ZN => 
                           n4349);
   U4196 : OAI21_X1 port map( B1 => n691, B2 => n4533, A => n4349, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U4197 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_27_port, 
                           ZN => n4350);
   U4198 : NAND2_X1 port map( A1 => n4513, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, ZN => 
                           n4512);
   U4199 : NOR2_X1 port map( A1 => n4350, A2 => n4512, ZN => n4519);
   U4200 : AOI211_X1 port map( C1 => n4350, C2 => n4512, A => n4490, B => n4519
                           , ZN => n4352);
   U4201 : NAND2_X1 port map( A1 => n4515, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n4514);
   U4202 : NOR2_X1 port map( A1 => n751, A2 => n4514, ZN => n4521);
   U4203 : AOI211_X1 port map( C1 => n751, C2 => n4514, A => n4521, B => n4442,
                           ZN => n4351);
   U4204 : OR2_X1 port map( A1 => n4352, A2 => n4351, ZN => 
                           datapath_i_fetch_stage_dp_n10);
   U4205 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_29_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_29_port, ZN => 
                           n4353);
   U4206 : OAI21_X1 port map( B1 => n726, B2 => n4533, A => n4353, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_29_port);
   U4207 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_28_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_28_port, ZN => 
                           n4354);
   U4208 : OAI21_X1 port map( B1 => n725, B2 => n4533, A => n4354, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U4209 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_29_port, 
                           ZN => n4355);
   U4210 : NAND2_X1 port map( A1 => n4519, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, ZN => 
                           n4518);
   U4211 : NOR2_X1 port map( A1 => n4355, A2 => n4518, ZN => n4526);
   U4212 : AOI211_X1 port map( C1 => n4355, C2 => n4518, A => n4490, B => n4526
                           , ZN => n4357);
   U4213 : NAND2_X1 port map( A1 => n4521, A2 => IRAM_ADDRESS_28_port, ZN => 
                           n4520);
   U4214 : NOR2_X1 port map( A1 => n753, A2 => n4520, ZN => n4527);
   U4215 : AOI211_X1 port map( C1 => n753, C2 => n4520, A => n4527, B => n4536,
                           ZN => n4356);
   U4216 : OR2_X1 port map( A1 => n4357, A2 => n4356, ZN => 
                           datapath_i_fetch_stage_dp_n4);
   U4217 : AOI221_X1 port map( B1 => n4541, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n4542, C2 =>
                           curr_instruction_to_cu_i_15_port, A => n4674, ZN => 
                           n4358);
   U4218 : INV_X1 port map( A => n4358, ZN => n4279);
   U4219 : INV_X1 port map( A => n4363, ZN => n4432);
   U4220 : NOR3_X1 port map( A1 => n737, A2 => curr_instruction_to_cu_i_31_port
                           , A3 => n4368, ZN => n4406);
   U4221 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           n4658, A3 => n4655, A4 => n4669, ZN => n4366);
   U4222 : AOI21_X1 port map( B1 => n4664, B2 => n4656, A => n4366, ZN => n4386
                           );
   U4223 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           curr_instruction_to_cu_i_30_port, A3 => n4359, ZN =>
                           n4401);
   U4224 : NAND3_X1 port map( A1 => n4360, A2 => n4655, A3 => n4656, ZN => 
                           n4419);
   U4225 : NAND2_X1 port map( A1 => n4401, A2 => n4419, ZN => n4396);
   U4226 : NOR3_X1 port map( A1 => n4406, A2 => n4386, A3 => n4396, ZN => n4423
                           );
   U4227 : OAI222_X1 port map( A1 => n4656, A2 => n4586, B1 => n4390, B2 => 
                           n4374, C1 => n4432, C2 => n4423, ZN => n311);
   U4228 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n311, ZN => 
                           cu_i_cmd_word_1_port);
   U4229 : OAI22_X1 port map( A1 => n4663, A2 => cu_i_cw3_6_port, B1 => 
                           cu_i_cw2_6_port, B2 => n704, ZN => n4361);
   U4230 : INV_X1 port map( A => n4361, ZN => n4282);
   U4231 : NOR2_X1 port map( A1 => n4587, A2 => n4656, ZN => 
                           cu_i_cmd_word_7_port);
   U4232 : OAI21_X1 port map( B1 => n4368, B2 => n4362, A => n4423, ZN => n4421
                           );
   U4233 : AOI211_X1 port map( C1 => n4363, C2 => n4421, A => 
                           cu_i_cmd_word_4_port, B => cu_i_cmd_word_7_port, ZN 
                           => n4373);
   U4234 : AND2_X1 port map( A1 => n4373, A2 => n4586, ZN => n4612);
   U4235 : INV_X1 port map( A => n4612, ZN => n4675);
   U4236 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_2_port, B1
                           => cu_i_cw1_2_port, B2 => n4663, ZN => n4381);
   U4237 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_1_port, B1
                           => cu_i_cw1_1_port, B2 => n4436, ZN => n4379);
   U4238 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_3_port, B1
                           => cu_i_cw1_3_port, B2 => n4663, ZN => n4376);
   U4239 : AOI21_X1 port map( B1 => n4381, B2 => n4379, A => n4376, ZN => n4364
                           );
   U4240 : INV_X1 port map( A => n4376, ZN => n4380);
   U4241 : OAI211_X1 port map( C1 => n4377, C2 => n4379, A => n4380, B => n4381
                           , ZN => n4365);
   U4242 : INV_X1 port map( A => n4365, ZN => n4281);
   U4243 : INV_X1 port map( A => n4426, ZN => n4428);
   U4244 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_1_port, A2 => 
                           curr_instruction_to_cu_i_4_port, A3 => n4672, A4 => 
                           n4428, ZN => n4400);
   U4245 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           n4400, ZN => n4388);
   U4246 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => n4666
                           , A3 => n4388, ZN => n4372);
   U4247 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n4656, A3 => n4366, ZN => n4371);
   U4248 : OAI21_X1 port map( B1 => n4368, B2 => n4419, A => n4367, ZN => n4370
                           );
   U4249 : NAND2_X1 port map( A1 => n4670, A2 => n4660, ZN => n4394);
   U4250 : NOR4_X1 port map( A1 => n4661, A2 => n4428, A3 => n4394, A4 => 
                           curr_instruction_to_cu_i_0_port, ZN => n4397);
   U4251 : INV_X1 port map( A => n4397, ZN => n4402);
   U4252 : OAI221_X1 port map( B1 => n4402, B2 => 
                           curr_instruction_to_cu_i_5_port, C1 => n4402, C2 => 
                           curr_instruction_to_cu_i_1_port, A => n4401, ZN => 
                           n4369);
   U4253 : OR4_X1 port map( A1 => n4372, A2 => n4371, A3 => n4370, A4 => n4369,
                           ZN => cu_i_N265);
   U4254 : NAND2_X1 port map( A1 => n4373, A2 => n4541, ZN => enable_rf_i);
   U4255 : INV_X1 port map( A => n4390, ZN => n4416);
   U4256 : NAND2_X1 port map( A1 => n4374, A2 => n4416, ZN => n4414);
   U4257 : INV_X1 port map( A => n4612, ZN => n4676);
   U4258 : AND2_X1 port map( A1 => n4676, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U4259 : INV_X1 port map( A => n4375, ZN => DRAM_READNOTWRITE);
   U4260 : AOI22_X1 port map( A1 => n704, A2 => n4612, B1 => n2319, B2 => n4436
                           , ZN => n4615);
   U4261 : CLKBUF_X1 port map( A => n4615, Z => n4617);
   U4262 : MUX2_X1 port map( A => datapath_i_val_b_i_2_port, B => 
                           datapath_i_val_immediate_i_2_port, S => n4617, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U4263 : AOI21_X1 port map( B1 => n4381, B2 => n4377, A => n4376, ZN => n4378
                           );
   U4264 : NOR2_X1 port map( A1 => n4379, A2 => n4378, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U4265 : NOR2_X1 port map( A1 => n4381, A2 => n4380, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U4266 : NOR2_X1 port map( A1 => n4659, A2 => n4414, ZN => cu_i_N273);
   U4267 : INV_X1 port map( A => n4414, ZN => n4544);
   U4268 : AOI221_X1 port map( B1 => cu_i_n25, B2 => n4544, C1 => cu_i_n26, C2 
                           => n4544, A => cu_i_N273, ZN => n4382);
   U4269 : INV_X1 port map( A => n4382, ZN => n4385);
   U4270 : NOR2_X1 port map( A1 => cu_i_n125, A2 => n4414, ZN => n4383);
   U4271 : NAND2_X1 port map( A1 => n4383, A2 => n4665, ZN => n4412);
   U4272 : NOR2_X1 port map( A1 => cu_i_n25, A2 => n4412, ZN => n4384);
   U4273 : MUX2_X1 port map( A => n4385, B => n4384, S => cu_i_n124, Z => 
                           cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U4275 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => 
                           curr_instruction_to_cu_i_0_port, ZN => n4389);
   U4276 : INV_X1 port map( A => n4386, ZN => n4387);
   U4277 : OAI21_X1 port map( B1 => n4389, B2 => n4388, A => n4387, ZN => 
                           cu_i_N267);
   U4278 : MUX2_X1 port map( A => datapath_i_val_b_i_0_port, B => 
                           datapath_i_val_immediate_i_0_port, S => n4615, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U4279 : MUX2_X1 port map( A => datapath_i_val_b_i_1_port, B => 
                           datapath_i_val_immediate_i_1_port, S => n4617, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U4280 : NAND2_X1 port map( A1 => n4612, A2 => n4390, ZN => cu_i_N278);
   U4281 : MUX2_X1 port map( A => datapath_i_val_b_i_3_port, B => 
                           datapath_i_val_immediate_i_3_port, S => n4615, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U4282 : NOR2_X1 port map( A1 => n4663, A2 => n1152, ZN => n4391);
   U4283 : NOR2_X1 port map( A1 => n704, A2 => cu_i_cw1_4_port, ZN => n4420);
   U4284 : NOR2_X1 port map( A1 => n4391, A2 => n4420, ZN => n4392);
   U4285 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n4392, ZN => n4654);
   U4286 : INV_X1 port map( A => n4392, ZN => n4639);
   U4287 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n4639, ZN => n4652);
   U4288 : CLKBUF_X1 port map( A => n4652, Z => n4641);
   U4289 : CLKBUF_X1 port map( A => n4639, Z => n4651);
   U4290 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_26_port, B2 => 
                           n4651, ZN => n4393);
   U4291 : OAI21_X1 port map( B1 => n691, B2 => n4643, A => n4393, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U4292 : NOR2_X1 port map( A1 => n4395, A2 => n4394, ZN => n4415);
   U4293 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => 
                           n4400, B1 => n4426, B2 => n4415, ZN => n4399);
   U4294 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n4396, B1 => n4406, B2 => n4656, ZN => n4398);
   U4295 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_1_port, A2 => 
                           n4397, ZN => n4407);
   U4296 : OAI211_X1 port map( C1 => curr_instruction_to_cu_i_0_port, C2 => 
                           n4399, A => n4398, B => n4407, ZN => cu_i_N264);
   U4297 : NAND2_X1 port map( A1 => n4400, A2 => n4660, ZN => n4409);
   U4298 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           n4656, ZN => n4405);
   U4299 : NOR3_X1 port map( A1 => n4664, A2 => n4658, A3 => n4419, ZN => n4404
                           );
   U4300 : OAI21_X1 port map( B1 => curr_instruction_to_cu_i_5_port, B2 => 
                           n4402, A => n4401, ZN => n4403);
   U4301 : AOI211_X1 port map( C1 => n4406, C2 => n4405, A => n4404, B => n4403
                           , ZN => n4408);
   U4302 : OAI211_X1 port map( C1 => n4410, C2 => n4409, A => n4408, B => n4407
                           , ZN => cu_i_N266);
   U4303 : NAND2_X1 port map( A1 => n704, A2 => n4414, ZN => cu_i_N274);
   U4304 : AOI221_X1 port map( B1 => cu_i_n125, B2 => cu_i_n26, C1 => n4659, C2
                           => n4665, A => n4414, ZN => cu_i_N275);
   U4305 : OAI21_X1 port map( B1 => cu_i_n26, B2 => cu_i_n125, A => n4544, ZN 
                           => n4411);
   U4306 : AOI22_X1 port map( A1 => cu_i_n25, A2 => n4412, B1 => n4411, B2 => 
                           n4671, ZN => cu_i_N276);
   U4307 : INV_X1 port map( A => n4413, ZN => n4545);
   U4308 : AOI211_X1 port map( C1 => n704, C2 => cu_i_n145, A => n4545, B => 
                           n4414, ZN => cu_i_N279);
   U4309 : NAND4_X1 port map( A1 => n4416, A2 => n4415, A3 => n4661, A4 => 
                           n4666, ZN => n4417);
   U4310 : OAI21_X1 port map( B1 => n4419, B2 => n4418, A => n4417, ZN => 
                           cu_i_cmd_word_8_port);
   U4311 : MUX2_X1 port map( A => cu_i_cmd_word_8_port, B => cu_i_cw1_12_port, 
                           S => n4436, Z => alu_cin_i);
   U4312 : AOI21_X1 port map( B1 => n756, B2 => n704, A => n4420, ZN => 
                           cu_i_cw1_i_4_port);
   U4313 : MUX2_X1 port map( A => cu_i_cw2_7_port, B => cu_i_cw1_7_port, S => 
                           n4663, Z => cu_i_cw1_i_7_port);
   U4314 : MUX2_X1 port map( A => cu_i_cw2_8_port, B => cu_i_cw1_8_port, S => 
                           n4663, Z => cu_i_cw1_i_8_port);
   U4315 : INV_X1 port map( A => n4421, ZN => n4429);
   U4316 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_14_port, A2 => 
                           curr_instruction_to_cu_i_15_port, A3 => 
                           curr_instruction_to_cu_i_11_port, A4 => 
                           curr_instruction_to_cu_i_12_port, ZN => n4422);
   U4317 : NAND2_X1 port map( A1 => n740, A2 => n4422, ZN => n4427);
   U4318 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_19_port, A2 => 
                           curr_instruction_to_cu_i_20_port, A3 => 
                           curr_instruction_to_cu_i_16_port, A4 => 
                           curr_instruction_to_cu_i_17_port, ZN => n4424);
   U4319 : AOI21_X1 port map( B1 => n697, B2 => n4424, A => n4423, ZN => n4425)
                           ;
   U4320 : AOI221_X1 port map( B1 => n4429, B2 => n4428, C1 => n4427, C2 => 
                           n4426, A => n4425, ZN => n4433);
   U4321 : OAI211_X1 port map( C1 => n4433, C2 => n4432, A => n4431, B => n4430
                           , ZN => cu_i_n209);
   U4322 : NOR2_X1 port map( A1 => cu_i_n123, A2 => cu_i_n23, ZN => cu_i_n210);
   U4323 : AOI22_X1 port map( A1 => n704, A2 => n699, B1 => n4673, B2 => n4663,
                           ZN => cu_i_n131);
   U4324 : MUX2_X1 port map( A => cu_i_cw2_6_port, B => cu_i_cw1_6_port, S => 
                           n4436, Z => cu_i_n127);
   U4325 : MUX2_X1 port map( A => cu_i_cw2_5_port, B => cu_i_cw1_5_port, S => 
                           n4436, Z => cu_i_n126);
   U4326 : MUX2_X1 port map( A => curr_instruction_to_cu_i_31_port, B => 
                           IRAM_DATA(31), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n69);
   U4327 : MUX2_X1 port map( A => curr_instruction_to_cu_i_30_port, B => 
                           IRAM_DATA(30), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n68);
   U4328 : MUX2_X1 port map( A => n4655, B => IRAM_DATA(29), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n67);
   U4329 : MUX2_X1 port map( A => curr_instruction_to_cu_i_28_port, B => 
                           IRAM_DATA(28), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n66);
   U4330 : MUX2_X1 port map( A => curr_instruction_to_cu_i_27_port, B => 
                           IRAM_DATA(27), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n65);
   U4331 : MUX2_X1 port map( A => curr_instruction_to_cu_i_26_port, B => 
                           IRAM_DATA(26), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n64);
   U4332 : MUX2_X1 port map( A => datapath_i_n9, B => IRAM_DATA(25), S => n4436
                           , Z => datapath_i_fetch_stage_dp_n63);
   U4333 : MUX2_X1 port map( A => datapath_i_n10, B => IRAM_DATA(24), S => 
                           n4436, Z => datapath_i_fetch_stage_dp_n62);
   U4334 : MUX2_X1 port map( A => datapath_i_n11, B => IRAM_DATA(23), S => 
                           n4436, Z => datapath_i_fetch_stage_dp_n61);
   U4335 : MUX2_X1 port map( A => datapath_i_n12, B => IRAM_DATA(22), S => 
                           n4663, Z => datapath_i_fetch_stage_dp_n60);
   U4336 : MUX2_X1 port map( A => datapath_i_n13, B => IRAM_DATA(21), S => 
                           n4663, Z => datapath_i_fetch_stage_dp_n59);
   U4337 : MUX2_X1 port map( A => curr_instruction_to_cu_i_20_port, B => 
                           IRAM_DATA(20), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n58);
   U4338 : MUX2_X1 port map( A => curr_instruction_to_cu_i_19_port, B => 
                           IRAM_DATA(19), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n57);
   U4339 : NAND2_X1 port map( A1 => n4663, A2 => IRAM_DATA(18), ZN => n4434);
   U4340 : OAI21_X1 port map( B1 => n4663, B2 => n697, A => n4434, ZN => 
                           datapath_i_fetch_stage_dp_n56);
   U4341 : MUX2_X1 port map( A => curr_instruction_to_cu_i_17_port, B => 
                           IRAM_DATA(17), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n55);
   U4342 : MUX2_X1 port map( A => curr_instruction_to_cu_i_16_port, B => 
                           IRAM_DATA(16), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n54);
   U4343 : MUX2_X1 port map( A => curr_instruction_to_cu_i_15_port, B => 
                           IRAM_DATA(15), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n53);
   U4344 : MUX2_X1 port map( A => curr_instruction_to_cu_i_14_port, B => 
                           IRAM_DATA(14), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n52);
   U4345 : NAND2_X1 port map( A1 => n4663, A2 => IRAM_DATA(13), ZN => n4435);
   U4346 : OAI21_X1 port map( B1 => n4436, B2 => n740, A => n4435, ZN => 
                           datapath_i_fetch_stage_dp_n51);
   U4347 : MUX2_X1 port map( A => curr_instruction_to_cu_i_12_port, B => 
                           IRAM_DATA(12), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n50);
   U4348 : MUX2_X1 port map( A => curr_instruction_to_cu_i_11_port, B => 
                           IRAM_DATA(11), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n49);
   U4349 : MUX2_X1 port map( A => datapath_i_n14, B => IRAM_DATA(10), S => 
                           n4436, Z => datapath_i_fetch_stage_dp_n48);
   U4350 : MUX2_X1 port map( A => datapath_i_n15, B => IRAM_DATA(9), S => n4436
                           , Z => datapath_i_fetch_stage_dp_n47);
   U4351 : MUX2_X1 port map( A => datapath_i_n16, B => IRAM_DATA(8), S => n4663
                           , Z => datapath_i_fetch_stage_dp_n46);
   U4352 : MUX2_X1 port map( A => datapath_i_n17, B => IRAM_DATA(7), S => n4436
                           , Z => datapath_i_fetch_stage_dp_n45);
   U4353 : MUX2_X1 port map( A => datapath_i_n18, B => IRAM_DATA(6), S => n4436
                           , Z => datapath_i_fetch_stage_dp_n44);
   U4354 : MUX2_X1 port map( A => curr_instruction_to_cu_i_5_port, B => 
                           IRAM_DATA(5), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n43);
   U4355 : MUX2_X1 port map( A => curr_instruction_to_cu_i_4_port, B => 
                           IRAM_DATA(4), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n42);
   U4356 : MUX2_X1 port map( A => curr_instruction_to_cu_i_3_port, B => 
                           IRAM_DATA(3), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n41);
   U4357 : MUX2_X1 port map( A => curr_instruction_to_cu_i_2_port, B => 
                           IRAM_DATA(2), S => n4663, Z => 
                           datapath_i_fetch_stage_dp_n40);
   U4358 : MUX2_X1 port map( A => curr_instruction_to_cu_i_1_port, B => 
                           IRAM_DATA(1), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n39);
   U4359 : MUX2_X1 port map( A => curr_instruction_to_cu_i_0_port, B => 
                           IRAM_DATA(0), S => n4436, Z => 
                           datapath_i_fetch_stage_dp_n38);
   U4360 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_0_port, ZN => 
                           n4437);
   U4361 : OAI21_X1 port map( B1 => n733, B2 => n4533, A => n4437, ZN => 
                           datapath_i_fetch_stage_dp_N5);
   U4362 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N39_port, B => 
                           datapath_i_fetch_stage_dp_N5, S => n4442, Z => 
                           datapath_i_fetch_stage_dp_n37);
   U4363 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_1_port, B1 => n4524, B2 
                           => datapath_i_new_pc_value_decode_1_port, ZN => 
                           n4438);
   U4364 : OAI21_X1 port map( B1 => n734, B2 => n4533, A => n4438, ZN => 
                           datapath_i_fetch_stage_dp_N6);
   U4365 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N40_port, B => 
                           datapath_i_fetch_stage_dp_N6, S => n4442, Z => 
                           datapath_i_fetch_stage_dp_n36);
   U4366 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port
                           , A => n4439, ZN => n4440);
   U4367 : AOI22_X1 port map( A1 => n4539, A2 => n4440, B1 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B2 => 
                           n4536, ZN => datapath_i_fetch_stage_dp_n35);
   U4368 : OAI21_X1 port map( B1 => n4441, B2 => IRAM_ADDRESS_3_port, A => 
                           n4490, ZN => n4444);
   U4369 : AND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_2_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, ZN
                           => n4446);
   U4370 : OAI21_X1 port map( B1 => datapath_i_new_pc_value_mem_stage_i_2_port,
                           B2 => datapath_i_new_pc_value_mem_stage_i_3_port, A 
                           => n4442, ZN => n4443);
   U4371 : OAI22_X1 port map( A1 => n4448, A2 => n4444, B1 => n4446, B2 => 
                           n4443, ZN => datapath_i_fetch_stage_dp_n34);
   U4372 : OAI211_X1 port map( C1 => n4446, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n4536, B => n4445, ZN => n4450);
   U4373 : OAI211_X1 port map( C1 => n4448, C2 => IRAM_ADDRESS_4_port, A => 
                           n4539, B => n4447, ZN => n4449);
   U4374 : NAND2_X1 port map( A1 => n4450, A2 => n4449, ZN => 
                           datapath_i_fetch_stage_dp_n33);
   U4375 : OAI211_X1 port map( C1 => n4452, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, A => 
                           n4536, B => n4451, ZN => n4456);
   U4376 : OAI211_X1 port map( C1 => n4454, C2 => IRAM_ADDRESS_6_port, A => 
                           n4539, B => n4453, ZN => n4455);
   U4377 : NAND2_X1 port map( A1 => n4456, A2 => n4455, ZN => 
                           datapath_i_fetch_stage_dp_n31);
   U4378 : OAI211_X1 port map( C1 => n4458, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, A => 
                           n4536, B => n4457, ZN => n4462);
   U4379 : OAI211_X1 port map( C1 => n4460, C2 => IRAM_ADDRESS_8_port, A => 
                           n4539, B => n4459, ZN => n4461);
   U4380 : NAND2_X1 port map( A1 => n4462, A2 => n4461, ZN => 
                           datapath_i_fetch_stage_dp_n29);
   U4381 : OAI211_X1 port map( C1 => n4464, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, A => 
                           n4536, B => n4463, ZN => n4468);
   U4382 : OAI211_X1 port map( C1 => n4466, C2 => IRAM_ADDRESS_10_port, A => 
                           n4539, B => n4465, ZN => n4467);
   U4383 : NAND2_X1 port map( A1 => n4468, A2 => n4467, ZN => 
                           datapath_i_fetch_stage_dp_n27);
   U4384 : OAI211_X1 port map( C1 => n4470, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, A => 
                           n4536, B => n4469, ZN => n4474);
   U4385 : OAI211_X1 port map( C1 => n4472, C2 => IRAM_ADDRESS_12_port, A => 
                           n4490, B => n4471, ZN => n4473);
   U4386 : NAND2_X1 port map( A1 => n4474, A2 => n4473, ZN => 
                           datapath_i_fetch_stage_dp_n25);
   U4387 : OAI211_X1 port map( C1 => n4476, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, A => 
                           n4536, B => n4475, ZN => n4480);
   U4388 : OAI211_X1 port map( C1 => n4478, C2 => IRAM_ADDRESS_14_port, A => 
                           n4490, B => n4477, ZN => n4479);
   U4389 : NAND2_X1 port map( A1 => n4480, A2 => n4479, ZN => 
                           datapath_i_fetch_stage_dp_n23);
   U4390 : OAI211_X1 port map( C1 => n4482, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, A => 
                           n4536, B => n4481, ZN => n4486);
   U4391 : OAI211_X1 port map( C1 => n4484, C2 => IRAM_ADDRESS_16_port, A => 
                           n4490, B => n4483, ZN => n4485);
   U4392 : NAND2_X1 port map( A1 => n4486, A2 => n4485, ZN => 
                           datapath_i_fetch_stage_dp_n21);
   U4393 : OAI211_X1 port map( C1 => n4488, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, A => 
                           n4536, B => n4487, ZN => n4493);
   U4394 : OAI211_X1 port map( C1 => n4491, C2 => IRAM_ADDRESS_18_port, A => 
                           n4490, B => n4489, ZN => n4492);
   U4395 : NAND2_X1 port map( A1 => n4493, A2 => n4492, ZN => 
                           datapath_i_fetch_stage_dp_n19);
   U4396 : OAI211_X1 port map( C1 => n4495, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, A => 
                           n4536, B => n4494, ZN => n4499);
   U4397 : OAI211_X1 port map( C1 => n4497, C2 => IRAM_ADDRESS_20_port, A => 
                           n4539, B => n4496, ZN => n4498);
   U4398 : NAND2_X1 port map( A1 => n4499, A2 => n4498, ZN => 
                           datapath_i_fetch_stage_dp_n17);
   U4399 : OAI211_X1 port map( C1 => n4501, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, A => 
                           n4536, B => n4500, ZN => n4505);
   U4400 : OAI211_X1 port map( C1 => n4503, C2 => IRAM_ADDRESS_22_port, A => 
                           n4539, B => n4502, ZN => n4504);
   U4401 : NAND2_X1 port map( A1 => n4505, A2 => n4504, ZN => 
                           datapath_i_fetch_stage_dp_n15);
   U4402 : OAI211_X1 port map( C1 => n4507, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, A => 
                           n4536, B => n4506, ZN => n4511);
   U4403 : OAI211_X1 port map( C1 => n4509, C2 => IRAM_ADDRESS_24_port, A => 
                           n4539, B => n4508, ZN => n4510);
   U4404 : NAND2_X1 port map( A1 => n4511, A2 => n4510, ZN => 
                           datapath_i_fetch_stage_dp_n13);
   U4405 : OAI211_X1 port map( C1 => n4513, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, A => 
                           n4536, B => n4512, ZN => n4517);
   U4406 : OAI211_X1 port map( C1 => n4515, C2 => IRAM_ADDRESS_26_port, A => 
                           n4539, B => n4514, ZN => n4516);
   U4407 : NAND2_X1 port map( A1 => n4517, A2 => n4516, ZN => 
                           datapath_i_fetch_stage_dp_n11);
   U4408 : OAI211_X1 port map( C1 => n4519, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, A => 
                           n4536, B => n4518, ZN => n4523);
   U4409 : OAI211_X1 port map( C1 => n4521, C2 => IRAM_ADDRESS_28_port, A => 
                           n4539, B => n4520, ZN => n4522);
   U4410 : NAND2_X1 port map( A1 => n4523, A2 => n4522, ZN => 
                           datapath_i_fetch_stage_dp_n9);
   U4411 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_30_port, B1 => n4524, B2
                           => datapath_i_new_pc_value_decode_30_port, ZN => 
                           n4525);
   U4412 : OAI21_X1 port map( B1 => n727, B2 => n4533, A => n4525, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   U4413 : NAND2_X1 port map( A1 => n4526, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, ZN => 
                           n4535);
   U4414 : OAI211_X1 port map( C1 => n4526, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, A => 
                           n4536, B => n4535, ZN => n4529);
   U4415 : NAND2_X1 port map( A1 => n4527, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n4534);
   U4416 : OAI211_X1 port map( C1 => n4527, C2 => IRAM_ADDRESS_30_port, A => 
                           n4539, B => n4534, ZN => n4528);
   U4417 : NAND2_X1 port map( A1 => n4529, A2 => n4528, ZN => 
                           datapath_i_fetch_stage_dp_n3);
   U4418 : AOI22_X1 port map( A1 => n4531, A2 => 
                           datapath_i_alu_output_val_i_31_port, B1 => 
                           datapath_i_new_pc_value_decode_31_port, B2 => n4530,
                           ZN => n4532);
   U4419 : OAI21_X1 port map( B1 => n703, B2 => n4533, A => n4532, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_31_port);
   U4420 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n4534, Z => n4538)
                           ;
   U4421 : XOR2_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_31_port, 
                           B => n4535, Z => n4537);
   U4422 : AOI22_X1 port map( A1 => n4539, A2 => n4538, B1 => n4537, B2 => 
                           n4536, ZN => datapath_i_fetch_stage_dp_n2);
   U4423 : OAI21_X1 port map( B1 => n737, B2 => n4540, A => n4541, ZN => 
                           read_rf_p2_i);
   U4424 : OAI221_X1 port map( B1 => n4542, B2 => n697, C1 => n4541, C2 => n740
                           , A => n4586, ZN => datapath_i_decode_stage_dp_n78);
   U4425 : AND4_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           A2 => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           A3 => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           A4 => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ZN => n4543);
   U4426 : AND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           A2 => n4543, ZN => n4559);
   U4427 : INV_X1 port map( A => n4559, ZN => n4568);
   U4428 : CLKBUF_X1 port map( A => n4583, Z => n4573);
   U4429 : NOR2_X1 port map( A1 => n4559, A2 => n4546, ZN => n4582);
   U4430 : CLKBUF_X1 port map( A => n4582, Z => n4572);
   U4431 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_0_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_0_port, ZN => n4547
                           );
   U4432 : OAI21_X1 port map( B1 => n733, B2 => n4568, A => n4547, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U4433 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_1_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_1_port, ZN => n4548
                           );
   U4434 : OAI21_X1 port map( B1 => n734, B2 => n4568, A => n4548, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U4435 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_2_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_2_port, ZN => n4549
                           );
   U4436 : OAI21_X1 port map( B1 => n728, B2 => n4568, A => n4549, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U4437 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_3_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_3_port, ZN => n4550
                           );
   U4438 : OAI21_X1 port map( B1 => n729, B2 => n4568, A => n4550, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U4439 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_4_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_4_port, ZN => n4551
                           );
   U4440 : OAI21_X1 port map( B1 => n730, B2 => n4568, A => n4551, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U4441 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_5_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_5_port, ZN => n4552
                           );
   U4442 : OAI21_X1 port map( B1 => n731, B2 => n4568, A => n4552, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U4443 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_6_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_6_port, ZN => n4553
                           );
   U4444 : OAI21_X1 port map( B1 => n732, B2 => n4568, A => n4553, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U4445 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_7_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_7_port, ZN => n4554
                           );
   U4446 : OAI21_X1 port map( B1 => n705, B2 => n4568, A => n4554, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U4447 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_8_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_8_port, ZN => n4555
                           );
   U4448 : OAI21_X1 port map( B1 => n706, B2 => n4568, A => n4555, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U4449 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_9_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_9_port, ZN => n4556
                           );
   U4450 : OAI21_X1 port map( B1 => n707, B2 => n4568, A => n4556, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U4451 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_10_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_10_port, ZN => 
                           n4557);
   U4452 : OAI21_X1 port map( B1 => n708, B2 => n4568, A => n4557, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U4453 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_11_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_11_port, ZN => 
                           n4558);
   U4454 : OAI21_X1 port map( B1 => n709, B2 => n4568, A => n4558, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U4455 : INV_X1 port map( A => n4559, ZN => n4585);
   U4456 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_12_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_12_port, ZN => 
                           n4560);
   U4457 : OAI21_X1 port map( B1 => n710, B2 => n4585, A => n4560, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U4458 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_13_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_13_port, ZN => 
                           n4561);
   U4459 : OAI21_X1 port map( B1 => n711, B2 => n4568, A => n4561, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U4460 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_14_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_14_port, ZN => 
                           n4562);
   U4461 : OAI21_X1 port map( B1 => n712, B2 => n4585, A => n4562, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U4462 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_15_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_15_port, ZN => 
                           n4563);
   U4463 : OAI21_X1 port map( B1 => n713, B2 => n4568, A => n4563, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U4464 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_16_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_16_port, ZN => 
                           n4564);
   U4465 : OAI21_X1 port map( B1 => n714, B2 => n4585, A => n4564, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U4466 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_17_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_17_port, ZN => 
                           n4565);
   U4467 : OAI21_X1 port map( B1 => n715, B2 => n4568, A => n4565, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U4468 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_18_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_18_port, ZN => 
                           n4566);
   U4469 : OAI21_X1 port map( B1 => n716, B2 => n4585, A => n4566, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U4470 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_19_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_19_port, ZN => 
                           n4567);
   U4471 : OAI21_X1 port map( B1 => n717, B2 => n4568, A => n4567, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U4472 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_20_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_20_port, ZN => 
                           n4569);
   U4473 : OAI21_X1 port map( B1 => n718, B2 => n4585, A => n4569, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U4474 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_21_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_21_port, ZN => 
                           n4570);
   U4475 : OAI21_X1 port map( B1 => n719, B2 => n4585, A => n4570, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U4476 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_22_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_22_port, ZN => 
                           n4571);
   U4477 : OAI21_X1 port map( B1 => n720, B2 => n4585, A => n4571, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U4478 : AOI22_X1 port map( A1 => n4573, A2 => 
                           datapath_i_data_from_memory_i_23_port, B1 => n4572, 
                           B2 => datapath_i_data_from_alu_i_23_port, ZN => 
                           n4574);
   U4479 : OAI21_X1 port map( B1 => n721, B2 => n4585, A => n4574, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U4480 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_24_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_24_port, ZN => 
                           n4575);
   U4481 : OAI21_X1 port map( B1 => n722, B2 => n4585, A => n4575, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U4482 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_25_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_25_port, ZN => 
                           n4576);
   U4483 : OAI21_X1 port map( B1 => n723, B2 => n4585, A => n4576, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U4484 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_26_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_26_port, ZN => 
                           n4577);
   U4485 : OAI21_X1 port map( B1 => n691, B2 => n4585, A => n4577, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U4486 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_27_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_27_port, ZN => 
                           n4578);
   U4487 : OAI21_X1 port map( B1 => n724, B2 => n4585, A => n4578, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U4488 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_28_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_28_port, ZN => 
                           n4579);
   U4489 : OAI21_X1 port map( B1 => n725, B2 => n4585, A => n4579, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U4490 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_29_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_29_port, ZN => 
                           n4580);
   U4491 : OAI21_X1 port map( B1 => n726, B2 => n4585, A => n4580, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U4492 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_30_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_30_port, ZN => 
                           n4581);
   U4493 : OAI21_X1 port map( B1 => n727, B2 => n4585, A => n4581, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U4494 : AOI22_X1 port map( A1 => n4583, A2 => 
                           datapath_i_data_from_memory_i_31_port, B1 => n4582, 
                           B2 => datapath_i_data_from_alu_i_31_port, ZN => 
                           n4584);
   U4495 : OAI21_X1 port map( B1 => n703, B2 => n4585, A => n4584, ZN => 
                           datapath_i_decode_stage_dp_n12);
   U4496 : OAI21_X1 port map( B1 => curr_instruction_to_cu_i_26_port, B2 => 
                           n4587, A => n4586, ZN => cu_i_cmd_word_6_port);
   U4497 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_6_port, B1 => 
                           cu_i_cw1_10_port, B2 => n4663, ZN => n4601);
   U4498 : NOR4_X1 port map( A1 => datapath_i_val_a_i_14_port, A2 => 
                           datapath_i_val_a_i_15_port, A3 => 
                           datapath_i_val_a_i_16_port, A4 => 
                           datapath_i_val_a_i_17_port, ZN => n4591);
   U4499 : NOR4_X1 port map( A1 => datapath_i_val_a_i_18_port, A2 => 
                           datapath_i_val_a_i_19_port, A3 => 
                           datapath_i_val_a_i_20_port, A4 => 
                           datapath_i_val_a_i_21_port, ZN => n4590);
   U4500 : NOR4_X1 port map( A1 => datapath_i_val_a_i_26_port, A2 => 
                           datapath_i_val_a_i_7_port, A3 => 
                           datapath_i_val_a_i_8_port, A4 => 
                           datapath_i_val_a_i_9_port, ZN => n4589);
   U4501 : NOR4_X1 port map( A1 => datapath_i_val_a_i_10_port, A2 => 
                           datapath_i_val_a_i_11_port, A3 => 
                           datapath_i_val_a_i_12_port, A4 => 
                           datapath_i_val_a_i_13_port, ZN => n4588);
   U4502 : NAND4_X1 port map( A1 => n4591, A2 => n4590, A3 => n4589, A4 => 
                           n4588, ZN => n4597);
   U4503 : NOR4_X1 port map( A1 => datapath_i_val_a_i_30_port, A2 => 
                           datapath_i_val_a_i_31_port, A3 => 
                           datapath_i_val_a_i_1_port, A4 => 
                           datapath_i_val_a_i_2_port, ZN => n4595);
   U4504 : NOR4_X1 port map( A1 => datapath_i_val_a_i_3_port, A2 => 
                           datapath_i_val_a_i_4_port, A3 => 
                           datapath_i_val_a_i_5_port, A4 => 
                           datapath_i_val_a_i_6_port, ZN => n4594);
   U4505 : NOR4_X1 port map( A1 => datapath_i_val_a_i_22_port, A2 => 
                           datapath_i_val_a_i_23_port, A3 => 
                           datapath_i_val_a_i_24_port, A4 => 
                           datapath_i_val_a_i_25_port, ZN => n4593);
   U4506 : NOR4_X1 port map( A1 => datapath_i_val_a_i_0_port, A2 => 
                           datapath_i_val_a_i_27_port, A3 => 
                           datapath_i_val_a_i_28_port, A4 => 
                           datapath_i_val_a_i_29_port, ZN => n4592);
   U4507 : NAND4_X1 port map( A1 => n4595, A2 => n4594, A3 => n4593, A4 => 
                           n4592, ZN => n4596);
   U4508 : NOR2_X1 port map( A1 => n4597, A2 => n4596, ZN => n4599);
   U4509 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_7_port, B1 => 
                           cu_i_cw1_11_port, B2 => n4663, ZN => n4598);
   U4510 : NAND2_X1 port map( A1 => n4599, A2 => n4598, ZN => n4600);
   U4511 : OAI22_X1 port map( A1 => n4601, A2 => n4600, B1 => n4599, B2 => 
                           n4598, ZN => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port);
   U4512 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, S 
                           => n4676, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port)
                           ;
   U4513 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port)
                           ;
   U4514 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, S 
                           => n4676, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port)
                           ;
   U4515 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           );
   U4516 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, S 
                           => n4676, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           );
   U4517 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           );
   U4518 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           );
   U4519 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           );
   U4520 : NAND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
                           A2 => n4676, ZN => n4614);
   U4521 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
                           ZN => n4602);
   U4522 : NAND2_X1 port map( A1 => n4614, A2 => n4602, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           );
   U4523 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
                           ZN => n4603);
   U4524 : NAND2_X1 port map( A1 => n4614, A2 => n4603, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           );
   U4525 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
                           ZN => n4604);
   U4526 : NAND2_X1 port map( A1 => n4614, A2 => n4604, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           );
   U4527 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
                           ZN => n4605);
   U4528 : NAND2_X1 port map( A1 => n4614, A2 => n4605, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           );
   U4529 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
                           ZN => n4606);
   U4530 : NAND2_X1 port map( A1 => n4614, A2 => n4606, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           );
   U4531 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
                           ZN => n4607);
   U4532 : NAND2_X1 port map( A1 => n4614, A2 => n4607, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           );
   U4533 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
                           ZN => n4608);
   U4534 : NAND2_X1 port map( A1 => n4614, A2 => n4608, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           );
   U4535 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
                           ZN => n4609);
   U4536 : NAND2_X1 port map( A1 => n4614, A2 => n4609, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           );
   U4537 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
                           ZN => n4610);
   U4538 : NAND2_X1 port map( A1 => n4614, A2 => n4610, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           );
   U4539 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
                           ZN => n4611);
   U4540 : NAND2_X1 port map( A1 => n4614, A2 => n4611, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           );
   U4541 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port)
                           ;
   U4542 : NAND2_X1 port map( A1 => n4612, A2 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
                           ZN => n4613);
   U4543 : NAND2_X1 port map( A1 => n4614, A2 => n4613, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           );
   U4544 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port)
                           ;
   U4545 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port)
                           ;
   U4546 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port)
                           ;
   U4547 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port)
                           ;
   U4548 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port)
                           ;
   U4549 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, S 
                           => n4675, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port)
                           ;
   U4550 : MUX2_X1 port map( A => datapath_i_val_b_i_7_port, B => 
                           datapath_i_val_immediate_i_7_port, S => n4615, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U4551 : MUX2_X1 port map( A => datapath_i_val_b_i_8_port, B => 
                           datapath_i_val_immediate_i_8_port, S => n4615, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U4552 : MUX2_X1 port map( A => datapath_i_val_b_i_9_port, B => 
                           datapath_i_val_immediate_i_9_port, S => n4615, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U4553 : MUX2_X1 port map( A => datapath_i_val_b_i_10_port, B => 
                           datapath_i_val_immediate_i_10_port, S => n4615, Z =>
                           datapath_i_execute_stage_dp_opb_10_port);
   U4554 : MUX2_X1 port map( A => datapath_i_val_b_i_11_port, B => 
                           datapath_i_val_immediate_i_11_port, S => n4615, Z =>
                           datapath_i_execute_stage_dp_opb_11_port);
   U4555 : MUX2_X1 port map( A => datapath_i_val_b_i_12_port, B => 
                           datapath_i_val_immediate_i_12_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_12_port);
   U4556 : MUX2_X1 port map( A => datapath_i_val_b_i_13_port, B => 
                           datapath_i_val_immediate_i_13_port, S => n4615, Z =>
                           datapath_i_execute_stage_dp_opb_13_port);
   U4557 : MUX2_X1 port map( A => datapath_i_val_b_i_14_port, B => 
                           datapath_i_val_immediate_i_14_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_14_port);
   U4558 : MUX2_X1 port map( A => datapath_i_val_b_i_15_port, B => 
                           datapath_i_val_immediate_i_15_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_15_port);
   U4559 : MUX2_X1 port map( A => datapath_i_val_b_i_16_port, B => 
                           datapath_i_val_immediate_i_16_port, S => n4615, Z =>
                           datapath_i_execute_stage_dp_opb_16_port);
   U4560 : MUX2_X1 port map( A => datapath_i_val_b_i_17_port, B => 
                           datapath_i_val_immediate_i_17_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_17_port);
   U4561 : MUX2_X1 port map( A => datapath_i_val_b_i_18_port, B => 
                           datapath_i_val_immediate_i_18_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_18_port);
   U4562 : MUX2_X1 port map( A => datapath_i_val_b_i_19_port, B => 
                           datapath_i_val_immediate_i_19_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_19_port);
   U4563 : MUX2_X1 port map( A => datapath_i_val_b_i_20_port, B => 
                           datapath_i_val_immediate_i_20_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_20_port);
   U4564 : MUX2_X1 port map( A => datapath_i_val_b_i_21_port, B => 
                           datapath_i_val_immediate_i_21_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_21_port);
   U4565 : MUX2_X1 port map( A => datapath_i_val_b_i_22_port, B => 
                           datapath_i_val_immediate_i_22_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_22_port);
   U4566 : MUX2_X1 port map( A => datapath_i_val_b_i_23_port, B => 
                           datapath_i_val_immediate_i_23_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_23_port);
   U4567 : MUX2_X1 port map( A => datapath_i_val_b_i_24_port, B => 
                           datapath_i_val_immediate_i_24_port, S => n4617, Z =>
                           datapath_i_execute_stage_dp_opb_24_port);
   U4568 : NAND2_X1 port map( A1 => n4617, A2 => 
                           datapath_i_val_immediate_i_25_port, ZN => n4616);
   U4569 : OAI21_X1 port map( B1 => n4617, B2 => n758, A => n4616, ZN => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U4570 : OAI21_X1 port map( B1 => n4617, B2 => n759, A => n4616, ZN => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U4571 : OAI21_X1 port map( B1 => n4617, B2 => n760, A => n4616, ZN => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U4572 : OAI21_X1 port map( B1 => n4617, B2 => n761, A => n4616, ZN => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U4573 : OAI21_X1 port map( B1 => n4617, B2 => n762, A => n4616, ZN => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U4574 : OAI21_X1 port map( B1 => n4617, B2 => n763, A => n4616, ZN => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U4575 : OAI21_X1 port map( B1 => n4617, B2 => n764, A => n4616, ZN => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U4576 : MUX2_X1 port map( A => datapath_i_val_b_i_4_port, B => 
                           datapath_i_val_immediate_i_4_port, S => n4617, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U4577 : MUX2_X1 port map( A => datapath_i_val_b_i_5_port, B => 
                           datapath_i_val_immediate_i_5_port, S => n4617, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U4578 : MUX2_X1 port map( A => datapath_i_val_b_i_6_port, B => 
                           datapath_i_val_immediate_i_6_port, S => n4617, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U4579 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_7_port, B2 => 
                           n4639, ZN => n4618);
   U4580 : OAI21_X1 port map( B1 => n705, B2 => n4654, A => n4618, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U4581 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_8_port, B2 => 
                           n4651, ZN => n4619);
   U4582 : OAI21_X1 port map( B1 => n706, B2 => n4643, A => n4619, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U4583 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_9_port, B2 => 
                           n4639, ZN => n4620);
   U4584 : OAI21_X1 port map( B1 => n707, B2 => n4654, A => n4620, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U4585 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_10_port, B2 => 
                           n4651, ZN => n4621);
   U4586 : OAI21_X1 port map( B1 => n708, B2 => n4643, A => n4621, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U4587 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_11_port, B2 => 
                           n4639, ZN => n4622);
   U4588 : OAI21_X1 port map( B1 => n709, B2 => n4654, A => n4622, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U4589 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_12_port, B2 => 
                           n4651, ZN => n4623);
   U4590 : OAI21_X1 port map( B1 => n710, B2 => n4643, A => n4623, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U4591 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_13_port, B2 => 
                           n4639, ZN => n4624);
   U4592 : OAI21_X1 port map( B1 => n711, B2 => n4654, A => n4624, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U4593 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_14_port, B2 => 
                           n4651, ZN => n4625);
   U4594 : OAI21_X1 port map( B1 => n712, B2 => n4643, A => n4625, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U4595 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_15_port, B2 => 
                           n4639, ZN => n4626);
   U4596 : OAI21_X1 port map( B1 => n713, B2 => n4654, A => n4626, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U4597 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_16_port, B2 => 
                           n4639, ZN => n4627);
   U4598 : OAI21_X1 port map( B1 => n714, B2 => n4654, A => n4627, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U4599 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_17_port, B2 => 
                           n4651, ZN => n4628);
   U4600 : OAI21_X1 port map( B1 => n715, B2 => n4654, A => n4628, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U4601 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_18_port, B2 => 
                           n4639, ZN => n4629);
   U4602 : OAI21_X1 port map( B1 => n716, B2 => n4643, A => n4629, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U4603 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_19_port, B2 => 
                           n4651, ZN => n4630);
   U4604 : OAI21_X1 port map( B1 => n717, B2 => n4643, A => n4630, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U4605 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_20_port, B2 => 
                           n4639, ZN => n4631);
   U4606 : OAI21_X1 port map( B1 => n718, B2 => n4643, A => n4631, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U4607 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_21_port, B2 => 
                           n4651, ZN => n4632);
   U4608 : OAI21_X1 port map( B1 => n719, B2 => n4643, A => n4632, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U4609 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_22_port, B2 => 
                           n4639, ZN => n4633);
   U4610 : OAI21_X1 port map( B1 => n720, B2 => n4643, A => n4633, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U4611 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_23_port, B2 => 
                           n4639, ZN => n4634);
   U4612 : OAI21_X1 port map( B1 => n721, B2 => n4643, A => n4634, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U4613 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_24_port, B2 => 
                           n4639, ZN => n4635);
   U4614 : OAI21_X1 port map( B1 => n722, B2 => n4643, A => n4635, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U4615 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_25_port, B2 => 
                           n4639, ZN => n4636);
   U4616 : OAI21_X1 port map( B1 => n723, B2 => n4643, A => n4636, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U4617 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_0_port, B2 => 
                           n4639, ZN => n4637);
   U4618 : OAI21_X1 port map( B1 => n733, B2 => n4643, A => n4637, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U4619 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_27_port, B2 => 
                           n4639, ZN => n4638);
   U4620 : OAI21_X1 port map( B1 => n724, B2 => n4643, A => n4638, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U4621 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_28_port, B2 => 
                           n4639, ZN => n4640);
   U4622 : OAI21_X1 port map( B1 => n725, B2 => n4643, A => n4640, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U4623 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n4641, B1 => datapath_i_val_a_i_29_port, B2 => 
                           n4651, ZN => n4642);
   U4624 : OAI21_X1 port map( B1 => n726, B2 => n4643, A => n4642, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U4625 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_30_port, B2 => 
                           n4651, ZN => n4644);
   U4626 : OAI21_X1 port map( B1 => n727, B2 => n4654, A => n4644, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U4627 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_31_port, B2 => 
                           n4651, ZN => n4645);
   U4628 : OAI21_X1 port map( B1 => n703, B2 => n4654, A => n4645, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U4629 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_1_port, B2 => 
                           n4651, ZN => n4646);
   U4630 : OAI21_X1 port map( B1 => n734, B2 => n4654, A => n4646, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U4631 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_2_port, B2 => 
                           n4651, ZN => n4647);
   U4632 : OAI21_X1 port map( B1 => n728, B2 => n4654, A => n4647, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U4633 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_3_port, B2 => 
                           n4651, ZN => n4648);
   U4634 : OAI21_X1 port map( B1 => n729, B2 => n4654, A => n4648, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U4635 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_4_port, B2 => 
                           n4651, ZN => n4649);
   U4636 : OAI21_X1 port map( B1 => n730, B2 => n4654, A => n4649, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U4637 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_5_port, B2 => 
                           n4651, ZN => n4650);
   U4638 : OAI21_X1 port map( B1 => n731, B2 => n4654, A => n4650, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U4639 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n4652, B1 => datapath_i_val_a_i_6_port, B2 => 
                           n4651, ZN => n4653);
   U4640 : OAI21_X1 port map( B1 => n732, B2 => n4654, A => n4653, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);

end SYN_dlx_rtl;
