`ifndef implemented_instructions.svh
`def implemented_instructions.svh


enum integer [4:0] {
	
} instructions;



`endif // implemented_instructions.svh