
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, dataout_mul_31_port, dataout_mul_30_port, 
      dataout_mul_29_port, dataout_mul_28_port, dataout_mul_27_port, 
      dataout_mul_26_port, dataout_mul_25_port, dataout_mul_24_port, 
      dataout_mul_23_port, dataout_mul_22_port, dataout_mul_21_port, 
      dataout_mul_20_port, dataout_mul_19_port, dataout_mul_18_port, 
      dataout_mul_17_port, dataout_mul_16_port, dataout_mul_15_port, 
      dataout_mul_13_port, dataout_mul_12_port, dataout_mul_11_port, 
      dataout_mul_10_port, dataout_mul_9_port, dataout_mul_8_port, 
      dataout_mul_7_port, dataout_mul_6_port, dataout_mul_5_port, 
      dataout_mul_4_port, dataout_mul_3_port, dataout_mul_2_port, 
      dataout_mul_1_port, dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521
      , N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n553, 
      boothmul_pipelined_i_muxes_in_7_233_port, 
      boothmul_pipelined_i_muxes_in_7_232_port, 
      boothmul_pipelined_i_muxes_in_7_231_port, 
      boothmul_pipelined_i_muxes_in_7_230_port, 
      boothmul_pipelined_i_muxes_in_7_229_port, 
      boothmul_pipelined_i_muxes_in_7_228_port, 
      boothmul_pipelined_i_muxes_in_7_227_port, 
      boothmul_pipelined_i_muxes_in_7_226_port, 
      boothmul_pipelined_i_muxes_in_7_225_port, 
      boothmul_pipelined_i_muxes_in_7_224_port, 
      boothmul_pipelined_i_muxes_in_7_223_port, 
      boothmul_pipelined_i_muxes_in_7_222_port, 
      boothmul_pipelined_i_muxes_in_7_221_port, 
      boothmul_pipelined_i_muxes_in_7_220_port, 
      boothmul_pipelined_i_muxes_in_7_219_port, 
      boothmul_pipelined_i_muxes_in_7_218_port, 
      boothmul_pipelined_i_muxes_in_7_217_port, 
      boothmul_pipelined_i_muxes_in_7_77_port, 
      boothmul_pipelined_i_muxes_in_7_76_port, 
      boothmul_pipelined_i_muxes_in_7_75_port, 
      boothmul_pipelined_i_muxes_in_7_74_port, 
      boothmul_pipelined_i_muxes_in_7_73_port, 
      boothmul_pipelined_i_muxes_in_7_72_port, 
      boothmul_pipelined_i_muxes_in_7_71_port, 
      boothmul_pipelined_i_muxes_in_7_70_port, 
      boothmul_pipelined_i_muxes_in_7_69_port, 
      boothmul_pipelined_i_muxes_in_7_68_port, 
      boothmul_pipelined_i_muxes_in_7_67_port, 
      boothmul_pipelined_i_muxes_in_7_66_port, 
      boothmul_pipelined_i_muxes_in_7_65_port, 
      boothmul_pipelined_i_muxes_in_7_64_port, 
      boothmul_pipelined_i_muxes_in_7_63_port, 
      boothmul_pipelined_i_muxes_in_7_62_port, 
      boothmul_pipelined_i_muxes_in_6_218_port, 
      boothmul_pipelined_i_muxes_in_6_217_port, 
      boothmul_pipelined_i_muxes_in_6_216_port, 
      boothmul_pipelined_i_muxes_in_6_215_port, 
      boothmul_pipelined_i_muxes_in_6_214_port, 
      boothmul_pipelined_i_muxes_in_6_213_port, 
      boothmul_pipelined_i_muxes_in_6_212_port, 
      boothmul_pipelined_i_muxes_in_6_211_port, 
      boothmul_pipelined_i_muxes_in_6_210_port, 
      boothmul_pipelined_i_muxes_in_6_209_port, 
      boothmul_pipelined_i_muxes_in_6_208_port, 
      boothmul_pipelined_i_muxes_in_6_207_port, 
      boothmul_pipelined_i_muxes_in_6_206_port, 
      boothmul_pipelined_i_muxes_in_6_205_port, 
      boothmul_pipelined_i_muxes_in_6_204_port, 
      boothmul_pipelined_i_muxes_in_6_203_port, 
      boothmul_pipelined_i_muxes_in_6_73_port, 
      boothmul_pipelined_i_muxes_in_6_72_port, 
      boothmul_pipelined_i_muxes_in_6_71_port, 
      boothmul_pipelined_i_muxes_in_6_70_port, 
      boothmul_pipelined_i_muxes_in_6_69_port, 
      boothmul_pipelined_i_muxes_in_6_68_port, 
      boothmul_pipelined_i_muxes_in_6_67_port, 
      boothmul_pipelined_i_muxes_in_6_66_port, 
      boothmul_pipelined_i_muxes_in_6_65_port, 
      boothmul_pipelined_i_muxes_in_6_64_port, 
      boothmul_pipelined_i_muxes_in_6_63_port, 
      boothmul_pipelined_i_muxes_in_6_62_port, 
      boothmul_pipelined_i_muxes_in_6_61_port, 
      boothmul_pipelined_i_muxes_in_6_60_port, 
      boothmul_pipelined_i_muxes_in_6_59_port, 
      boothmul_pipelined_i_muxes_in_6_58_port, 
      boothmul_pipelined_i_muxes_in_5_205_port, 
      boothmul_pipelined_i_muxes_in_5_204_port, 
      boothmul_pipelined_i_muxes_in_5_203_port, 
      boothmul_pipelined_i_muxes_in_5_202_port, 
      boothmul_pipelined_i_muxes_in_5_201_port, 
      boothmul_pipelined_i_muxes_in_5_200_port, 
      boothmul_pipelined_i_muxes_in_5_199_port, 
      boothmul_pipelined_i_muxes_in_5_198_port, 
      boothmul_pipelined_i_muxes_in_5_197_port, 
      boothmul_pipelined_i_muxes_in_5_196_port, 
      boothmul_pipelined_i_muxes_in_5_195_port, 
      boothmul_pipelined_i_muxes_in_5_194_port, 
      boothmul_pipelined_i_muxes_in_5_193_port, 
      boothmul_pipelined_i_muxes_in_5_192_port, 
      boothmul_pipelined_i_muxes_in_5_191_port, 
      boothmul_pipelined_i_muxes_in_5_190_port, 
      boothmul_pipelined_i_muxes_in_5_189_port, 
      boothmul_pipelined_i_muxes_in_5_68_port, 
      boothmul_pipelined_i_muxes_in_5_67_port, 
      boothmul_pipelined_i_muxes_in_5_66_port, 
      boothmul_pipelined_i_muxes_in_5_65_port, 
      boothmul_pipelined_i_muxes_in_5_64_port, 
      boothmul_pipelined_i_muxes_in_5_63_port, 
      boothmul_pipelined_i_muxes_in_5_62_port, 
      boothmul_pipelined_i_muxes_in_5_61_port, 
      boothmul_pipelined_i_muxes_in_5_60_port, 
      boothmul_pipelined_i_muxes_in_5_59_port, 
      boothmul_pipelined_i_muxes_in_5_58_port, 
      boothmul_pipelined_i_muxes_in_5_57_port, 
      boothmul_pipelined_i_muxes_in_5_56_port, 
      boothmul_pipelined_i_muxes_in_5_55_port, 
      boothmul_pipelined_i_muxes_in_5_54_port, 
      boothmul_pipelined_i_muxes_in_4_190_port, 
      boothmul_pipelined_i_muxes_in_4_189_port, 
      boothmul_pipelined_i_muxes_in_4_188_port, 
      boothmul_pipelined_i_muxes_in_4_187_port, 
      boothmul_pipelined_i_muxes_in_4_186_port, 
      boothmul_pipelined_i_muxes_in_4_185_port, 
      boothmul_pipelined_i_muxes_in_4_184_port, 
      boothmul_pipelined_i_muxes_in_4_183_port, 
      boothmul_pipelined_i_muxes_in_4_182_port, 
      boothmul_pipelined_i_muxes_in_4_181_port, 
      boothmul_pipelined_i_muxes_in_4_180_port, 
      boothmul_pipelined_i_muxes_in_4_179_port, 
      boothmul_pipelined_i_muxes_in_4_178_port, 
      boothmul_pipelined_i_muxes_in_4_177_port, 
      boothmul_pipelined_i_muxes_in_4_176_port, 
      boothmul_pipelined_i_muxes_in_4_175_port, 
      boothmul_pipelined_i_muxes_in_4_65_port, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_58_port, 
      boothmul_pipelined_i_muxes_in_4_57_port, 
      boothmul_pipelined_i_muxes_in_4_56_port, 
      boothmul_pipelined_i_muxes_in_4_55_port, 
      boothmul_pipelined_i_muxes_in_4_54_port, 
      boothmul_pipelined_i_muxes_in_4_53_port, 
      boothmul_pipelined_i_muxes_in_4_52_port, 
      boothmul_pipelined_i_muxes_in_4_51_port, 
      boothmul_pipelined_i_muxes_in_4_50_port, 
      boothmul_pipelined_i_muxes_in_3_177_port, 
      boothmul_pipelined_i_muxes_in_3_176_port, 
      boothmul_pipelined_i_muxes_in_3_175_port, 
      boothmul_pipelined_i_muxes_in_3_174_port, 
      boothmul_pipelined_i_muxes_in_3_173_port, 
      boothmul_pipelined_i_muxes_in_3_172_port, 
      boothmul_pipelined_i_muxes_in_3_171_port, 
      boothmul_pipelined_i_muxes_in_3_170_port, 
      boothmul_pipelined_i_muxes_in_3_169_port, 
      boothmul_pipelined_i_muxes_in_3_168_port, 
      boothmul_pipelined_i_muxes_in_3_167_port, 
      boothmul_pipelined_i_muxes_in_3_166_port, 
      boothmul_pipelined_i_muxes_in_3_165_port, 
      boothmul_pipelined_i_muxes_in_3_164_port, 
      boothmul_pipelined_i_muxes_in_3_163_port, 
      boothmul_pipelined_i_muxes_in_3_162_port, 
      boothmul_pipelined_i_muxes_in_3_161_port, 
      boothmul_pipelined_i_muxes_in_3_60_port, 
      boothmul_pipelined_i_muxes_in_3_59_port, 
      boothmul_pipelined_i_muxes_in_3_58_port, 
      boothmul_pipelined_i_muxes_in_3_57_port, 
      boothmul_pipelined_i_muxes_in_3_56_port, 
      boothmul_pipelined_i_muxes_in_3_55_port, 
      boothmul_pipelined_i_muxes_in_3_54_port, 
      boothmul_pipelined_i_muxes_in_3_53_port, 
      boothmul_pipelined_i_muxes_in_3_52_port, 
      boothmul_pipelined_i_muxes_in_3_51_port, 
      boothmul_pipelined_i_muxes_in_3_50_port, 
      boothmul_pipelined_i_muxes_in_3_49_port, 
      boothmul_pipelined_i_muxes_in_3_48_port, 
      boothmul_pipelined_i_muxes_in_3_47_port, 
      boothmul_pipelined_i_muxes_in_3_46_port, 
      boothmul_pipelined_i_sum_out_6_0_port, 
      boothmul_pipelined_i_sum_out_6_1_port, 
      boothmul_pipelined_i_sum_out_6_2_port, 
      boothmul_pipelined_i_sum_out_6_3_port, 
      boothmul_pipelined_i_sum_out_6_4_port, 
      boothmul_pipelined_i_sum_out_6_5_port, 
      boothmul_pipelined_i_sum_out_6_6_port, 
      boothmul_pipelined_i_sum_out_6_7_port, 
      boothmul_pipelined_i_sum_out_6_8_port, 
      boothmul_pipelined_i_sum_out_6_9_port, 
      boothmul_pipelined_i_sum_out_6_10_port, 
      boothmul_pipelined_i_sum_out_6_11_port, 
      boothmul_pipelined_i_sum_out_6_13_port, 
      boothmul_pipelined_i_sum_out_6_14_port, 
      boothmul_pipelined_i_sum_out_6_15_port, 
      boothmul_pipelined_i_sum_out_6_16_port, 
      boothmul_pipelined_i_sum_out_6_17_port, 
      boothmul_pipelined_i_sum_out_6_18_port, 
      boothmul_pipelined_i_sum_out_6_19_port, 
      boothmul_pipelined_i_sum_out_6_20_port, 
      boothmul_pipelined_i_sum_out_6_21_port, 
      boothmul_pipelined_i_sum_out_6_22_port, 
      boothmul_pipelined_i_sum_out_6_23_port, 
      boothmul_pipelined_i_sum_out_6_24_port, 
      boothmul_pipelined_i_sum_out_6_25_port, 
      boothmul_pipelined_i_sum_out_6_26_port, 
      boothmul_pipelined_i_sum_out_6_27_port, 
      boothmul_pipelined_i_sum_out_6_28_port, 
      boothmul_pipelined_i_sum_out_5_0_port, 
      boothmul_pipelined_i_sum_out_5_1_port, 
      boothmul_pipelined_i_sum_out_5_2_port, 
      boothmul_pipelined_i_sum_out_5_3_port, 
      boothmul_pipelined_i_sum_out_5_4_port, 
      boothmul_pipelined_i_sum_out_5_5_port, 
      boothmul_pipelined_i_sum_out_5_6_port, 
      boothmul_pipelined_i_sum_out_5_7_port, 
      boothmul_pipelined_i_sum_out_5_8_port, 
      boothmul_pipelined_i_sum_out_5_9_port, 
      boothmul_pipelined_i_sum_out_5_11_port, 
      boothmul_pipelined_i_sum_out_5_12_port, 
      boothmul_pipelined_i_sum_out_5_13_port, 
      boothmul_pipelined_i_sum_out_5_14_port, 
      boothmul_pipelined_i_sum_out_5_15_port, 
      boothmul_pipelined_i_sum_out_5_16_port, 
      boothmul_pipelined_i_sum_out_5_17_port, 
      boothmul_pipelined_i_sum_out_5_18_port, 
      boothmul_pipelined_i_sum_out_5_19_port, 
      boothmul_pipelined_i_sum_out_5_20_port, 
      boothmul_pipelined_i_sum_out_5_21_port, 
      boothmul_pipelined_i_sum_out_5_22_port, 
      boothmul_pipelined_i_sum_out_5_23_port, 
      boothmul_pipelined_i_sum_out_5_24_port, 
      boothmul_pipelined_i_sum_out_5_25_port, 
      boothmul_pipelined_i_sum_out_5_26_port, 
      boothmul_pipelined_i_sum_out_4_0_port, 
      boothmul_pipelined_i_sum_out_4_1_port, 
      boothmul_pipelined_i_sum_out_4_2_port, 
      boothmul_pipelined_i_sum_out_4_3_port, 
      boothmul_pipelined_i_sum_out_4_4_port, 
      boothmul_pipelined_i_sum_out_4_5_port, 
      boothmul_pipelined_i_sum_out_4_6_port, 
      boothmul_pipelined_i_sum_out_4_7_port, 
      boothmul_pipelined_i_sum_out_4_9_port, 
      boothmul_pipelined_i_sum_out_4_10_port, 
      boothmul_pipelined_i_sum_out_4_11_port, 
      boothmul_pipelined_i_sum_out_4_12_port, 
      boothmul_pipelined_i_sum_out_4_13_port, 
      boothmul_pipelined_i_sum_out_4_14_port, 
      boothmul_pipelined_i_sum_out_4_15_port, 
      boothmul_pipelined_i_sum_out_4_16_port, 
      boothmul_pipelined_i_sum_out_4_17_port, 
      boothmul_pipelined_i_sum_out_4_18_port, 
      boothmul_pipelined_i_sum_out_4_19_port, 
      boothmul_pipelined_i_sum_out_4_20_port, 
      boothmul_pipelined_i_sum_out_4_21_port, 
      boothmul_pipelined_i_sum_out_4_22_port, 
      boothmul_pipelined_i_sum_out_4_23_port, 
      boothmul_pipelined_i_sum_out_4_24_port, 
      boothmul_pipelined_i_sum_out_3_0_port, 
      boothmul_pipelined_i_sum_out_3_1_port, 
      boothmul_pipelined_i_sum_out_3_2_port, 
      boothmul_pipelined_i_sum_out_3_3_port, 
      boothmul_pipelined_i_sum_out_3_4_port, 
      boothmul_pipelined_i_sum_out_3_5_port, 
      boothmul_pipelined_i_sum_out_3_7_port, 
      boothmul_pipelined_i_sum_out_3_8_port, 
      boothmul_pipelined_i_sum_out_3_9_port, 
      boothmul_pipelined_i_sum_out_3_10_port, 
      boothmul_pipelined_i_sum_out_3_11_port, 
      boothmul_pipelined_i_sum_out_3_12_port, 
      boothmul_pipelined_i_sum_out_3_13_port, 
      boothmul_pipelined_i_sum_out_3_14_port, 
      boothmul_pipelined_i_sum_out_3_15_port, 
      boothmul_pipelined_i_sum_out_3_16_port, 
      boothmul_pipelined_i_sum_out_3_17_port, 
      boothmul_pipelined_i_sum_out_3_18_port, 
      boothmul_pipelined_i_sum_out_3_19_port, 
      boothmul_pipelined_i_sum_out_3_20_port, 
      boothmul_pipelined_i_sum_out_3_21_port, 
      boothmul_pipelined_i_sum_out_3_22_port, 
      boothmul_pipelined_i_sum_out_2_0_port, 
      boothmul_pipelined_i_sum_out_2_1_port, 
      boothmul_pipelined_i_sum_out_2_2_port, 
      boothmul_pipelined_i_sum_out_2_3_port, 
      boothmul_pipelined_i_sum_out_2_5_port, 
      boothmul_pipelined_i_sum_out_2_6_port, 
      boothmul_pipelined_i_sum_out_2_7_port, 
      boothmul_pipelined_i_sum_out_2_8_port, 
      boothmul_pipelined_i_sum_out_2_9_port, 
      boothmul_pipelined_i_sum_out_2_10_port, 
      boothmul_pipelined_i_sum_out_2_11_port, 
      boothmul_pipelined_i_sum_out_2_12_port, 
      boothmul_pipelined_i_sum_out_2_13_port, 
      boothmul_pipelined_i_sum_out_2_14_port, 
      boothmul_pipelined_i_sum_out_2_15_port, 
      boothmul_pipelined_i_sum_out_2_16_port, 
      boothmul_pipelined_i_sum_out_2_17_port, 
      boothmul_pipelined_i_sum_out_2_18_port, 
      boothmul_pipelined_i_sum_out_2_19_port, 
      boothmul_pipelined_i_sum_out_2_20_port, 
      boothmul_pipelined_i_sum_out_1_0_port, 
      boothmul_pipelined_i_sum_out_1_1_port, 
      boothmul_pipelined_i_sum_out_1_3_port, 
      boothmul_pipelined_i_sum_out_1_4_port, 
      boothmul_pipelined_i_sum_out_1_5_port, 
      boothmul_pipelined_i_sum_out_1_6_port, 
      boothmul_pipelined_i_sum_out_1_7_port, 
      boothmul_pipelined_i_sum_out_1_8_port, 
      boothmul_pipelined_i_sum_out_1_9_port, 
      boothmul_pipelined_i_sum_out_1_10_port, 
      boothmul_pipelined_i_sum_out_1_11_port, 
      boothmul_pipelined_i_sum_out_1_12_port, 
      boothmul_pipelined_i_sum_out_1_13_port, 
      boothmul_pipelined_i_sum_out_1_14_port, 
      boothmul_pipelined_i_sum_out_1_15_port, 
      boothmul_pipelined_i_sum_out_1_16_port, 
      boothmul_pipelined_i_sum_out_1_17_port, 
      boothmul_pipelined_i_sum_out_1_18_port, 
      boothmul_pipelined_i_sum_B_in_7_14_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_12_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_10_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_8_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_6_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_4_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_6_28_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_5_26_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_4_24_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_3_22_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_13_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_7_15_port, 
      boothmul_pipelined_i_multiplicand_pip_6_11_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_6_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_15_port, 
      boothmul_pipelined_i_multiplicand_pip_5_9_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_5_12_port, 
      boothmul_pipelined_i_multiplicand_pip_5_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_14_port, 
      boothmul_pipelined_i_multiplicand_pip_5_15_port, 
      boothmul_pipelined_i_multiplicand_pip_4_7_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_4_10_port, 
      boothmul_pipelined_i_multiplicand_pip_4_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_12_port, 
      boothmul_pipelined_i_multiplicand_pip_4_13_port, 
      boothmul_pipelined_i_multiplicand_pip_4_14_port, 
      boothmul_pipelined_i_multiplicand_pip_4_15_port, 
      boothmul_pipelined_i_multiplicand_pip_3_5_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_3_8_port, 
      boothmul_pipelined_i_multiplicand_pip_3_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_10_port, 
      boothmul_pipelined_i_multiplicand_pip_3_11_port, 
      boothmul_pipelined_i_multiplicand_pip_3_12_port, 
      boothmul_pipelined_i_multiplicand_pip_3_13_port, 
      boothmul_pipelined_i_multiplicand_pip_3_14_port, 
      boothmul_pipelined_i_multiplicand_pip_3_15_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_multiplicand_pip_2_6_port, 
      boothmul_pipelined_i_multiplicand_pip_2_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_8_port, 
      boothmul_pipelined_i_multiplicand_pip_2_9_port, 
      boothmul_pipelined_i_multiplicand_pip_2_10_port, 
      boothmul_pipelined_i_multiplicand_pip_2_11_port, 
      boothmul_pipelined_i_multiplicand_pip_2_12_port, 
      boothmul_pipelined_i_multiplicand_pip_2_13_port, 
      boothmul_pipelined_i_multiplicand_pip_2_14_port, 
      boothmul_pipelined_i_multiplicand_pip_2_15_port, 
      boothmul_pipelined_i_muxes_in_0_119_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n1035, 
      n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, 
      n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, 
      n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, 
      n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, 
      n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, 
      n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
      n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
      n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, 
      n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, 
      n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, 
      n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, 
      n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, 
      n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, 
      n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, 
      n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
      n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, 
      n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
      n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, 
      n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, 
      n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, 
      n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, 
      n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, 
      n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
      n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
      n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
      n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, 
      n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, 
      n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
      n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, 
      n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
      n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, 
      n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, 
      n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, 
      n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, 
      n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, 
      n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
      n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
      n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, 
      n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
      n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, 
      n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, 
      n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, 
      n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, 
      n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, 
      n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, 
      n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
      n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, 
      n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, 
      n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, 
      n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, 
      n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, 
      n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, 
      n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
      n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
      n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, 
      n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, 
      n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, 
      n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, 
      n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, 
      n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, 
      n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, 
      n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, 
      n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
      n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, 
      n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, 
      n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, 
      n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, 
      n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, 
      n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
      n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, 
      n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
      n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
      n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, 
      n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, 
      n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, 
      n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
      n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, 
      n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, 
      n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, 
      n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, 
      n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, 
      n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, 
      n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, 
      n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, 
      n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, 
      n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, 
      n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, 
      n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, 
      n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, 
      n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, 
      n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, 
      n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, 
      n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, 
      n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, 
      n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, 
      n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, 
      n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, 
      n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, 
      n2516, n2517_port, n2518_port, n2519_port, n2520_port, n2521_port, 
      n2522_port, n2523_port, n2524_port, n2525_port, n2526_port, n2527_port, 
      n2528_port, n2529_port, n2530_port, n2531_port, n2532_port, n2533_port, 
      n2534_port, n2535_port, n2536_port, n2537_port, n2538_port, n2539_port, 
      n2540_port, n2541_port, n2542_port, n2543_port, n2544_port, n2545_port, 
      n2546_port, n2547_port, n2548_port, n2549, n2550, n2551, n2552, n2553, 
      n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, 
      n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
      n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, 
      n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
      n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, 
      n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, 
      n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
      n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
      n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, 
      n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, 
      n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, 
      n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, 
      n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, 
      n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, 
      n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, 
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
      n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
      n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
      n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
      n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
      n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
      n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
      n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, 
      n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, 
      n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
      n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
      n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, 
      n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
      n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
      n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
      n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
      n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
      n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
      n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
      n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
      n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356 : 
      std_logic;

begin
   
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n3099, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n3099, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n3099, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n3100, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n3100, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n3100, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n3099, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n3100, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n3100, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n3099, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n3100, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n3099, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n3100, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n3099, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n3099, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n3099, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n3100, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n3100, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n3100, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n3100, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n3100, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n3100, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n3100, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n3100, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n3100, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n3100, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n3100, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n3100, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n3099, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n3100, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n3099, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => n3098, GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => n3097, GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => n3096, GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => DATA1(3), GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, CK 
                           => clk, RN => n1042, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, QN 
                           => n3081);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, CK 
                           => clk, RN => n1037, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, QN 
                           => n_1004);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => n1039, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, QN 
                           => n_1005);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, CK 
                           => clk, RN => n1048, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, QN 
                           => n_1006);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, CK 
                           => clk, RN => n1047, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, QN 
                           => n_1007);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, CK 
                           => clk, RN => n1046, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, QN 
                           => n3080);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, CK 
                           => clk, RN => n1045, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, QN 
                           => n_1008);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, QN 
                           => n_1009);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, CK 
                           => clk, RN => n1041, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, QN 
                           => n_1010);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, CK 
                           => clk, RN => n1041, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, QN 
                           => n_1011);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, CK 
                           => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, QN 
                           => n_1012);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, CK 
                           => clk, RN => n1039, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, QN 
                           => n_1013);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, CK 
                           => clk, RN => n1048, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, QN 
                           => n3079);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, CK 
                           => clk, RN => n1047, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, QN 
                           => n_1014);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => n1046, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, QN 
                           => n_1015);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, CK 
                           => clk, RN => n1045, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, QN 
                           => n_1016);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, CK 
                           => clk, RN => n1038, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, QN 
                           => n_1017);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, CK 
                           => clk, RN => n1049, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, QN 
                           => n_1018);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, CK 
                           => clk, RN => n1036, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, QN 
                           => n_1019);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, CK 
                           => clk, RN => n1037, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, QN 
                           => n_1020);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, CK 
                           => clk, RN => n1039, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, QN 
                           => n_1021);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, CK 
                           => clk, RN => n1039, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, QN 
                           => n3078);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, CK 
                           => clk, RN => n1039, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, QN 
                           => n_1022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, QN 
                           => n_1023);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, CK 
                           => clk, RN => n1038, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, QN 
                           => n_1024);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, CK 
                           => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, QN 
                           => n_1025);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, CK 
                           => clk, RN => n1049, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, QN 
                           => n_1026);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, CK 
                           => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, QN 
                           => n_1027);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, CK 
                           => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, QN 
                           => n_1028);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, QN 
                           => n_1029);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, CK 
                           => clk, RN => n1044, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, QN 
                           => n_1030);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, CK 
                           => clk, RN => n1043, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, QN 
                           => n_1031);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, CK 
                           => clk, RN => n1038, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, QN 
                           => n3082);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, CK 
                           => clk, RN => n1048, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, QN 
                           => n_1032);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, CK 
                           => clk, RN => n1047, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, QN 
                           => n_1033);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_15_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, QN 
                           => n_1034);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_14_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, QN 
                           => n_1035);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_13_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, QN 
                           => n_1036);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_12_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, QN 
                           => n_1037);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_11_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, QN 
                           => n_1038);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_10_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, QN 
                           => n_1039);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_9_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, QN 
                           => n_1040);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_8_port, CK => clk, RN => n1037, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, QN 
                           => n_1041);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_7_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, QN 
                           => n_1042);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_6_port, CK => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, QN 
                           => n_1043);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_5_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, QN 
                           => n3076);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_4_port, CK => clk, RN => n1038, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, QN 
                           => n_1044);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_3_port, CK => clk, RN => n1043, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, QN 
                           => n_1045);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_28_port, CK => clk
                           , RN => n1045, Q => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, QN => 
                           n_1046);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_27_port, CK => clk
                           , RN => n1049, Q => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, QN => 
                           n_1047);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_26_port, CK => clk
                           , RN => n1046, Q => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, QN => 
                           n_1048);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_25_port, CK => clk
                           , RN => n1039, Q => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, QN => 
                           n_1049);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_24_port, CK => clk
                           , RN => n1044, Q => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, QN => 
                           n_1050);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_23_port, CK => clk
                           , RN => n1048, Q => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, QN => 
                           n_1051);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_22_port, CK => clk
                           , RN => n1038, Q => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, QN => 
                           n_1052);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_21_port, CK => clk
                           , RN => n1040, Q => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, QN => 
                           n_1053);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_20_port, CK => clk
                           , RN => n1042, Q => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, QN => 
                           n_1054);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_19_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, QN => 
                           n_1055);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_18_port, CK => clk
                           , RN => n1036, Q => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, QN => 
                           n_1056);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_17_port, CK => clk
                           , RN => n1038, Q => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, QN => 
                           n_1057);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_16_port, CK => clk
                           , RN => n1044, Q => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, QN => 
                           n_1058);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_15_port, CK => clk
                           , RN => n1036, Q => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, QN => 
                           n_1059);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_14_port, CK => clk
                           , RN => n1047, Q => 
                           boothmul_pipelined_i_sum_B_in_7_14_port, QN => 
                           n_1060);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_13_port, CK => clk
                           , RN => n1043, Q => dataout_mul_13_port, QN => 
                           n_1061);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => n3095, CK => clk, RN => n1042, Q => 
                           dataout_mul_12_port, QN => n_1062);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_11_port, CK => clk
                           , RN => n1039, Q => dataout_mul_11_port, QN => 
                           n_1063);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_10_port, CK => clk
                           , RN => n1037, Q => dataout_mul_10_port, QN => 
                           n_1064);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_9_port, CK => clk, RN
                           => n1044, Q => dataout_mul_9_port, QN => n_1065);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_8_port, CK => clk, RN
                           => n1043, Q => dataout_mul_8_port, QN => n_1066);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_7_port, CK => clk, RN
                           => n1042, Q => dataout_mul_7_port, QN => n_1067);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_6_port, CK => clk, RN
                           => n1041, Q => dataout_mul_6_port, QN => n_1068);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_5_port, CK => clk, RN
                           => n1049, Q => dataout_mul_5_port, QN => n_1069);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_4_port, CK => clk, RN
                           => n1048, Q => dataout_mul_4_port, QN => n_1070);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_3_port, CK => clk, RN
                           => n1038, Q => dataout_mul_3_port, QN => n_1071);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_2_port, CK => clk, RN
                           => n1037, Q => dataout_mul_2_port, QN => n_1072);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_1_port, CK => clk, RN
                           => n1040, Q => dataout_mul_1_port, QN => n_1073);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_0_port, CK => clk, RN
                           => rst_BAR, Q => dataout_mul_0_port, QN => n_1074);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_58_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_7_62_port, QN => 
                           n_1075);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_59_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_7_63_port, QN => 
                           n_1076);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_60_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_7_64_port, QN => 
                           n_1077);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_61_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_7_65_port, QN => 
                           n_1078);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_62_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_7_66_port, QN => 
                           n_1079);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_63_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_7_67_port, QN => 
                           n_1080);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_64_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_7_68_port, QN => 
                           n_1081);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_65_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_7_69_port, QN => 
                           n_1082);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_66_port, CK => 
                           clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_7_70_port, QN => 
                           n_1083);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_67_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_7_71_port, QN => 
                           n_1084);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_68_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_7_72_port, QN => 
                           n_1085);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_69_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_7_73_port, QN => 
                           n_1086);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_178_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_70_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_7_74_port, QN => 
                           n_1087);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_177_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_71_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_7_75_port, QN => 
                           n_1088);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_176_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_72_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_7_76_port, QN => 
                           n_1089);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_175_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_7_77_port, QN => 
                           n_1090);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_203_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_7_217_port, QN => 
                           n_1091);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_204_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_7_218_port, QN => 
                           n_1092);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_205_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_7_219_port, QN => 
                           n_1093);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_42_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_206_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_7_220_port, QN => 
                           n_1094);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_41_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_207_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_221_port, QN => 
                           n_1095);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_40_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_208_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_7_222_port, QN => 
                           n_1096);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_39_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_209_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_7_223_port, QN => 
                           n_1097);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_38_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_210_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_7_224_port, QN => 
                           n_1098);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_37_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_211_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_7_225_port, QN => 
                           n_1099);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_36_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_212_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_7_226_port, QN => 
                           n_1100);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_35_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_213_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_7_227_port, QN => 
                           n_1101);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_34_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_214_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_7_228_port, QN => 
                           n_1102);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_33_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_215_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_7_229_port, QN => 
                           n_1103);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_216_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_7_230_port, QN => 
                           n_1104);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_217_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_7_231_port, QN => 
                           n_1105);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_218_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_7_232_port, QN => 
                           n_1106);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_7_233_port, QN => 
                           n_1107);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_26_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, QN => 
                           n_1108);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_25_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, QN => 
                           n_1109);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_24_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, QN => 
                           n_1110);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_23_port, CK => clk
                           , RN => n1038, Q => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, QN => 
                           n_1111);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_22_port, CK => clk
                           , RN => n1049, Q => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, QN => 
                           n_1112);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_21_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, QN => 
                           n_1113);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_20_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, QN => 
                           n_1114);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_19_port, CK => clk
                           , RN => n1043, Q => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, QN => 
                           n_1115);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_18_port, CK => clk
                           , RN => n1042, Q => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, QN => 
                           n_1116);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_17_port, CK => clk
                           , RN => n1042, Q => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, QN => 
                           n_1117);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_16_port, CK => clk
                           , RN => n1045, Q => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, QN => 
                           n_1118);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_15_port, CK => clk
                           , RN => n1040, Q => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, QN => 
                           n_1119);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_14_port, CK => clk
                           , RN => n1039, Q => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, QN => 
                           n_1120);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_13_port, CK => clk
                           , RN => n1042, Q => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, QN => 
                           n_1121);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_12_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_B_in_6_12_port, QN => 
                           n_1122);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_11_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_out_6_11_port, QN => n_1123
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => n3094, CK => clk, RN => n1039, Q => 
                           boothmul_pipelined_i_sum_out_6_10_port, QN => n_1124
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_9_port, CK => clk, RN
                           => n1048, Q => boothmul_pipelined_i_sum_out_6_9_port
                           , QN => n_1125);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_8_port, CK => clk, RN
                           => n1048, Q => boothmul_pipelined_i_sum_out_6_8_port
                           , QN => n_1126);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_7_port, CK => clk, RN
                           => n1038, Q => boothmul_pipelined_i_sum_out_6_7_port
                           , QN => n_1127);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_6_port, CK => clk, RN
                           => n1040, Q => boothmul_pipelined_i_sum_out_6_6_port
                           , QN => n_1128);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_5_port, CK => clk, RN
                           => n1046, Q => boothmul_pipelined_i_sum_out_6_5_port
                           , QN => n_1129);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_4_port, CK => clk, RN
                           => n1046, Q => boothmul_pipelined_i_sum_out_6_4_port
                           , QN => n_1130);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_3_port, CK => clk, RN
                           => n1047, Q => boothmul_pipelined_i_sum_out_6_3_port
                           , QN => n_1131);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_2_port, CK => clk, RN
                           => n1046, Q => boothmul_pipelined_i_sum_out_6_2_port
                           , QN => n_1132);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_1_port, CK => clk, RN
                           => n1042, Q => boothmul_pipelined_i_sum_out_6_1_port
                           , QN => n_1133);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_0_port, CK => clk, RN
                           => n1044, Q => boothmul_pipelined_i_sum_out_6_0_port
                           , QN => n_1134);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_54_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_6_58_port, QN => 
                           n_1135);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_55_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_6_59_port, QN => 
                           n_1136);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_56_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_6_60_port, QN => 
                           n_1137);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_57_port, CK => 
                           clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_6_61_port, QN => 
                           n_1138);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_58_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_6_62_port, QN => 
                           n_1139);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_59_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_6_63_port, QN => 
                           n_1140);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_60_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_6_64_port, QN => 
                           n_1141);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_61_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_6_65_port, QN => 
                           n_1142);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_62_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_6_66_port, QN => 
                           n_1143);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_63_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_6_67_port, QN => 
                           n_1144);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_64_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_6_68_port, QN => 
                           n_1145);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_65_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_6_69_port, QN => 
                           n_1146);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_66_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_6_70_port, QN => 
                           n_1147);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_67_port, CK => 
                           clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_6_71_port, QN => 
                           n_1148);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_68_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_6_72_port, QN => 
                           n_1149);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_205_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_6_73_port, QN => 
                           n_1150);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_189_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_6_203_port, QN => 
                           n_1151);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_190_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_6_204_port, QN => 
                           n_1152);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_191_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_6_205_port, QN => 
                           n_1153);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_56_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_192_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_6_206_port, QN => 
                           n_1154);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_55_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_193_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_6_207_port, QN => 
                           n_1155);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_54_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_194_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_6_208_port, QN => 
                           n_1156);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_53_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_195_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_6_209_port, QN => 
                           n_1157);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_52_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_196_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_6_210_port, QN => 
                           n_1158);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_51_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_197_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_6_211_port, QN => 
                           n_1159);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_50_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_198_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_6_212_port, QN => 
                           n_1160);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_49_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_199_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_6_213_port, QN => 
                           n_1161);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_48_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_200_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_6_214_port, QN => 
                           n_1162);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_47_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_201_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_6_215_port, QN => 
                           n_1163);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_46_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_202_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_6_216_port, QN => 
                           n_1164);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_203_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_6_217_port, QN => 
                           n_1165);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_204_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_6_218_port, QN => 
                           n_1166);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_24_port, CK => clk
                           , RN => n1047, Q => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, QN => 
                           n_1167);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_23_port, CK => clk
                           , RN => n1036, Q => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, QN => 
                           n_1168);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_22_port, CK => clk
                           , RN => n1037, Q => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, QN => 
                           n_1169);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_21_port, CK => clk
                           , RN => n1045, Q => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, QN => 
                           n_1170);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_20_port, CK => clk
                           , RN => n1037, Q => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, QN => 
                           n_1171);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_19_port, CK => clk
                           , RN => n1042, Q => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, QN => 
                           n_1172);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_18_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, QN => 
                           n_1173);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_17_port, CK => clk
                           , RN => n1038, Q => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, QN => 
                           n_1174);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_16_port, CK => clk
                           , RN => n1045, Q => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, QN => 
                           n_1175);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_15_port, CK => clk
                           , RN => n1049, Q => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, QN => 
                           n_1176);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_14_port, CK => clk
                           , RN => n1039, Q => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, QN => 
                           n_1177);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_13_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, QN => 
                           n_1178);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_12_port, CK => clk
                           , RN => n1048, Q => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, QN => 
                           n_1179);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_11_port, CK => clk
                           , RN => n1048, Q => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, QN => 
                           n_1180);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_10_port, CK => clk
                           , RN => n1048, Q => 
                           boothmul_pipelined_i_sum_B_in_5_10_port, QN => 
                           n_1181);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_9_port, CK => clk, RN
                           => n1047, Q => boothmul_pipelined_i_sum_out_5_9_port
                           , QN => n_1182);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           n3093, CK => clk, RN => n1046, Q => 
                           boothmul_pipelined_i_sum_out_5_8_port, QN => n_1183)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_7_port, CK => clk, RN
                           => n1049, Q => boothmul_pipelined_i_sum_out_5_7_port
                           , QN => n_1184);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_6_port, CK => clk, RN
                           => n1038, Q => boothmul_pipelined_i_sum_out_5_6_port
                           , QN => n_1185);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_5_port, CK => clk, RN
                           => n1046, Q => boothmul_pipelined_i_sum_out_5_5_port
                           , QN => n_1186);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_4_port, CK => clk, RN
                           => n1047, Q => boothmul_pipelined_i_sum_out_5_4_port
                           , QN => n_1187);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_3_port, CK => clk, RN
                           => n1037, Q => boothmul_pipelined_i_sum_out_5_3_port
                           , QN => n_1188);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_2_port, CK => clk, RN
                           => n1037, Q => boothmul_pipelined_i_sum_out_5_2_port
                           , QN => n_1189);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_1_port, CK => clk, RN
                           => n1041, Q => boothmul_pipelined_i_sum_out_5_1_port
                           , QN => n_1190);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_0_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_0_port, QN => n_1191)
                           ;
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_50_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_5_54_port, QN => 
                           n_1192);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_51_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_5_55_port, QN => 
                           n_1193);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_52_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_5_56_port, QN => 
                           n_1194);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_53_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_5_57_port, QN => 
                           n_1195);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_54_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_5_58_port, QN => 
                           n_1196);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_55_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_5_59_port, QN => 
                           n_1197);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_56_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_5_60_port, QN => 
                           n_1198);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_57_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_61_port, QN => 
                           n_1199);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_58_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_5_62_port, QN => 
                           n_1200);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_59_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_5_63_port, QN => 
                           n_1201);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_60_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_5_64_port, QN => 
                           n_1202);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_61_port, CK => 
                           clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_5_65_port, QN => 
                           n_1203);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_62_port, CK => 
                           clk, RN => n1038, Q => 
                           boothmul_pipelined_i_muxes_in_5_66_port, QN => 
                           n_1204);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_63_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_5_67_port, QN => 
                           n_1205);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_64_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_5_68_port, QN => 
                           n_1206);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_175_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_5_189_port, QN => 
                           n_1207);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_176_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_5_190_port, QN => 
                           n_1208);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_177_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_5_191_port, QN => 
                           n_1209);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_178_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_5_192_port, QN => 
                           n_1210);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_179_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_193_port, QN => 
                           n_1211);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_180_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_194_port, QN => 
                           n_1212);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_181_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_195_port, QN => 
                           n_1213);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_182_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_196_port, QN => 
                           n_1214);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_183_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_197_port, QN => 
                           n_1215);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_184_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_198_port, QN => 
                           n_1216);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_185_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_199_port, QN => 
                           n_1217);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_186_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_200_port, QN => 
                           n_1218);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_187_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_201_port, QN => 
                           n_1219);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_188_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_5_202_port, QN => 
                           n_1220);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_189_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_5_203_port, QN => 
                           n_1221);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_190_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_5_204_port, QN => 
                           n_1222);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_65_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_5_205_port, QN => 
                           n_1223);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_22_port, CK => clk
                           , RN => n1047, Q => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, QN => 
                           n_1224);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_21_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, QN => 
                           n_1225);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_20_port, CK => clk
                           , RN => n1035, Q => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, QN => 
                           n_1226);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_19_port, CK => clk
                           , RN => n1045, Q => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, QN => 
                           n_1227);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_18_port, CK => clk
                           , RN => n1039, Q => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, QN => 
                           n_1228);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_17_port, CK => clk
                           , RN => n1035, Q => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, QN => 
                           n_1229);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_16_port, CK => clk
                           , RN => n1049, Q => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, QN => 
                           n_1230);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_15_port, CK => clk
                           , RN => n1048, Q => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, QN => 
                           n_1231);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_14_port, CK => clk
                           , RN => n1039, Q => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, QN => 
                           n_1232);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_13_port, CK => clk
                           , RN => n1039, Q => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, QN => 
                           n_1233);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_12_port, CK => clk
                           , RN => n1046, Q => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, QN => 
                           n_1234);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, QN => 
                           n_1235);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_10_port, CK => clk
                           , RN => n1041, Q => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, QN => 
                           n_1236);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_9_port, CK => clk, RN
                           => n1049, Q => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, QN => n_1237
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_8_port, CK => clk, RN
                           => n1042, Q => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, QN => n_1238
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_7_port, CK => clk, RN
                           => n1047, Q => boothmul_pipelined_i_sum_out_4_7_port
                           , QN => n_1239);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           n3092, CK => clk, RN => n1043, Q => 
                           boothmul_pipelined_i_sum_out_4_6_port, QN => n_1240)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_5_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_5_port, QN => n_1241)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_4_port, CK => clk, RN
                           => n1047, Q => boothmul_pipelined_i_sum_out_4_4_port
                           , QN => n_1242);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_3_port, CK => clk, RN
                           => n1046, Q => boothmul_pipelined_i_sum_out_4_3_port
                           , QN => n_1243);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_2_port, CK => clk, RN
                           => n1049, Q => boothmul_pipelined_i_sum_out_4_2_port
                           , QN => n_1244);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_1_port, CK => clk, RN
                           => n1049, Q => boothmul_pipelined_i_sum_out_4_1_port
                           , QN => n_1245);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_0_port, CK => clk, RN
                           => n1038, Q => boothmul_pipelined_i_sum_out_4_0_port
                           , QN => n_1246);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_46_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_4_50_port, QN => 
                           n_1247);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_47_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_4_51_port, QN => 
                           n_1248);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_48_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_4_52_port, QN => 
                           n_1249);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_49_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_4_53_port, QN => 
                           n_1250);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_50_port, CK => 
                           clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_4_54_port, QN => 
                           n_1251);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_51_port, CK => 
                           clk, RN => n1038, Q => 
                           boothmul_pipelined_i_muxes_in_4_55_port, QN => 
                           n_1252);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_52_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_4_56_port, QN => 
                           n_1253);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_53_port, CK => 
                           clk, RN => n1038, Q => 
                           boothmul_pipelined_i_muxes_in_4_57_port, QN => 
                           n_1254);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_54_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_4_58_port, QN => 
                           n_1255);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_55_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port, QN => 
                           n_1256);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_56_port, CK => 
                           clk, RN => n1047, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port, QN => 
                           n_1257);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_57_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port, QN => 
                           n_1258);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_58_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port, QN => 
                           n_1259);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_59_port, CK => 
                           clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port, QN => 
                           n_1260);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_60_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port, QN => 
                           n_1261);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_177_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_4_65_port, QN => 
                           n_1262);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_161_port, CK => 
                           clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_4_175_port, QN => 
                           n_1263);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_162_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_4_176_port, QN => 
                           n_1264);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_163_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_4_177_port, QN => 
                           n_1265);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_164_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_4_178_port, QN => 
                           n_1266);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_165_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_4_179_port, QN => 
                           n_1267);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_166_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_4_180_port, QN => 
                           n_1268);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_167_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_4_181_port, QN => 
                           n_1269);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_168_port, CK => 
                           clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_4_182_port, QN => 
                           n_1270);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_169_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_4_183_port, QN => 
                           n_1271);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_170_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_4_184_port, QN => 
                           n_1272);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_171_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_4_185_port, QN => 
                           n_1273);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_172_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_4_186_port, QN => 
                           n_1274);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_173_port, CK => 
                           clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_4_187_port, QN => 
                           n_1275);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_174_port, CK => 
                           clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_4_188_port, QN => 
                           n_1276);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_175_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_4_189_port, QN => 
                           n_1277);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_176_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_4_190_port, QN => 
                           n_1278);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_20_port, CK => clk
                           , RN => n1035, Q => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, QN => 
                           n_1279);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_19_port, CK => clk
                           , RN => n1046, Q => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, QN => 
                           n_1280);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_18_port, CK => clk
                           , RN => n1036, Q => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, QN => 
                           n_1281);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_17_port, CK => clk
                           , RN => n1040, Q => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, QN => 
                           n_1282);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_16_port, CK => clk
                           , RN => n1036, Q => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, QN => 
                           n_1283);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_15_port, CK => clk
                           , RN => n1036, Q => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, QN => 
                           n_1284);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_14_port, CK => clk
                           , RN => n1035, Q => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, QN => 
                           n_1285);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_13_port, CK => clk
                           , RN => n1047, Q => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, QN => 
                           n_1286);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_12_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, QN => 
                           n_1287);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_11_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, QN => 
                           n_1288);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_10_port, CK => clk
                           , RN => n1044, Q => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, QN => 
                           n_1289);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_9_port, CK => clk, RN
                           => n1045, Q => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, QN => n_1290
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_8_port, CK => clk, RN
                           => n1039, Q => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, QN => n_1291
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_7_port, CK => clk, RN
                           => n1048, Q => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, QN => n_1292
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_6_port, CK => clk, RN
                           => n1048, Q => 
                           boothmul_pipelined_i_sum_B_in_3_6_port, QN => n_1293
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_5_port, CK => clk, RN
                           => n1036, Q => boothmul_pipelined_i_sum_out_3_5_port
                           , QN => n_1294);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           n3091, CK => clk, RN => n1037, Q => 
                           boothmul_pipelined_i_sum_out_3_4_port, QN => n_1295)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_3_port, CK => clk, RN
                           => n1045, Q => boothmul_pipelined_i_sum_out_3_3_port
                           , QN => n_1296);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_2_port, CK => clk, RN
                           => n1048, Q => boothmul_pipelined_i_sum_out_3_2_port
                           , QN => n_1297);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_1_port, CK => clk, RN
                           => n1048, Q => boothmul_pipelined_i_sum_out_3_1_port
                           , QN => n_1298);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_0_port, CK => clk, RN
                           => n1047, Q => boothmul_pipelined_i_sum_out_3_0_port
                           , QN => n_1299);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_3_46_port, QN => 
                           n_1300);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_3_47_port, QN => 
                           n_1301);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_3_48_port, QN => 
                           n_1302);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => rst_BAR, Q =>
                           boothmul_pipelined_i_muxes_in_3_49_port, QN => 
                           n_1303);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_3_50_port, QN => 
                           n_1304);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_3_51_port, QN => 
                           n_1305);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => n1038, Q => 
                           boothmul_pipelined_i_muxes_in_3_52_port, QN => 
                           n_1306);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_3_53_port, QN => 
                           n_1307);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => n1038, Q => 
                           boothmul_pipelined_i_muxes_in_3_54_port, QN => 
                           n_1308);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_3_55_port, QN => 
                           n_1309);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => n1035, Q => 
                           boothmul_pipelined_i_muxes_in_3_56_port, QN => 
                           n_1310);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_3_57_port, QN => 
                           n_1311);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_58_port, QN => 
                           n_1312);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => n1049, Q => 
                           boothmul_pipelined_i_muxes_in_3_59_port, QN => 
                           n_1313);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => n1038, Q => 
                           boothmul_pipelined_i_muxes_in_3_60_port, QN => 
                           n_1314);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_119_port, CK => 
                           clk, RN => n1044, Q => 
                           boothmul_pipelined_i_muxes_in_3_161_port, QN => 
                           n_1315);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => n1043, Q => 
                           boothmul_pipelined_i_muxes_in_3_162_port, QN => 
                           n_1316);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => n1042, Q => 
                           boothmul_pipelined_i_muxes_in_3_163_port, QN => 
                           n_1317);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_3_164_port, QN => 
                           n_1318);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => n1036, Q => 
                           boothmul_pipelined_i_muxes_in_3_165_port, QN => 
                           n_1319);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => n1037, Q => 
                           boothmul_pipelined_i_muxes_in_3_166_port, QN => 
                           n_1320);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => n1048, Q => 
                           boothmul_pipelined_i_muxes_in_3_167_port, QN => 
                           n_1321);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_3_168_port, QN => 
                           n_1322);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_3_169_port, QN => 
                           n_1323);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_3_170_port, QN => 
                           n_1324);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_3_171_port, QN => 
                           n_1325);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => n1040, Q => 
                           boothmul_pipelined_i_muxes_in_3_172_port, QN => 
                           n_1326);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => n1041, Q => 
                           boothmul_pipelined_i_muxes_in_3_173_port, QN => 
                           n_1327);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => n1038, Q => 
                           boothmul_pipelined_i_muxes_in_3_174_port, QN => 
                           n_1328);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => n1039, Q => 
                           boothmul_pipelined_i_muxes_in_3_175_port, QN => 
                           n_1329);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => n1046, Q => 
                           boothmul_pipelined_i_muxes_in_3_176_port, QN => 
                           n_1330);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_18_port, CK => clk
                           , RN => n1047, Q => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, QN => 
                           n_1331);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_17_port, CK => clk
                           , RN => n1043, Q => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, QN => 
                           n_1332);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_16_port, CK => clk
                           , RN => n1043, Q => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, QN => 
                           n_1333);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_15_port, CK => clk
                           , RN => n1043, Q => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, QN => 
                           n_1334);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_14_port, CK => clk
                           , RN => n1043, Q => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, QN => 
                           n_1335);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_13_port, CK => clk
                           , RN => n1043, Q => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, QN => 
                           n_1336);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_12_port, CK => clk
                           , RN => n1043, Q => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, QN => 
                           n_1337);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_11_port, CK => clk
                           , RN => n1042, Q => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, QN => 
                           n_1338);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_10_port, CK => clk
                           , RN => n1046, Q => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, QN => 
                           n_1339);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_9_port, CK => clk, RN
                           => n1036, Q => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, QN => n_1340
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_8_port, CK => clk, RN
                           => n1046, Q => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, QN => n_1341
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_7_port, CK => clk, RN
                           => n1046, Q => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, QN => n_1342
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_6_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, QN => n_1343
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_5_port, CK => clk, RN
                           => n1046, Q => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, QN => n_1344
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_4_port, CK => clk, RN
                           => n1044, Q => 
                           boothmul_pipelined_i_sum_B_in_2_4_port, QN => n_1345
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_3_port, CK => clk, RN
                           => n1037, Q => boothmul_pipelined_i_sum_out_2_3_port
                           , QN => n_1346);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           n3086, CK => clk, RN => n1037, Q => 
                           boothmul_pipelined_i_sum_out_2_2_port, QN => n_1347)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_1_port, CK => clk, RN
                           => n1038, Q => boothmul_pipelined_i_sum_out_2_1_port
                           , QN => n_1348);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_0_port, CK => clk, RN
                           => n1038, Q => boothmul_pipelined_i_sum_out_2_0_port
                           , QN => n_1349);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => n1045, Q => 
                           boothmul_pipelined_i_muxes_in_3_177_port, QN => 
                           n3077);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n3099, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3083,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => boothmul_pipelined_i_sum_out_1_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_out_1_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_1_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_1_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_1_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_1_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_1_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_1_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_1_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_1_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_1_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_1_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_1_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_1_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_1_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1350, S => 
                           boothmul_pipelined_i_sum_out_1_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CI => n3085,
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_2_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_2_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_2_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_2_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_2_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_2_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_2_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_2_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_2_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_2_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_2_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_2_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_2_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_2_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_2_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CO => n_1351, S => 
                           boothmul_pipelined_i_sum_out_2_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3084,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_3_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_3_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_3_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_3_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_3_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_3_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_3_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_3_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_3_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_3_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_3_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_3_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_3_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_3_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_3_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1352, S => 
                           boothmul_pipelined_i_sum_out_3_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CI => n3090,
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_4_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_4_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_4_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_4_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_4_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_4_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_4_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_4_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_4_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_4_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_4_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_4_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_4_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_4_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_4_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1353, S => 
                           boothmul_pipelined_i_sum_out_4_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CI => n3089
                           , CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_5_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_5_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_5_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_5_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_5_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_5_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_5_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_5_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_5_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_5_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_5_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_5_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_5_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_5_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_5_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1354, S => 
                           boothmul_pipelined_i_sum_out_5_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CI => n3088
                           , CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_6_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_6_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_6_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_6_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_6_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_6_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_6_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_6_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_6_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_6_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_6_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_6_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_6_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_out_6_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_out_6_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1355, S => 
                           boothmul_pipelined_i_sum_out_6_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CI => n3087
                           , CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_29_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1356, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   U3 : CLKBUF_X1 port map( A => n1038, Z => n1035);
   U4 : CLKBUF_X1 port map( A => n1038, Z => n1036);
   U5 : CLKBUF_X1 port map( A => n1038, Z => n1037);
   U6 : CLKBUF_X1 port map( A => rst_BAR, Z => n1038);
   U7 : CLKBUF_X1 port map( A => n1040, Z => n1039);
   U8 : CLKBUF_X1 port map( A => n1035, Z => n1040);
   U9 : CLKBUF_X1 port map( A => n1036, Z => n1041);
   U10 : CLKBUF_X1 port map( A => n1036, Z => n1042);
   U11 : CLKBUF_X1 port map( A => n1036, Z => n1043);
   U12 : CLKBUF_X1 port map( A => n1036, Z => n1044);
   U13 : CLKBUF_X1 port map( A => n1037, Z => n1045);
   U14 : CLKBUF_X1 port map( A => n1037, Z => n1046);
   U15 : CLKBUF_X1 port map( A => n1037, Z => n1047);
   U16 : CLKBUF_X1 port map( A => n1037, Z => n1048);
   U17 : CLKBUF_X1 port map( A => n1037, Z => n1049);
   U18 : AOI211_X4 port map( C1 => data2_mul_1_port, C2 => data2_mul_2_port, A 
                           => data2_mul_3_port, B => n2783, ZN => n2811);
   U19 : AOI211_X4 port map( C1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, C2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => boothmul_pipelined_i_multiplicand_pip_2_5_port, B
                           => n2823, ZN => n2852);
   U20 : NOR2_X2 port map( A1 => n1115, A2 => n1651, ZN => n2494);
   U21 : CLKBUF_X1 port map( A => n2779, Z => n2769);
   U22 : NOR2_X1 port map( A1 => FUNC(2), A2 => FUNC(0), ZN => n1093);
   U23 : INV_X1 port map( A => FUNC(1), ZN => n1919);
   U24 : AND2_X1 port map( A1 => n1093, A2 => n1919, ZN => n2744);
   U25 : INV_X1 port map( A => n2744, ZN => n3100);
   U26 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n1050);
   U27 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, A
                           => n1050, ZN => n1073);
   U28 : NOR2_X1 port map( A1 => boothmul_pipelined_i_multiplicand_pip_3_7_port
                           , A2 => n1073, ZN => n2879);
   U29 : CLKBUF_X1 port map( A => n2879, Z => n2897);
   U30 : NAND3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           A3 => n3082, ZN => n2865);
   U31 : INV_X1 port map( A => n2865, ZN => n2895);
   U32 : NOR2_X1 port map( A1 => boothmul_pipelined_i_multiplicand_pip_3_6_port
                           , A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, ZN 
                           => n1051);
   U33 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, A2 
                           => n1051, ZN => n2864);
   U34 : INV_X1 port map( A => n2864, ZN => n2894);
   U35 : NOR2_X1 port map( A1 => n3082, A2 => n1073, ZN => n2878);
   U36 : CLKBUF_X1 port map( A => n2878, Z => n2896);
   U37 : AOI22_X1 port map( A1 => n2894, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, B1 => 
                           n2896, B2 => 
                           boothmul_pipelined_i_muxes_in_3_161_port, ZN => 
                           n1052);
   U38 : INV_X1 port map( A => n1052, ZN => n1053);
   U39 : AOI221_X1 port map( B1 => boothmul_pipelined_i_muxes_in_3_46_port, B2 
                           => n2897, C1 => 
                           boothmul_pipelined_i_muxes_in_3_46_port, C2 => n2895
                           , A => n1053, ZN => n1054);
   U40 : INV_X1 port map( A => n1054, ZN => 
                           boothmul_pipelined_i_mux_out_3_22_port);
   U41 : INV_X1 port map( A => data1_mul_15_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port);
   U42 : XOR2_X1 port map( A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, B 
                           => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => boothmul_pipelined_i_muxes_in_0_119_port);
   U43 : INV_X1 port map( A => data1_mul_0_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port);
   U44 : INV_X1 port map( A => data1_mul_2_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port);
   U45 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n1055);
   U46 : OAI21_X1 port map( B1 => data2_mul_1_port, B2 => data2_mul_2_port, A 
                           => n1055, ZN => n2782);
   U47 : NOR2_X1 port map( A1 => n2782, A2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           ZN => n1078);
   U48 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n3070);
   U49 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_115_port, ZN => 
                           n3056);
   U50 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN =>
                           n2781);
   U51 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => n2781, ZN => n3069);
   U52 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n3055);
   U53 : OR2_X1 port map( A1 => n2781, A2 => data2_mul_1_port, ZN => n3075);
   U54 : OAI222_X1 port map( A1 => n3070, A2 => n3056, B1 => n3069, B2 => n3055
                           , C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, 
                           C2 => n3075, ZN => n1079);
   U55 : AND2_X1 port map( A1 => n1078, A2 => n1079, ZN => n3083);
   U56 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n1056);
   U57 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           A => n1056, ZN => n1057);
   U58 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, A2 
                           => n1057, ZN => n3011);
   U59 : CLKBUF_X1 port map( A => n3011, Z => n3005);
   U60 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, A2 
                           => n1056, ZN => n2988);
   U61 : NOR2_X1 port map( A1 => n3080, A2 => n1057, ZN => n3010);
   U62 : CLKBUF_X1 port map( A => n3010, Z => n2999);
   U63 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           A3 => n3080, ZN => n3008);
   U64 : CLKBUF_X1 port map( A => n3008, Z => n3004);
   U65 : AOI22_X1 port map( A1 => n2999, A2 => 
                           boothmul_pipelined_i_muxes_in_6_203_port, B1 => 
                           n3004, B2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, ZN => 
                           n1058);
   U66 : INV_X1 port map( A => n1058, ZN => n1059);
   U67 : AOI221_X1 port map( B1 => boothmul_pipelined_i_muxes_in_6_58_port, B2 
                           => n3005, C1 => 
                           boothmul_pipelined_i_muxes_in_6_58_port, C2 => n2988
                           , A => n1059, ZN => n1060);
   U68 : INV_X1 port map( A => n1060, ZN => 
                           boothmul_pipelined_i_mux_out_6_28_port);
   U69 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n1061);
   U70 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, A
                           => n1061, ZN => n1062);
   U71 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, A2 
                           => n1062, ZN => n2973);
   U72 : CLKBUF_X1 port map( A => n2973, Z => n2967);
   U73 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, A2 
                           => n1061, ZN => n2950);
   U74 : NOR2_X1 port map( A1 => n3079, A2 => n1062, ZN => n2972);
   U75 : CLKBUF_X1 port map( A => n2972, Z => n2961);
   U76 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           A3 => n3079, ZN => n2970);
   U77 : CLKBUF_X1 port map( A => n2970, Z => n2966);
   U78 : AOI22_X1 port map( A1 => n2961, A2 => 
                           boothmul_pipelined_i_muxes_in_5_189_port, B1 => 
                           n2966, B2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, ZN => 
                           n1063);
   U79 : INV_X1 port map( A => n1063, ZN => n1064);
   U80 : AOI221_X1 port map( B1 => boothmul_pipelined_i_muxes_in_5_54_port, B2 
                           => n2967, C1 => 
                           boothmul_pipelined_i_muxes_in_5_54_port, C2 => n2950
                           , A => n1064, ZN => n1065);
   U81 : INV_X1 port map( A => n1065, ZN => 
                           boothmul_pipelined_i_mux_out_5_26_port);
   U82 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n1066);
   U83 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, A
                           => n1066, ZN => n1067);
   U84 : NOR2_X1 port map( A1 => boothmul_pipelined_i_multiplicand_pip_4_9_port
                           , A2 => n1067, ZN => n2935);
   U85 : CLKBUF_X1 port map( A => n2935, Z => n2929);
   U86 : NOR2_X1 port map( A1 => boothmul_pipelined_i_multiplicand_pip_4_9_port
                           , A2 => n1066, ZN => n2912);
   U87 : NOR2_X1 port map( A1 => n3078, A2 => n1067, ZN => n2934);
   U88 : CLKBUF_X1 port map( A => n2934, Z => n2923);
   U89 : NOR3_X1 port map( A1 => boothmul_pipelined_i_multiplicand_pip_4_8_port
                           , A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, A3 
                           => n3078, ZN => n2932);
   U90 : CLKBUF_X1 port map( A => n2932, Z => n2928);
   U91 : AOI22_X1 port map( A1 => n2923, A2 => 
                           boothmul_pipelined_i_muxes_in_4_175_port, B1 => 
                           n2928, B2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, ZN => 
                           n1068);
   U92 : INV_X1 port map( A => n1068, ZN => n1069);
   U93 : AOI221_X1 port map( B1 => boothmul_pipelined_i_muxes_in_4_50_port, B2 
                           => n2929, C1 => 
                           boothmul_pipelined_i_muxes_in_4_50_port, C2 => n2912
                           , A => n1069, ZN => n1070);
   U94 : INV_X1 port map( A => n1070, ZN => 
                           boothmul_pipelined_i_mux_out_4_24_port);
   U95 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           ZN => n3014);
   U96 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A => n3014, ZN => n1071);
   U97 : NOR2_X1 port map( A1 => n3081, A2 => n1071, ZN => n3051);
   U98 : CLKBUF_X1 port map( A => n3051, Z => n3039);
   U99 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, A2 
                           => n1071, ZN => n3043);
   U100 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_7_233_port, A2
                           => n3039, B1 => 
                           boothmul_pipelined_i_muxes_in_7_77_port, B2 => n3043
                           , ZN => n1072);
   U101 : INV_X1 port map( A => n1072, ZN => n2352);
   U102 : AND2_X1 port map( A1 => n2352, A2 => 
                           boothmul_pipelined_i_sum_B_in_7_14_port, ZN => n3087
                           );
   U103 : CLKBUF_X1 port map( A => DATA1(8), Z => n3096);
   U104 : CLKBUF_X1 port map( A => DATA1(15), Z => n3098);
   U105 : CLKBUF_X1 port map( A => DATA1(9), Z => n3097);
   U106 : INV_X1 port map( A => n2744, ZN => n3099);
   U107 : NOR2_X1 port map( A1 => n1073, A2 => n3077, ZN => n1081);
   U108 : AND2_X1 port map( A1 => n1081, A2 => 
                           boothmul_pipelined_i_sum_B_in_3_6_port, ZN => n3084)
                           ;
   U109 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n1074);
   U110 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n1074, ZN => n2822);
   U111 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           A2 => n2822, ZN => n1080);
   U112 : AND2_X1 port map( A1 => n1080, A2 => 
                           boothmul_pipelined_i_sum_B_in_2_4_port, ZN => n3085)
                           ;
   U113 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_73_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_73_port, ZN 
                           => n1075);
   U114 : INV_X1 port map( A => n1075, ZN => n1084);
   U115 : AND2_X1 port map( A1 => n1084, A2 => 
                           boothmul_pipelined_i_sum_B_in_6_12_port, ZN => n3088
                           );
   U116 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_205_port, B1 => 
                           n2961, B2 => 
                           boothmul_pipelined_i_muxes_in_5_205_port, ZN => 
                           n1076);
   U117 : INV_X1 port map( A => n1076, ZN => n1083);
   U118 : AND2_X1 port map( A1 => n1083, A2 => 
                           boothmul_pipelined_i_sum_B_in_5_10_port, ZN => n3089
                           );
   U119 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_65_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_65_port, ZN 
                           => n1077);
   U120 : INV_X1 port map( A => n1077, ZN => n1082);
   U121 : AND2_X1 port map( A1 => n1082, A2 => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, ZN => n3090)
                           ;
   U122 : INV_X1 port map( A => data1_mul_14_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port);
   U123 : INV_X1 port map( A => data1_mul_13_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port);
   U124 : INV_X1 port map( A => data1_mul_12_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port);
   U125 : INV_X1 port map( A => data1_mul_11_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port);
   U126 : INV_X1 port map( A => data1_mul_10_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port);
   U127 : INV_X1 port map( A => data1_mul_9_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port);
   U128 : INV_X1 port map( A => data1_mul_8_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port);
   U129 : INV_X1 port map( A => data1_mul_7_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port);
   U130 : INV_X1 port map( A => data1_mul_6_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port);
   U131 : INV_X1 port map( A => data1_mul_5_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port);
   U132 : INV_X1 port map( A => data1_mul_4_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port);
   U133 : INV_X1 port map( A => data1_mul_3_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port);
   U134 : INV_X1 port map( A => data1_mul_1_port, ZN => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port);
   U135 : INV_X1 port map( A => FUNC(2), ZN => n2730);
   U136 : NOR2_X1 port map( A1 => n2730, A2 => FUNC(0), ZN => n1094);
   U137 : AND2_X1 port map( A1 => n1919, A2 => n1094, ZN => n1267);
   U138 : INV_X1 port map( A => FUNC(3), ZN => n2743);
   U139 : NAND2_X1 port map( A1 => n1267, A2 => n2743, ZN => n553);
   U140 : XOR2_X1 port map( A => n1079, B => n1078, Z => n3086);
   U141 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_2_4_port, B => 
                           n1080, Z => n3091);
   U142 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_3_6_port, B => 
                           n1081, Z => n3092);
   U143 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_4_8_port, B => 
                           n1082, Z => n3093);
   U144 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_5_10_port, B => 
                           n1083, Z => n3094);
   U145 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_6_12_port, B => 
                           n1084, Z => n3095);
   U146 : NOR4_X1 port map( A1 => DATA2(6), A2 => DATA2(7), A3 => DATA2(8), A4 
                           => DATA2(9), ZN => n1092);
   U147 : INV_X1 port map( A => DATA2(0), ZN => n2778);
   U148 : INV_X1 port map( A => DATA2(1), ZN => n2777);
   U149 : NAND2_X1 port map( A1 => n2778, A2 => n2777, ZN => n1205);
   U150 : INV_X1 port map( A => n1205, ZN => n1465);
   U151 : INV_X1 port map( A => DATA2(3), ZN => n2775);
   U152 : INV_X1 port map( A => DATA2(5), ZN => n2773);
   U153 : INV_X1 port map( A => DATA2(4), ZN => n2774);
   U154 : NAND2_X1 port map( A1 => n2773, A2 => n2774, ZN => n1938);
   U155 : INV_X1 port map( A => n1938, ZN => n2512);
   U156 : NAND2_X1 port map( A1 => n2775, A2 => n2512, ZN => n1115);
   U157 : NOR2_X1 port map( A1 => n1115, A2 => DATA2(2), ZN => n1710);
   U158 : NAND2_X1 port map( A1 => n1465, A2 => n1710, ZN => n2474);
   U159 : INV_X1 port map( A => DATA2(10), ZN => n2766);
   U160 : INV_X1 port map( A => DATA2(11), ZN => n2765);
   U161 : INV_X1 port map( A => DATA2(12), ZN => n2764);
   U162 : INV_X1 port map( A => DATA2(13), ZN => n2763);
   U163 : NAND4_X1 port map( A1 => n2766, A2 => n2765, A3 => n2764, A4 => n2763
                           , ZN => n1085);
   U164 : NOR4_X1 port map( A1 => DATA2(15), A2 => DATA2(14), A3 => n2474, A4 
                           => n1085, ZN => n1091);
   U165 : NOR4_X1 port map( A1 => DATA1(15), A2 => DATA1(14), A3 => DATA1(13), 
                           A4 => DATA1(12), ZN => n1089);
   U166 : NOR4_X1 port map( A1 => DATA1(11), A2 => DATA1(10), A3 => DATA1(9), 
                           A4 => n3096, ZN => n1088);
   U167 : CLKBUF_X1 port map( A => DATA1(6), Z => n2582);
   U168 : CLKBUF_X1 port map( A => DATA1(4), Z => n1277);
   U169 : NOR4_X1 port map( A1 => DATA1(7), A2 => n2582, A3 => DATA1(5), A4 => 
                           n1277, ZN => n1087);
   U170 : NOR4_X1 port map( A1 => DATA1(3), A2 => DATA1(2), A3 => DATA1(1), A4 
                           => DATA1(0), ZN => n1086);
   U171 : AND4_X1 port map( A1 => n1089, A2 => n1088, A3 => n1087, A4 => n1086,
                           ZN => n1090);
   U172 : AOI211_X1 port map( C1 => n1092, C2 => n1091, A => n1090, B => n553, 
                           ZN => n2354);
   U173 : CLKBUF_X1 port map( A => n2354, Z => n2468);
   U174 : NAND2_X1 port map( A1 => FUNC(1), A2 => n1093, ZN => n2462);
   U175 : INV_X1 port map( A => n2462, ZN => n2438);
   U176 : INV_X1 port map( A => DATA2(9), ZN => n2767);
   U177 : NOR2_X1 port map( A1 => n2767, A2 => n3097, ZN => n2673);
   U178 : INV_X1 port map( A => n2673, ZN => n2611);
   U179 : NAND2_X1 port map( A1 => n3097, A2 => n2767, ZN => n2674);
   U180 : NAND2_X1 port map( A1 => n2611, A2 => n2674, ZN => n2565);
   U181 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_9_port, B1 => n2438
                           , B2 => n2565, ZN => n1286);
   U182 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(4), ZN => n1414);
   U183 : NOR2_X1 port map( A1 => n2777, A2 => n2775, ZN => n1096);
   U184 : INV_X1 port map( A => n1096, ZN => n1118);
   U185 : NOR2_X1 port map( A1 => n1414, A2 => n1118, ZN => n2552);
   U186 : NAND2_X1 port map( A1 => n1094, A2 => n2773, ZN => n1916);
   U187 : AOI211_X1 port map( C1 => n2552, C2 => DATA2(0), A => n1919, B => 
                           n1916, ZN => n1280);
   U188 : NAND2_X1 port map( A1 => FUNC(3), A2 => n1280, ZN => n2455);
   U189 : INV_X1 port map( A => n2455, ZN => n2736);
   U190 : NAND2_X1 port map( A1 => n1938, A2 => DATA2(3), ZN => n1994);
   U191 : NAND2_X1 port map( A1 => n2777, A2 => n1994, ZN => n1095);
   U192 : NAND2_X1 port map( A1 => n1414, A2 => n1994, ZN => n2521_port);
   U193 : NOR2_X1 port map( A1 => n2778, A2 => n1414, ZN => n1306);
   U194 : AOI21_X1 port map( B1 => n1095, B2 => n2521_port, A => n1306, ZN => 
                           n2526_port);
   U195 : INV_X1 port map( A => n2526_port, ZN => n2420);
   U196 : NOR2_X1 port map( A1 => n2778, A2 => n1118, ZN => n1415);
   U197 : AOI21_X1 port map( B1 => DATA2(2), B2 => n1415, A => n1938, ZN => 
                           n2357);
   U198 : INV_X1 port map( A => n2357, ZN => n2508);
   U199 : NAND2_X1 port map( A1 => n2508, A2 => n2512, ZN => n2510);
   U200 : INV_X1 port map( A => DATA2(2), ZN => n2776);
   U201 : OAI21_X1 port map( B1 => n2775, B2 => n2776, A => n2512, ZN => n1127)
                           ;
   U202 : NOR2_X1 port map( A1 => n1096, A2 => n1127, ZN => n2489);
   U203 : CLKBUF_X1 port map( A => n2489, Z => n1631);
   U204 : INV_X1 port map( A => n1631, ZN => n1843);
   U205 : INV_X1 port map( A => n1115, ZN => n1097);
   U206 : OAI21_X1 port map( B1 => n2777, B2 => n2776, A => n1097, ZN => n1975)
                           ;
   U207 : INV_X1 port map( A => n1975, ZN => n1694);
   U208 : CLKBUF_X1 port map( A => n1694, Z => n1752);
   U209 : INV_X1 port map( A => n1752, ZN => n2480);
   U210 : AOI21_X1 port map( B1 => DATA2(2), B2 => DATA2(0), A => n2480, ZN => 
                           n2211);
   U211 : CLKBUF_X1 port map( A => n2211, Z => n2483);
   U212 : INV_X1 port map( A => n2483, ZN => n2083);
   U213 : NAND3_X1 port map( A1 => n2778, A2 => DATA2(1), A3 => n1710, ZN => 
                           n2025);
   U214 : INV_X1 port map( A => DATA1(22), ZN => n2161);
   U215 : NOR2_X1 port map( A1 => n2025, A2 => n2161, ZN => n1550);
   U216 : NAND3_X1 port map( A1 => n2777, A2 => DATA2(0), A3 => n1710, ZN => 
                           n1968);
   U217 : INV_X1 port map( A => n1968, ZN => n2242);
   U218 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(21), ZN => n1543);
   U219 : INV_X1 port map( A => n2474, ZN => n1145);
   U220 : CLKBUF_X1 port map( A => n1145, Z => n2205);
   U221 : NAND2_X1 port map( A1 => DATA1(20), A2 => n2205, ZN => n1529);
   U222 : CLKBUF_X1 port map( A => n1710, Z => n1548);
   U223 : INV_X1 port map( A => n1548, ZN => n1829);
   U224 : OR3_X1 port map( A1 => n2778, A2 => n2777, A3 => n1829, ZN => n1691);
   U225 : INV_X1 port map( A => n1691, ZN => n2039);
   U226 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(23), ZN => n1577);
   U227 : NAND2_X1 port map( A1 => DATA1(24), A2 => n1829, ZN => n1098);
   U228 : NAND4_X1 port map( A1 => n1543, A2 => n1529, A3 => n1577, A4 => n1098
                           , ZN => n1099);
   U229 : NOR2_X1 port map( A1 => n1550, A2 => n1099, ZN => n1113);
   U230 : NOR4_X1 port map( A1 => n2776, A2 => n2778, A3 => n1115, A4 => 
                           DATA2(1), ZN => n1533);
   U231 : CLKBUF_X1 port map( A => n1533, Z => n1626);
   U232 : INV_X1 port map( A => n1626, ZN => n2081);
   U233 : INV_X1 port map( A => n1548, ZN => n2477);
   U234 : INV_X1 port map( A => DATA1(23), ZN => n2128);
   U235 : NOR2_X1 port map( A1 => n2025, A2 => n2128, ZN => n1556);
   U236 : INV_X1 port map( A => DATA1(21), ZN => n2700);
   U237 : NOR2_X1 port map( A1 => n2474, A2 => n2700, ZN => n1524);
   U238 : AOI211_X1 port map( C1 => DATA1(25), C2 => n2477, A => n1556, B => 
                           n1524, ZN => n1100);
   U239 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(22), ZN => n1539);
   U240 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(24), ZN => n1587);
   U241 : AND3_X1 port map( A1 => n1100, A2 => n1539, A3 => n1587, ZN => n1133)
                           ;
   U242 : INV_X1 port map( A => n1691, ZN => n1830);
   U243 : INV_X1 port map( A => DATA1(24), ZN => n2709);
   U244 : NOR2_X1 port map( A1 => n2025, A2 => n2709, ZN => n1579);
   U245 : INV_X1 port map( A => DATA1(26), ZN => n2557);
   U246 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(23), ZN => n1546);
   U247 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(22), ZN => n1542);
   U248 : OAI211_X1 port map( C1 => n1548, C2 => n2557, A => n1546, B => n1542,
                           ZN => n1101);
   U249 : AOI211_X1 port map( C1 => DATA1(25), C2 => n1830, A => n1579, B => 
                           n1101, ZN => n1138);
   U250 : OAI222_X1 port map( A1 => n2083, A2 => n1113, B1 => n2081, B2 => 
                           n1133, C1 => n1694, C2 => n1138, ZN => n1227);
   U251 : OAI21_X1 port map( B1 => n1115, B2 => DATA2(0), A => n2480, ZN => 
                           n1651);
   U252 : CLKBUF_X1 port map( A => n1651, Z => n2156);
   U253 : INV_X1 port map( A => n2156, ZN => n2213);
   U254 : INV_X1 port map( A => n2025, ZN => n2040);
   U255 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(20), ZN => n1544);
   U256 : NAND2_X1 port map( A1 => DATA1(21), A2 => n2039, ZN => n1547);
   U257 : CLKBUF_X1 port map( A => DATA1(18), Z => n2284);
   U258 : NAND2_X1 port map( A1 => n1145, A2 => n2284, ZN => n1102);
   U259 : AND3_X1 port map( A1 => n1544, A2 => n1547, A3 => n1102, ZN => n1103)
                           ;
   U260 : CLKBUF_X1 port map( A => DATA1(19), Z => n2256);
   U261 : NAND2_X1 port map( A1 => n2256, A2 => n2242, ZN => n1530);
   U262 : OAI211_X1 port map( C1 => n1548, C2 => n2161, A => n1103, B => n1530,
                           ZN => n1104);
   U263 : INV_X1 port map( A => n1104, ZN => n1112);
   U264 : INV_X1 port map( A => DATA1(16), ZN => n2691);
   U265 : NOR2_X1 port map( A1 => n2474, A2 => n2691, ZN => n1106);
   U266 : INV_X1 port map( A => DATA1(20), ZN => n2701);
   U267 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(17), ZN => n1500);
   U268 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(18), ZN => n1531);
   U269 : OAI211_X1 port map( C1 => n1548, C2 => n2701, A => n1500, B => n1531,
                           ZN => n1105);
   U270 : AOI211_X1 port map( C1 => n2039, C2 => DATA1(19), A => n1106, B => 
                           n1105, ZN => n1124);
   U271 : INV_X1 port map( A => DATA1(17), ZN => n2292);
   U272 : NOR2_X1 port map( A1 => n2474, A2 => n2292, ZN => n1108);
   U273 : NAND2_X1 port map( A1 => n2242, A2 => n2284, ZN => n1520);
   U274 : NAND2_X1 port map( A1 => n2040, A2 => n2256, ZN => n1527);
   U275 : OAI211_X1 port map( C1 => n1548, C2 => n2700, A => n1520, B => n1527,
                           ZN => n1107);
   U276 : AOI211_X1 port map( C1 => n2039, C2 => DATA1(20), A => n1108, B => 
                           n1107, ZN => n1123);
   U277 : INV_X1 port map( A => n1533, ZN => n1754);
   U278 : OAI222_X1 port map( A1 => n1112, A2 => n1694, B1 => n1124, B2 => 
                           n2083, C1 => n1123, C2 => n1754, ZN => n1151);
   U279 : INV_X1 port map( A => n1151, ZN => n1177);
   U280 : INV_X1 port map( A => n2211, ZN => n1174);
   U281 : NAND2_X1 port map( A1 => n2256, A2 => n2205, ZN => n1519);
   U282 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(20), ZN => n1526);
   U283 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(21), ZN => n1540);
   U284 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(22), ZN => n1554);
   U285 : AND3_X1 port map( A1 => n1526, A2 => n1540, A3 => n1554, ZN => n1109)
                           ;
   U286 : OAI211_X1 port map( C1 => n2128, C2 => n1548, A => n1519, B => n1109,
                           ZN => n1110);
   U287 : INV_X1 port map( A => n1110, ZN => n1114);
   U288 : OAI222_X1 port map( A1 => n1174, A2 => n1112, B1 => n2081, B2 => 
                           n1114, C1 => n1752, C2 => n1113, ZN => n1139);
   U289 : INV_X1 port map( A => n1139, ZN => n1111);
   U290 : NOR4_X1 port map( A1 => n2775, A2 => n1938, A3 => n1205, A4 => 
                           DATA2(2), ZN => n2127);
   U291 : INV_X1 port map( A => n2127, ZN => n2487);
   U292 : OAI22_X1 port map( A1 => n2213, A2 => n1177, B1 => n1111, B2 => n2487
                           , ZN => n1117);
   U293 : OAI222_X1 port map( A1 => n1114, A2 => n1752, B1 => n1123, B2 => 
                           n2083, C1 => n1112, C2 => n1754, ZN => n1150);
   U294 : INV_X1 port map( A => n1150, ZN => n1136);
   U295 : INV_X1 port map( A => n2494, ZN => n1977);
   U296 : OAI222_X1 port map( A1 => n1133, A2 => n1694, B1 => n1114, B2 => 
                           n2083, C1 => n1113, C2 => n1754, ZN => n1140);
   U297 : INV_X1 port map( A => n1140, ZN => n1161);
   U298 : NAND3_X1 port map( A1 => n1205, A2 => n1115, A3 => n2489, ZN => n2491
                           );
   U299 : OAI22_X1 port map( A1 => n1136, A2 => n1977, B1 => n1161, B2 => n2491
                           , ZN => n1116);
   U300 : AOI211_X1 port map( C1 => n1843, C2 => n1227, A => n1117, B => n1116,
                           ZN => n1242);
   U301 : NAND3_X1 port map( A1 => DATA2(0), A2 => DATA2(2), A3 => DATA2(3), ZN
                           => n1131);
   U302 : OAI21_X1 port map( B1 => n2776, B2 => n1118, A => n2512, ZN => n1848)
                           ;
   U303 : INV_X1 port map( A => n1848, ZN => n2501);
   U304 : NAND3_X1 port map( A1 => n1131, A2 => n2501, A3 => n1127, ZN => n2497
                           );
   U305 : OR2_X1 port map( A1 => n1415, A2 => n1127, ZN => n2499);
   U306 : INV_X1 port map( A => n2499, ZN => n2442);
   U307 : CLKBUF_X1 port map( A => n1843, Z => n1925);
   U308 : INV_X1 port map( A => n1651, ZN => n2485);
   U309 : INV_X1 port map( A => DATA1(14), ZN => n2578);
   U310 : NOR2_X1 port map( A1 => n2474, A2 => n2578, ZN => n1120);
   U311 : CLKBUF_X1 port map( A => DATA1(16), Z => n2315);
   U312 : NAND2_X1 port map( A1 => n2040, A2 => n2315, ZN => n1501);
   U313 : NAND2_X1 port map( A1 => n2242, A2 => n3098, ZN => n1511);
   U314 : OAI211_X1 port map( C1 => n1691, C2 => n2292, A => n1501, B => n1511,
                           ZN => n1119);
   U315 : AOI211_X1 port map( C1 => DATA1(18), C2 => n2477, A => n1120, B => 
                           n1119, ZN => n1171);
   U316 : NAND2_X1 port map( A1 => n2256, A2 => n1829, ZN => n1121);
   U317 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(17), ZN => n1521);
   U318 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(16), ZN => n1505);
   U319 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(15), ZN => n1516);
   U320 : NAND4_X1 port map( A1 => n1121, A2 => n1521, A3 => n1505, A4 => n1516
                           , ZN => n1122);
   U321 : AOI21_X1 port map( B1 => n2039, B2 => n2284, A => n1122, ZN => n1149)
                           ;
   U322 : OAI222_X1 port map( A1 => n1174, A2 => n1171, B1 => n2081, B2 => 
                           n1149, C1 => n1694, C2 => n1124, ZN => n1197);
   U323 : INV_X1 port map( A => n1197, ZN => n1154);
   U324 : OAI22_X1 port map( A1 => n2485, A2 => n1154, B1 => n1177, B2 => n2487
                           , ZN => n1126);
   U325 : OAI222_X1 port map( A1 => n1174, A2 => n1149, B1 => n2081, B2 => 
                           n1124, C1 => n1694, C2 => n1123, ZN => n1187);
   U326 : INV_X1 port map( A => n1187, ZN => n1128);
   U327 : CLKBUF_X1 port map( A => n1977, Z => n2214);
   U328 : OAI22_X1 port map( A1 => n1128, A2 => n2214, B1 => n1136, B2 => n2491
                           , ZN => n1125);
   U329 : AOI211_X1 port map( C1 => n1925, C2 => n1139, A => n1126, B => n1125,
                           ZN => n1202);
   U330 : INV_X1 port map( A => n1202, ZN => n1188);
   U331 : OR2_X1 port map( A1 => n1127, A2 => n2442, ZN => n1779);
   U332 : INV_X1 port map( A => n1779, ZN => n2506);
   U333 : INV_X1 port map( A => n2491, ZN => n1790);
   U334 : OAI22_X1 port map( A1 => n2485, A2 => n1128, B1 => n1136, B2 => n2487
                           , ZN => n1130);
   U335 : OAI22_X1 port map( A1 => n1631, A2 => n1161, B1 => n1177, B2 => n1977
                           , ZN => n1129);
   U336 : AOI211_X1 port map( C1 => n1790, C2 => n1139, A => n1130, B => n1129,
                           ZN => n1157);
   U337 : INV_X1 port map( A => n1157, ZN => n1189);
   U338 : AOI22_X1 port map( A1 => n2442, A2 => n1188, B1 => n2506, B2 => n1189
                           , ZN => n1144);
   U339 : NOR2_X1 port map( A1 => n1848, A2 => n1131, ZN => n1932);
   U340 : CLKBUF_X1 port map( A => n2127, Z => n2160);
   U341 : AOI22_X1 port map( A1 => n2160, A2 => n1140, B1 => n2494, B2 => n1139
                           , ZN => n1135);
   U342 : INV_X1 port map( A => DATA1(25), ZN => n2716);
   U343 : NOR2_X1 port map( A1 => n2025, A2 => n2716, ZN => n1589);
   U344 : INV_X1 port map( A => DATA1(27), ZN => n2059);
   U345 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(24), ZN => n1553);
   U346 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(23), ZN => n1538);
   U347 : OAI211_X1 port map( C1 => n1548, C2 => n2059, A => n1553, B => n1538,
                           ZN => n1132);
   U348 : AOI211_X1 port map( C1 => DATA1(26), C2 => n1830, A => n1589, B => 
                           n1132, ZN => n1160);
   U349 : OAI222_X1 port map( A1 => n1174, A2 => n1133, B1 => n2081, B2 => 
                           n1138, C1 => n1694, C2 => n1160, ZN => n1235);
   U350 : AOI22_X1 port map( A1 => n1790, A2 => n1227, B1 => n1925, B2 => n1235
                           , ZN => n1134);
   U351 : OAI211_X1 port map( C1 => n2213, C2 => n1136, A => n1135, B => n1134,
                           ZN => n1244);
   U352 : CLKBUF_X1 port map( A => n1848, Z => n1931);
   U353 : AOI22_X1 port map( A1 => DATA1(24), A2 => n2205, B1 => DATA1(28), B2 
                           => n1829, ZN => n1137);
   U354 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(25), ZN => n1576);
   U355 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(26), ZN => n1611);
   U356 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(27), ZN => n1709);
   U357 : AND4_X1 port map( A1 => n1137, A2 => n1576, A3 => n1611, A4 => n1709,
                           ZN => n1226);
   U358 : OAI222_X1 port map( A1 => n1226, A2 => n1752, B1 => n1138, B2 => 
                           n2083, C1 => n1160, C2 => n2081, ZN => n2155);
   U359 : INV_X1 port map( A => n2155, ZN => n1162);
   U360 : AOI22_X1 port map( A1 => n2160, A2 => n1227, B1 => n2156, B2 => n1139
                           , ZN => n1142);
   U361 : AOI22_X1 port map( A1 => n1790, A2 => n1235, B1 => n2494, B2 => n1140
                           , ZN => n1141);
   U362 : OAI211_X1 port map( C1 => n2489, C2 => n1162, A => n1142, B => n1141,
                           ZN => n2277);
   U363 : AOI22_X1 port map( A1 => n1932, A2 => n1244, B1 => n1931, B2 => n2277
                           , ZN => n1143);
   U364 : OAI211_X1 port map( C1 => n1242, C2 => n2497, A => n1144, B => n1143,
                           ZN => n1249);
   U365 : INV_X1 port map( A => n1249, ZN => n1220);
   U366 : AOI22_X1 port map( A1 => n2242, A2 => DATA1(14), B1 => n2039, B2 => 
                           n2315, ZN => n1148);
   U367 : NAND2_X1 port map( A1 => DATA1(17), A2 => n2477, ZN => n1147);
   U368 : NAND2_X1 port map( A1 => n2040, A2 => n3098, ZN => n1506);
   U369 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(13), ZN => n1146);
   U370 : NAND4_X1 port map( A1 => n1148, A2 => n1147, A3 => n1506, A4 => n1146
                           , ZN => n1183);
   U371 : INV_X1 port map( A => n1183, ZN => n1172);
   U372 : OAI222_X1 port map( A1 => n1174, A2 => n1172, B1 => n2081, B2 => 
                           n1171, C1 => n1694, C2 => n1149, ZN => n1212);
   U373 : AOI22_X1 port map( A1 => n2160, A2 => n1187, B1 => n2156, B2 => n1212
                           , ZN => n1153);
   U374 : AOI22_X1 port map( A1 => n1790, A2 => n1151, B1 => n1925, B2 => n1150
                           , ZN => n1152);
   U375 : OAI211_X1 port map( C1 => n1154, C2 => n2214, A => n1153, B => n1152,
                           ZN => n1213);
   U376 : INV_X1 port map( A => n1213, ZN => n1192);
   U377 : OAI22_X1 port map( A1 => n1192, A2 => n2499, B1 => n1202, B2 => n1779
                           , ZN => n1156);
   U378 : INV_X1 port map( A => n1932, ZN => n2503);
   U379 : OAI22_X1 port map( A1 => n1157, A2 => n2497, B1 => n1242, B2 => n2503
                           , ZN => n1155);
   U380 : AOI211_X1 port map( C1 => n1848, C2 => n1244, A => n1156, B => n1155,
                           ZN => n1219);
   U381 : INV_X1 port map( A => n2497, ZN => n2383);
   U382 : INV_X1 port map( A => n2277, ZN => n1247);
   U383 : OAI22_X1 port map( A1 => n1157, A2 => n2499, B1 => n1247, B2 => n2503
                           , ZN => n1167);
   U384 : AOI22_X1 port map( A1 => DATA1(25), A2 => n2205, B1 => DATA1(29), B2 
                           => n1829, ZN => n1159);
   U385 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(26), ZN => n1586);
   U386 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(27), ZN => n1624);
   U387 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(28), ZN => n1158);
   U388 : AND4_X1 port map( A1 => n1159, A2 => n1586, A3 => n1624, A4 => n1158,
                           ZN => n1234);
   U389 : OAI222_X1 port map( A1 => n1234, A2 => n1752, B1 => n1160, B2 => 
                           n2083, C1 => n1226, C2 => n2081, ZN => n2157);
   U390 : INV_X1 port map( A => n2157, ZN => n1230);
   U391 : OAI22_X1 port map( A1 => n1631, A2 => n1230, B1 => n2485, B2 => n1161
                           , ZN => n1165);
   U392 : INV_X1 port map( A => n1235, ZN => n1163);
   U393 : OAI22_X1 port map( A1 => n1163, A2 => n2487, B1 => n1162, B2 => n2491
                           , ZN => n1164);
   U394 : AOI211_X1 port map( C1 => n2494, C2 => n1227, A => n1165, B => n1164,
                           ZN => n1231);
   U395 : OAI22_X1 port map( A1 => n2501, A2 => n1231, B1 => n1242, B2 => n1779
                           , ZN => n1166);
   U396 : AOI211_X1 port map( C1 => n2383, C2 => n1244, A => n1167, B => n1166,
                           ZN => n1248);
   U397 : OAI222_X1 port map( A1 => n2510, A2 => n1220, B1 => n2508, B2 => 
                           n1219, C1 => n1248, C2 => n2512, ZN => n2392);
   U398 : INV_X1 port map( A => DATA1(15), ZN => n2577);
   U399 : NOR2_X1 port map( A1 => n1691, A2 => n2577, ZN => n1503);
   U400 : NOR2_X1 port map( A1 => n2025, A2 => n2578, ZN => n1513);
   U401 : NOR2_X1 port map( A1 => n1503, A2 => n1513, ZN => n1170);
   U402 : NAND2_X1 port map( A1 => DATA1(16), A2 => n1829, ZN => n1169);
   U403 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(13), ZN => n1601);
   U404 : CLKBUF_X1 port map( A => DATA1(12), Z => n2397);
   U405 : NAND2_X1 port map( A1 => n1145, A2 => n2397, ZN => n1168);
   U406 : NAND4_X1 port map( A1 => n1170, A2 => n1169, A3 => n1601, A4 => n1168
                           , ZN => n1196);
   U407 : INV_X1 port map( A => n1196, ZN => n1173);
   U408 : OAI222_X1 port map( A1 => n1174, A2 => n1173, B1 => n2081, B2 => 
                           n1172, C1 => n1752, C2 => n1171, ZN => n1294);
   U409 : AOI22_X1 port map( A1 => n2160, A2 => n1197, B1 => n2156, B2 => n1294
                           , ZN => n1176);
   U410 : AOI22_X1 port map( A1 => n1790, A2 => n1187, B1 => n2494, B2 => n1212
                           , ZN => n1175);
   U411 : OAI211_X1 port map( C1 => n1631, C2 => n1177, A => n1176, B => n1175,
                           ZN => n1295);
   U412 : AOI22_X1 port map( A1 => n2442, A2 => n1295, B1 => n2506, B2 => n1213
                           , ZN => n1179);
   U413 : CLKBUF_X1 port map( A => n1932, Z => n2373);
   U414 : AOI22_X1 port map( A1 => n2383, A2 => n1188, B1 => n2373, B2 => n1189
                           , ZN => n1178);
   U415 : OAI211_X1 port map( C1 => n2501, C2 => n1242, A => n1179, B => n1178,
                           ZN => n1180);
   U416 : INV_X1 port map( A => n1180, ZN => n1218);
   U417 : INV_X1 port map( A => DATA1(11), ZN => n2411);
   U418 : NOR2_X1 port map( A1 => n2474, A2 => n2411, ZN => n1181);
   U419 : NOR2_X1 port map( A1 => n1691, A2 => n2578, ZN => n1508);
   U420 : AOI211_X1 port map( C1 => n3098, C2 => n2477, A => n1181, B => n1508,
                           ZN => n1182);
   U421 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(13), ZN => n1517);
   U422 : NAND2_X1 port map( A1 => n2242, A2 => n2397, ZN => n1644);
   U423 : NAND3_X1 port map( A1 => n1182, A2 => n1517, A3 => n1644, ZN => n1208
                           );
   U424 : AOI222_X1 port map( A1 => n1183, A2 => n2480, B1 => n1208, B2 => 
                           n2483, C1 => n1196, C2 => n1626, ZN => n1332);
   U425 : INV_X1 port map( A => n1294, ZN => n1209);
   U426 : OAI22_X1 port map( A1 => n2485, A2 => n1332, B1 => n1209, B2 => n1977
                           , ZN => n1186);
   U427 : CLKBUF_X1 port map( A => n1790, Z => n2219);
   U428 : AOI22_X1 port map( A1 => n1212, A2 => n2160, B1 => n1197, B2 => n2219
                           , ZN => n1184);
   U429 : INV_X1 port map( A => n1184, ZN => n1185);
   U430 : AOI211_X1 port map( C1 => n1843, C2 => n1187, A => n1186, B => n1185,
                           ZN => n1335);
   U431 : INV_X1 port map( A => n1335, ZN => n1296);
   U432 : CLKBUF_X1 port map( A => n2442, Z => n2385);
   U433 : INV_X1 port map( A => n1779, ZN => n2384);
   U434 : AOI22_X1 port map( A1 => n1296, A2 => n2385, B1 => n1295, B2 => n2384
                           , ZN => n1191);
   U435 : AOI22_X1 port map( A1 => n1848, A2 => n1189, B1 => n1188, B2 => n1932
                           , ZN => n1190);
   U436 : OAI211_X1 port map( C1 => n2497, C2 => n1192, A => n1191, B => n1190,
                           ZN => n1193);
   U437 : INV_X1 port map( A => n1193, ZN => n1217);
   U438 : CLKBUF_X1 port map( A => DATA1(10), Z => n2576);
   U439 : INV_X1 port map( A => n2576, ZN => n2561);
   U440 : NOR2_X1 port map( A1 => n2474, A2 => n2561, ZN => n1693);
   U441 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(13), ZN => n1510);
   U442 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(12), ZN => n1600);
   U443 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(11), ZN => n1663);
   U444 : NAND3_X1 port map( A1 => n1510, A2 => n1600, A3 => n1663, ZN => n1194
                           );
   U445 : AOI211_X1 port map( C1 => DATA1(14), C2 => n2477, A => n1693, B => 
                           n1194, ZN => n1195);
   U446 : INV_X1 port map( A => n1195, ZN => n1290);
   U447 : AOI222_X1 port map( A1 => n2211, A2 => n1290, B1 => n1626, B2 => 
                           n1208, C1 => n2480, C2 => n1196, ZN => n1291);
   U448 : INV_X1 port map( A => n1291, ZN => n1367);
   U449 : AOI22_X1 port map( A1 => n2160, A2 => n1294, B1 => n2156, B2 => n1367
                           , ZN => n1199);
   U450 : AOI22_X1 port map( A1 => n2219, A2 => n1212, B1 => n1925, B2 => n1197
                           , ZN => n1198);
   U451 : OAI211_X1 port map( C1 => n1332, C2 => n2214, A => n1199, B => n1198,
                           ZN => n1370);
   U452 : AOI22_X1 port map( A1 => n2442, A2 => n1370, B1 => n2383, B2 => n1295
                           , ZN => n1201);
   U453 : AOI22_X1 port map( A1 => n2506, A2 => n1296, B1 => n2373, B2 => n1213
                           , ZN => n1200);
   U454 : OAI211_X1 port map( C1 => n2501, C2 => n1202, A => n1201, B => n1200,
                           ZN => n1203);
   U455 : INV_X1 port map( A => n1203, ZN => n1300);
   U456 : OAI222_X1 port map( A1 => n1218, A2 => n2512, B1 => n1217, B2 => 
                           n2510, C1 => n1300, C2 => n2508, ZN => n1372);
   U457 : INV_X1 port map( A => n1372, ZN => n1342);
   U458 : NAND2_X1 port map( A1 => n2776, A2 => n2775, ZN => n1204);
   U459 : OAI21_X1 port map( B1 => n1204, B2 => DATA2(1), A => n1938, ZN => 
                           n1206);
   U460 : OAI21_X1 port map( B1 => n1205, B2 => n1204, A => n1938, ZN => n2391)
                           ;
   U461 : CLKBUF_X1 port map( A => n2391, Z => n2517_port);
   U462 : INV_X1 port map( A => n2517_port, ZN => n2323);
   U463 : NAND2_X1 port map( A1 => n1206, A2 => n2323, ZN => n2293);
   U464 : OAI222_X1 port map( A1 => n2510, A2 => n1218, B1 => n2508, B2 => 
                           n1217, C1 => n1219, C2 => n2512, ZN => n1339);
   U465 : INV_X1 port map( A => n1339, ZN => n1302);
   U466 : NOR3_X1 port map( A1 => n2778, A2 => n2774, A3 => n2777, ZN => n1221)
                           ;
   U467 : NOR3_X1 port map( A1 => n2521_port, A2 => n1206, A3 => n1221, ZN => 
                           n2514);
   U468 : INV_X1 port map( A => n2514, ZN => n2268);
   U469 : OAI22_X1 port map( A1 => n1342, A2 => n2293, B1 => n1302, B2 => n2268
                           , ZN => n1223);
   U470 : INV_X1 port map( A => DATA1(13), ZN => n2649);
   U471 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(12), ZN => n1515);
   U472 : CLKBUF_X1 port map( A => DATA1(11), Z => n2678);
   U473 : NAND2_X1 port map( A1 => n2040, A2 => n2678, ZN => n1643);
   U474 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(10), ZN => n1676);
   U475 : AND3_X1 port map( A1 => n1515, A2 => n1643, A3 => n1676, ZN => n1207)
                           ;
   U476 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(9), ZN => n1268);
   U477 : OAI211_X1 port map( C1 => n1548, C2 => n2649, A => n1207, B => n1268,
                           ZN => n1331);
   U478 : AOI222_X1 port map( A1 => n1208, A2 => n2480, B1 => n1331, B2 => 
                           n2483, C1 => n1290, C2 => n1626, ZN => n1397);
   U479 : OAI22_X1 port map( A1 => n2485, A2 => n1397, B1 => n1332, B2 => n2487
                           , ZN => n1211);
   U480 : OAI22_X1 port map( A1 => n1291, A2 => n2214, B1 => n1209, B2 => n2491
                           , ZN => n1210);
   U481 : AOI211_X1 port map( C1 => n1925, C2 => n1212, A => n1211, B => n1210,
                           ZN => n1400);
   U482 : OAI22_X1 port map( A1 => n2499, A2 => n1400, B1 => n2497, B2 => n1335
                           , ZN => n1216);
   U483 : AOI22_X1 port map( A1 => n1932, A2 => n1295, B1 => n1931, B2 => n1213
                           , ZN => n1214);
   U484 : INV_X1 port map( A => n1214, ZN => n1215);
   U485 : AOI211_X1 port map( C1 => n1370, C2 => n2384, A => n1216, B => n1215,
                           ZN => n1338);
   U486 : OAI222_X1 port map( A1 => n2510, A2 => n1300, B1 => n2508, B2 => 
                           n1338, C1 => n1217, C2 => n2512, ZN => n1406);
   U487 : INV_X1 port map( A => n1406, ZN => n1301);
   U488 : OAI222_X1 port map( A1 => n1220, A2 => n2512, B1 => n1219, B2 => 
                           n2510, C1 => n1218, C2 => n2508, ZN => n2390);
   U489 : INV_X1 port map( A => n2390, ZN => n1303);
   U490 : INV_X1 port map( A => n2521_port, ZN => n1990);
   U491 : NAND2_X1 port map( A1 => n1990, A2 => n1221, ZN => n2525_port);
   U492 : OAI22_X1 port map( A1 => n2323, A2 => n1301, B1 => n1303, B2 => 
                           n2525_port, ZN => n1222);
   U493 : AOI211_X1 port map( C1 => n2521_port, C2 => n2392, A => n1223, B => 
                           n1222, ZN => n1409);
   U494 : INV_X1 port map( A => n1994, ZN => n2532_port);
   U495 : NOR4_X1 port map( A1 => n1414, A2 => n2777, A3 => DATA2(0), A4 => 
                           n2532_port, ZN => n2228);
   U496 : CLKBUF_X1 port map( A => n2228, Z => n2528_port);
   U497 : INV_X1 port map( A => n2528_port, ZN => n2153);
   U498 : INV_X1 port map( A => DATA1(28), ZN => n2723);
   U499 : NOR2_X1 port map( A1 => n2025, A2 => n2723, ZN => n1712);
   U500 : INV_X1 port map( A => DATA1(30), ZN => n2581);
   U501 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(27), ZN => n1610);
   U502 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(26), ZN => n1224);
   U503 : OAI211_X1 port map( C1 => n1548, C2 => n2581, A => n1610, B => n1224,
                           ZN => n1225);
   U504 : AOI211_X1 port map( C1 => DATA1(29), C2 => n2039, A => n1712, B => 
                           n1225, ZN => n2084);
   U505 : OAI222_X1 port map( A1 => n1174, A2 => n1226, B1 => n1754, B2 => 
                           n1234, C1 => n1752, C2 => n2084, ZN => n2159);
   U506 : AOI22_X1 port map( A1 => n2494, A2 => n1235, B1 => n1925, B2 => n2159
                           , ZN => n1229);
   U507 : AOI22_X1 port map( A1 => n2127, A2 => n2155, B1 => n1651, B2 => n1227
                           , ZN => n1228);
   U508 : OAI211_X1 port map( C1 => n1230, C2 => n2491, A => n1229, B => n1228,
                           ZN => n2274);
   U509 : INV_X1 port map( A => n2274, ZN => n1241);
   U510 : INV_X1 port map( A => n1231, ZN => n2275);
   U511 : INV_X1 port map( A => n2159, ZN => n1238);
   U512 : NOR2_X1 port map( A1 => n2474, A2 => n2059, ZN => n1233);
   U513 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(28), ZN => n1623);
   U514 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(29), ZN => n1831);
   U515 : OAI211_X1 port map( C1 => n1691, C2 => n2581, A => n1623, B => n1831,
                           ZN => n1232);
   U516 : AOI211_X1 port map( C1 => DATA1(31), C2 => n2477, A => n1233, B => 
                           n1232, ZN => n2082);
   U517 : OAI222_X1 port map( A1 => n1174, A2 => n1234, B1 => n1754, B2 => 
                           n2084, C1 => n1752, C2 => n2082, ZN => n2158);
   U518 : AOI22_X1 port map( A1 => n2494, A2 => n2155, B1 => n1843, B2 => n2158
                           , ZN => n1237);
   U519 : AOI22_X1 port map( A1 => n2160, A2 => n2157, B1 => n1651, B2 => n1235
                           , ZN => n1236);
   U520 : OAI211_X1 port map( C1 => n1238, C2 => n2491, A => n1237, B => n1236,
                           ZN => n2276);
   U521 : AOI22_X1 port map( A1 => n2383, A2 => n2275, B1 => n1931, B2 => n2276
                           , ZN => n1240);
   U522 : AOI22_X1 port map( A1 => n2442, A2 => n1244, B1 => n2384, B2 => n2277
                           , ZN => n1239);
   U523 : OAI211_X1 port map( C1 => n1241, C2 => n2503, A => n1240, B => n1239,
                           ZN => n2308);
   U524 : OAI22_X1 port map( A1 => n2499, A2 => n1242, B1 => n2501, B2 => n1241
                           , ZN => n1243);
   U525 : INV_X1 port map( A => n1243, ZN => n1246);
   U526 : AOI22_X1 port map( A1 => n2506, A2 => n1244, B1 => n2373, B2 => n2275
                           , ZN => n1245);
   U527 : OAI211_X1 port map( C1 => n1247, C2 => n2497, A => n1246, B => n1245,
                           ZN => n2309);
   U528 : INV_X1 port map( A => n2510, ZN => n2321);
   U529 : INV_X1 port map( A => n1248, ZN => n1250);
   U530 : CLKBUF_X1 port map( A => n2357, Z => n1936);
   U531 : AOI222_X1 port map( A1 => n2308, A2 => n1938, B1 => n2309, B2 => 
                           n2321, C1 => n1250, C2 => n1936, ZN => n2343);
   U532 : INV_X1 port map( A => n2293, ZN => n2518_port);
   U533 : AOI22_X1 port map( A1 => n2518_port, A2 => n2390, B1 => n2514, B2 => 
                           n2392, ZN => n1252);
   U534 : INV_X1 port map( A => n2525_port, ZN => n2388);
   U535 : AOI222_X1 port map( A1 => n2309, A2 => n1938, B1 => n1250, B2 => 
                           n2321, C1 => n1249, C2 => n2357, ZN => n1255);
   U536 : INV_X1 port map( A => n1255, ZN => n2389);
   U537 : AOI22_X1 port map( A1 => n2388, A2 => n2389, B1 => n2517_port, B2 => 
                           n1339, ZN => n1251);
   U538 : OAI211_X1 port map( C1 => n1990, C2 => n2343, A => n1252, B => n1251,
                           ZN => n2430);
   U539 : INV_X1 port map( A => n2430, ZN => n2421);
   U540 : NAND3_X1 port map( A1 => n2777, A2 => n1994, A3 => n1306, ZN => 
                           n2537_port);
   U541 : CLKBUF_X1 port map( A => n2514, Z => n2366);
   U542 : AOI22_X1 port map( A1 => n2366, A2 => n2390, B1 => n2391, B2 => n1372
                           , ZN => n1254);
   U543 : AOI22_X1 port map( A1 => n2518_port, A2 => n1339, B1 => n2388, B2 => 
                           n2392, ZN => n1253);
   U544 : OAI211_X1 port map( C1 => n1990, C2 => n1255, A => n1254, B => n1253,
                           ZN => n2429);
   U545 : INV_X1 port map( A => n2429, ZN => n1326);
   U546 : OAI222_X1 port map( A1 => n2420, A2 => n1409, B1 => n2153, B2 => 
                           n2421, C1 => n2537_port, C2 => n1326, ZN => n1266);
   U547 : NOR2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n1262);
   U548 : NAND2_X1 port map( A1 => n3097, A2 => DATA2_I_9_port, ZN => n2436);
   U549 : OAI21_X1 port map( B1 => DATA1(9), B2 => DATA2_I_9_port, A => n2436, 
                           ZN => n1880);
   U550 : NOR2_X1 port map( A1 => n1262, A2 => n1880, ZN => n2452);
   U551 : INV_X1 port map( A => DATA1(7), ZN => n2667);
   U552 : XNOR2_X1 port map( A => n2667, B => DATA2_I_7_port, ZN => n1352);
   U553 : INV_X1 port map( A => DATA1(5), ZN => n2600);
   U554 : XOR2_X1 port map( A => n2600, B => DATA2_I_5_port, Z => n1418);
   U555 : INV_X1 port map( A => n1418, ZN => n1420);
   U556 : INV_X1 port map( A => DATA1(3), ZN => n1463);
   U557 : XNOR2_X1 port map( A => n1463, B => DATA2_I_3_port, ZN => n1495);
   U558 : NAND2_X1 port map( A1 => DATA1(2), A2 => DATA2_I_2_port, ZN => n1320)
                           ;
   U559 : OAI21_X1 port map( B1 => DATA1(2), B2 => DATA2_I_2_port, A => n1320, 
                           ZN => n2006);
   U560 : NAND2_X1 port map( A1 => DATA1(1), A2 => DATA2_I_1_port, ZN => n1318)
                           ;
   U561 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n2244)
                           ;
   U562 : INV_X1 port map( A => n2244, ZN => n2460);
   U563 : NOR2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n2459);
   U564 : OAI21_X1 port map( B1 => DATA1(1), B2 => DATA2_I_1_port, A => n1318, 
                           ZN => n2243);
   U565 : NOR2_X1 port map( A1 => n2459, A2 => n2243, ZN => n2202);
   U566 : OAI21_X1 port map( B1 => cin, B2 => n2460, A => n2202, ZN => n1256);
   U567 : OAI221_X1 port map( B1 => n2006, B2 => n1318, C1 => n2006, C2 => 
                           n1256, A => n1320, ZN => n1257);
   U568 : AND2_X1 port map( A1 => DATA1(3), A2 => DATA2_I_3_port, ZN => n1322);
   U569 : AOI21_X1 port map( B1 => n1495, B2 => n1257, A => n1322, ZN => n1258)
                           ;
   U570 : NAND2_X1 port map( A1 => n1277, A2 => DATA2_I_4_port, ZN => n1323);
   U571 : OAI21_X1 port map( B1 => n1277, B2 => DATA2_I_4_port, A => n1323, ZN 
                           => n1459);
   U572 : OAI21_X1 port map( B1 => n1258, B2 => n1459, A => n1323, ZN => n1259)
                           ;
   U573 : AND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n1324);
   U574 : AOI21_X1 port map( B1 => n1420, B2 => n1259, A => n1324, ZN => n1260)
                           ;
   U575 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n1325)
                           ;
   U576 : OAI21_X1 port map( B1 => DATA1(6), B2 => DATA2_I_6_port, A => n1325, 
                           ZN => n1383);
   U577 : OAI21_X1 port map( B1 => n1260, B2 => n1383, A => n1325, ZN => n1261)
                           ;
   U578 : AOI22_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, B1 => n1352,
                           B2 => n1261, ZN => n1881);
   U579 : NOR2_X1 port map( A1 => n3099, A2 => n1881, ZN => n2451);
   U580 : INV_X1 port map( A => n2451, ZN => n2347);
   U581 : AOI211_X1 port map( C1 => n1262, C2 => n1880, A => n2452, B => n2347,
                           ZN => n1265);
   U582 : NAND2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n1287)
                           ;
   U583 : INV_X1 port map( A => DATA1(8), ZN => n2609);
   U584 : INV_X1 port map( A => DATA2_I_8_port, ZN => n1263);
   U585 : NOR3_X1 port map( A1 => n2609, A2 => n1880, A3 => n1263, ZN => n1884)
                           ;
   U586 : NAND2_X1 port map( A1 => n2744, A2 => n1881, ZN => n2433);
   U587 : AOI211_X1 port map( C1 => n1880, C2 => n1287, A => n1884, B => n2433,
                           ZN => n1264);
   U588 : AOI211_X1 port map( C1 => n2736, C2 => n1266, A => n1265, B => n1264,
                           ZN => n1285);
   U589 : OR2_X1 port map( A1 => n2462, A2 => FUNC(3), ZN => n2437);
   U590 : INV_X1 port map( A => n2437, ZN => n2410);
   U591 : NAND2_X1 port map( A1 => FUNC(3), A2 => n1267, ZN => n2458);
   U592 : INV_X1 port map( A => n2458, ZN => n2412);
   U593 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => n3097, B => 
                           DATA2(9), ZN => n1284);
   U594 : NOR2_X1 port map( A1 => n2025, A2 => n2667, ZN => n1392);
   U595 : NAND2_X1 port map( A1 => n2242, A2 => n3096, ZN => n1329);
   U596 : OAI211_X1 port map( C1 => n1548, C2 => n2600, A => n1268, B => n1329,
                           ZN => n1269);
   U597 : AOI211_X1 port map( C1 => n2582, C2 => n2039, A => n1392, B => n1269,
                           ZN => n1753);
   U598 : NOR2_X1 port map( A1 => n2474, A2 => n2609, ZN => n1288);
   U599 : NAND2_X1 port map( A1 => n2040, A2 => n2582, ZN => n1428);
   U600 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(5), ZN => n1973);
   U601 : OAI211_X1 port map( C1 => n2667, C2 => n1968, A => n1428, B => n1973,
                           ZN => n1270);
   U602 : AOI211_X1 port map( C1 => n1277, C2 => n2477, A => n1288, B => n1270,
                           ZN => n1751);
   U603 : INV_X1 port map( A => n2582, ZN => n2580);
   U604 : NOR2_X1 port map( A1 => n1968, A2 => n2580, ZN => n1391);
   U605 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(7), ZN => n1327);
   U606 : NAND2_X1 port map( A1 => n2039, A2 => n1277, ZN => n2209);
   U607 : OAI211_X1 port map( C1 => n1548, C2 => n1463, A => n1327, B => n2209,
                           ZN => n1271);
   U608 : AOI211_X1 port map( C1 => DATA1(5), C2 => n2040, A => n1391, B => 
                           n1271, ZN => n1276);
   U609 : OAI222_X1 port map( A1 => n1174, A2 => n1753, B1 => n1754, B2 => 
                           n1751, C1 => n1752, C2 => n1276, ZN => n1791);
   U610 : INV_X1 port map( A => n1791, ZN => n1930);
   U611 : NOR2_X1 port map( A1 => n1968, A2 => n2600, ZN => n1431);
   U612 : INV_X1 port map( A => DATA1(2), ZN => n2658);
   U613 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(6), ZN => n1361);
   U614 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(3), ZN => n2472);
   U615 : OAI211_X1 port map( C1 => n1710, C2 => n2658, A => n1361, B => n2472,
                           ZN => n1272);
   U616 : AOI211_X1 port map( C1 => DATA1(4), C2 => n2040, A => n1431, B => 
                           n1272, ZN => n1279);
   U617 : OAI222_X1 port map( A1 => n1174, A2 => n1751, B1 => n1754, B2 => 
                           n1276, C1 => n1752, C2 => n1279, ZN => n1927);
   U618 : INV_X1 port map( A => n1927, ZN => n1273);
   U619 : OAI22_X1 port map( A1 => n2485, A2 => n1930, B1 => n1273, B2 => n1977
                           , ZN => n1282);
   U620 : INV_X1 port map( A => DATA1(1), ZN => n2651);
   U621 : INV_X1 port map( A => n1277, ZN => n2660);
   U622 : NOR2_X1 port map( A1 => n1968, A2 => n2660, ZN => n1467);
   U623 : NOR2_X1 port map( A1 => n2025, A2 => n1463, ZN => n2207);
   U624 : AOI211_X1 port map( C1 => DATA1(2), C2 => n1830, A => n1467, B => 
                           n2207, ZN => n1274);
   U625 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(5), ZN => n1393);
   U626 : OAI211_X1 port map( C1 => n1548, C2 => n2651, A => n1274, B => n1393,
                           ZN => n1275);
   U627 : INV_X1 port map( A => n1275, ZN => n1385);
   U628 : OAI222_X1 port map( A1 => n1385, A2 => n1694, B1 => n1276, B2 => 
                           n2083, C1 => n1279, C2 => n2081, ZN => n1926);
   U629 : INV_X1 port map( A => n1926, ZN => n1315);
   U630 : NOR2_X1 port map( A1 => n1968, A2 => n1463, ZN => n1971);
   U631 : INV_X1 port map( A => DATA1(0), ZN => n2650);
   U632 : NAND2_X1 port map( A1 => n1145, A2 => n1277, ZN => n1429);
   U633 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(2), ZN => n2473);
   U634 : OAI211_X1 port map( C1 => n1548, C2 => n2650, A => n1429, B => n2473,
                           ZN => n1278);
   U635 : AOI211_X1 port map( C1 => DATA1(1), C2 => n2039, A => n1971, B => 
                           n1278, ZN => n1424);
   U636 : OAI222_X1 port map( A1 => n1174, A2 => n1279, B1 => n1754, B2 => 
                           n1385, C1 => n1752, C2 => n1424, ZN => n1924);
   U637 : INV_X1 port map( A => n1924, ZN => n1356);
   U638 : OAI22_X1 port map( A1 => n1315, A2 => n2487, B1 => n1356, B2 => n2491
                           , ZN => n1281);
   U639 : NAND2_X1 port map( A1 => n1280, A2 => n2743, ZN => n2427);
   U640 : INV_X1 port map( A => n2427, ZN => n2441);
   U641 : OAI21_X1 port map( B1 => n1282, B2 => n1281, A => n2441, ZN => n1283)
                           ;
   U642 : NAND4_X1 port map( A1 => n1286, A2 => n1285, A3 => n1284, A4 => n1283
                           , ZN => OUTALU(9));
   U643 : OAI21_X1 port map( B1 => DATA1(8), B2 => DATA2_I_8_port, A => n1287, 
                           ZN => n1879);
   U644 : INV_X1 port map( A => n1879, ZN => n1314);
   U645 : OAI22_X1 port map( A1 => n1409, A2 => n2537_port, B1 => n1326, B2 => 
                           n2153, ZN => n1312);
   U646 : AOI21_X1 port map( B1 => DATA1(12), B2 => n2477, A => n1288, ZN => 
                           n1289);
   U647 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(11), ZN => n1599);
   U648 : NAND2_X1 port map( A1 => n2040, A2 => n2576, ZN => n1662);
   U649 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(9), ZN => n1690);
   U650 : NAND4_X1 port map( A1 => n1289, A2 => n1599, A3 => n1662, A4 => n1690
                           , ZN => n1364);
   U651 : AOI222_X1 port map( A1 => n1290, A2 => n2480, B1 => n1364, B2 => 
                           n2483, C1 => n1331, C2 => n1626, ZN => n1435);
   U652 : OAI22_X1 port map( A1 => n2485, A2 => n1435, B1 => n1291, B2 => n2487
                           , ZN => n1293);
   U653 : OAI22_X1 port map( A1 => n1332, A2 => n2491, B1 => n1397, B2 => n1977
                           , ZN => n1292);
   U654 : AOI211_X1 port map( C1 => n1925, C2 => n1294, A => n1293, B => n1292,
                           ZN => n1439);
   U655 : INV_X1 port map( A => n1439, ZN => n1403);
   U656 : AOI22_X1 port map( A1 => n2442, A2 => n1403, B1 => n2383, B2 => n1370
                           , ZN => n1298);
   U657 : AOI22_X1 port map( A1 => n1932, A2 => n1296, B1 => n1931, B2 => n1295
                           , ZN => n1297);
   U658 : OAI211_X1 port map( C1 => n1400, C2 => n1779, A => n1298, B => n1297,
                           ZN => n1299);
   U659 : INV_X1 port map( A => n1299, ZN => n1371);
   U660 : OAI222_X1 port map( A1 => n1300, A2 => n2512, B1 => n1338, B2 => 
                           n2510, C1 => n1371, C2 => n2508, ZN => n1405);
   U661 : INV_X1 port map( A => n1405, ZN => n1445);
   U662 : OAI22_X1 port map( A1 => n2323, A2 => n1445, B1 => n1301, B2 => n2293
                           , ZN => n1305);
   U663 : OAI22_X1 port map( A1 => n1990, A2 => n1303, B1 => n1302, B2 => 
                           n2525_port, ZN => n1304);
   U664 : AOI211_X1 port map( C1 => n2366, C2 => n1372, A => n1305, B => n1304,
                           ZN => n1448);
   U665 : NAND3_X1 port map( A1 => DATA2(1), A2 => n1306, A3 => n1994, ZN => 
                           n2147);
   U666 : OAI22_X1 port map( A1 => n1448, A2 => n2420, B1 => n2421, B2 => n2147
                           , ZN => n1311);
   U667 : AOI222_X1 port map( A1 => n1927, A2 => n1651, B1 => n1926, B2 => 
                           n2494, C1 => n1924, C2 => n2160, ZN => n1309);
   U668 : CLKBUF_X1 port map( A => n2354, Z => n2449);
   U669 : INV_X1 port map( A => DATA2(8), ZN => n2768);
   U670 : OAI22_X1 port map( A1 => n2609, A2 => DATA2(8), B1 => n2768, B2 => 
                           n3096, ZN => n2604);
   U671 : AOI22_X1 port map( A1 => n2449, A2 => dataout_mul_8_port, B1 => n2438
                           , B2 => n2604, ZN => n1308);
   U672 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => n3096, B => 
                           DATA2(8), ZN => n1307);
   U673 : OAI211_X1 port map( C1 => n1309, C2 => n2427, A => n1308, B => n1307,
                           ZN => n1310);
   U674 : AOI221_X1 port map( B1 => n1312, B2 => n2736, C1 => n1311, C2 => 
                           n2736, A => n1310, ZN => n1313);
   U675 : OAI221_X1 port map( B1 => n1314, B2 => n2347, C1 => n1879, C2 => 
                           n2433, A => n1313, ZN => OUTALU(8));
   U676 : OAI22_X1 port map( A1 => n2485, A2 => n1315, B1 => n1356, B2 => n2214
                           , ZN => n1317);
   U677 : OAI221_X1 port map( B1 => DATA1(7), B2 => n2462, C1 => n2667, C2 => 
                           n2458, A => n2437, ZN => n1316);
   U678 : AOI22_X1 port map( A1 => n2441, A2 => n1317, B1 => DATA2(7), B2 => 
                           n1316, ZN => n1355);
   U679 : NOR2_X1 port map( A1 => DATA2(7), A2 => n2667, ZN => n2605);
   U680 : AOI22_X1 port map( A1 => n2449, A2 => dataout_mul_7_port, B1 => n2438
                           , B2 => n2605, ZN => n1354);
   U681 : NOR2_X1 port map( A1 => cin, A2 => n3099, ZN => n2466);
   U682 : INV_X1 port map( A => n2466, ZN => n1969);
   U683 : INV_X1 port map( A => n2243, ZN => n2245);
   U684 : INV_X1 port map( A => n1318, ZN => n1319);
   U685 : AOI21_X1 port map( B1 => n2460, B2 => n2245, A => n1319, ZN => n2005)
                           ;
   U686 : OAI21_X1 port map( B1 => n2005, B2 => n2006, A => n1320, ZN => n1490)
                           ;
   U687 : AOI21_X1 port map( B1 => n1495, B2 => n1490, A => n1322, ZN => n1454)
                           ;
   U688 : OAI21_X1 port map( B1 => n1454, B2 => n1459, A => n1323, ZN => n1389)
                           ;
   U689 : AOI21_X1 port map( B1 => n1420, B2 => n1389, A => n1324, ZN => n1378)
                           ;
   U690 : OAI21_X1 port map( B1 => n1378, B2 => n1383, A => n1325, ZN => n1347)
                           ;
   U691 : NAND2_X1 port map( A1 => n2744, A2 => cin, ZN => n2461);
   U692 : NOR2_X1 port map( A1 => n1319, A2 => n2202, ZN => n2003);
   U693 : OAI21_X1 port map( B1 => n2003, B2 => n2006, A => n1320, ZN => n1494)
                           ;
   U694 : NAND2_X1 port map( A1 => n1495, A2 => n1494, ZN => n1493);
   U695 : INV_X1 port map( A => n1493, ZN => n1321);
   U696 : NOR2_X1 port map( A1 => n1322, A2 => n1321, ZN => n1453);
   U697 : OAI21_X1 port map( B1 => n1453, B2 => n1459, A => n1323, ZN => n1388)
                           ;
   U698 : AOI21_X1 port map( B1 => n1420, B2 => n1388, A => n1324, ZN => n1377)
                           ;
   U699 : OAI21_X1 port map( B1 => n1377, B2 => n1383, A => n1325, ZN => n1346)
                           ;
   U700 : OAI22_X1 port map( A1 => n1969, A2 => n1347, B1 => n2461, B2 => n1346
                           , ZN => n1351);
   U701 : OAI22_X1 port map( A1 => n1448, A2 => n2537_port, B1 => n1326, B2 => 
                           n2147, ZN => n1344);
   U702 : INV_X1 port map( A => n1327, ZN => n1328);
   U703 : AOI21_X1 port map( B1 => n2678, B2 => n2477, A => n1328, ZN => n1330)
                           ;
   U704 : NAND2_X1 port map( A1 => n2039, A2 => DATA1(10), ZN => n1642);
   U705 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(9), ZN => n1675);
   U706 : NAND4_X1 port map( A1 => n1330, A2 => n1642, A3 => n1675, A4 => n1329
                           , ZN => n1396);
   U707 : AOI222_X1 port map( A1 => n1331, A2 => n2480, B1 => n1396, B2 => 
                           n2483, C1 => n1364, C2 => n1626, ZN => n1471);
   U708 : OAI22_X1 port map( A1 => n2213, A2 => n1471, B1 => n1397, B2 => n2487
                           , ZN => n1334);
   U709 : OAI22_X1 port map( A1 => n1631, A2 => n1332, B1 => n1435, B2 => n1977
                           , ZN => n1333);
   U710 : AOI211_X1 port map( C1 => n2219, C2 => n1367, A => n1334, B => n1333,
                           ZN => n1474);
   U711 : OAI22_X1 port map( A1 => n1400, A2 => n2497, B1 => n1474, B2 => n2499
                           , ZN => n1337);
   U712 : OAI22_X1 port map( A1 => n2501, A2 => n1335, B1 => n1439, B2 => n1779
                           , ZN => n1336);
   U713 : AOI211_X1 port map( C1 => n2373, C2 => n1370, A => n1337, B => n1336,
                           ZN => n1404);
   U714 : OAI222_X1 port map( A1 => n1338, A2 => n2512, B1 => n1371, B2 => 
                           n2510, C1 => n1404, C2 => n2508, ZN => n1360);
   U715 : AOI22_X1 port map( A1 => n2518_port, A2 => n1405, B1 => n2517_port, 
                           B2 => n1360, ZN => n1341);
   U716 : AOI22_X1 port map( A1 => n2514, A2 => n1406, B1 => n2521_port, B2 => 
                           n1339, ZN => n1340);
   U717 : OAI211_X1 port map( C1 => n1342, C2 => n2525_port, A => n1341, B => 
                           n1340, ZN => n1484);
   U718 : INV_X1 port map( A => n1484, ZN => n1449);
   U719 : OAI22_X1 port map( A1 => n1449, A2 => n2420, B1 => n1409, B2 => n2153
                           , ZN => n1343);
   U720 : AOI211_X1 port map( C1 => n2532_port, C2 => n2430, A => n1344, B => 
                           n1343, ZN => n1413);
   U721 : NAND2_X1 port map( A1 => DATA2(0), A2 => DATA2(3), ZN => n1345);
   U722 : AOI211_X1 port map( C1 => n2776, C2 => n2777, A => n2775, B => n2774,
                           ZN => n2538_port);
   U723 : INV_X1 port map( A => n2538_port, ZN => n1996);
   U724 : OAI21_X1 port map( B1 => n2774, B2 => n1345, A => n1996, ZN => n1999)
                           ;
   U725 : NOR3_X1 port map( A1 => n1413, A2 => n2455, A3 => n1999, ZN => n1350)
                           ;
   U726 : INV_X1 port map( A => n2461, ZN => n2004);
   U727 : AOI22_X1 port map( A1 => n2466, A2 => n1347, B1 => n2004, B2 => n1346
                           , ZN => n1348);
   U728 : NOR2_X1 port map( A1 => n1348, A2 => n1352, ZN => n1349);
   U729 : AOI211_X1 port map( C1 => n1352, C2 => n1351, A => n1350, B => n1349,
                           ZN => n1353);
   U730 : NAND3_X1 port map( A1 => n1355, A2 => n1354, A3 => n1353, ZN => 
                           OUTALU(7));
   U731 : AOI22_X1 port map( A1 => n2466, A2 => n1378, B1 => n2004, B2 => n1377
                           , ZN => n1384);
   U732 : NOR3_X1 port map( A1 => n2213, A2 => n1356, A3 => n2427, ZN => n1359)
                           ;
   U733 : INV_X1 port map( A => DATA2(6), ZN => n2772);
   U734 : AOI22_X1 port map( A1 => n2582, A2 => n2772, B1 => DATA2(6), B2 => 
                           n2580, ZN => n2664);
   U735 : AOI21_X1 port map( B1 => n2582, B2 => n2412, A => n2410, ZN => n1357)
                           ;
   U736 : OAI22_X1 port map( A1 => n2664, A2 => n2462, B1 => n1357, B2 => n2772
                           , ZN => n1358);
   U737 : AOI211_X1 port map( C1 => dataout_mul_6_port, C2 => n2449, A => n1359
                           , B => n1358, ZN => n1382);
   U738 : CLKBUF_X1 port map( A => n1999, Z => n2113);
   U739 : INV_X1 port map( A => n2113, ZN => n2541_port);
   U740 : NOR2_X1 port map( A1 => n2538_port, A2 => n2541_port, ZN => 
                           n2543_port);
   U741 : INV_X1 port map( A => n2543_port, ZN => n2100);
   U742 : OAI22_X1 port map( A1 => n1449, A2 => n2537_port, B1 => n1409, B2 => 
                           n2147, ZN => n1376);
   U743 : INV_X1 port map( A => n1360, ZN => n1482);
   U744 : NAND2_X1 port map( A1 => DATA1(10), A2 => n2477, ZN => n1362);
   U745 : NAND2_X1 port map( A1 => n2039, A2 => n3097, ZN => n1661);
   U746 : NAND2_X1 port map( A1 => n2040, A2 => DATA1(8), ZN => n1689);
   U747 : AND4_X1 port map( A1 => n1362, A2 => n1661, A3 => n1689, A4 => n1361,
                           ZN => n1363);
   U748 : OAI21_X1 port map( B1 => n1968, B2 => n2667, A => n1363, ZN => n1433)
                           ;
   U749 : AOI222_X1 port map( A1 => n1364, A2 => n2480, B1 => n1433, B2 => 
                           n2483, C1 => n1396, C2 => n1626, ZN => n1978);
   U750 : OAI22_X1 port map( A1 => n2213, A2 => n1978, B1 => n1435, B2 => n2487
                           , ZN => n1366);
   U751 : OAI22_X1 port map( A1 => n1397, A2 => n2491, B1 => n1471, B2 => n1977
                           , ZN => n1365);
   U752 : AOI211_X1 port map( C1 => n1843, C2 => n1367, A => n1366, B => n1365,
                           ZN => n1982);
   U753 : OAI22_X1 port map( A1 => n1439, A2 => n2497, B1 => n1982, B2 => n2499
                           , ZN => n1369);
   U754 : OAI22_X1 port map( A1 => n1400, A2 => n2503, B1 => n1474, B2 => n1779
                           , ZN => n1368);
   U755 : AOI211_X1 port map( C1 => n1848, C2 => n1370, A => n1369, B => n1368,
                           ZN => n1443);
   U756 : OAI222_X1 port map( A1 => n1371, A2 => n2512, B1 => n1404, B2 => 
                           n2510, C1 => n1443, C2 => n2508, ZN => n1479);
   U757 : AOI22_X1 port map( A1 => n2366, A2 => n1405, B1 => n2391, B2 => n1479
                           , ZN => n1374);
   U758 : AOI22_X1 port map( A1 => n2388, A2 => n1406, B1 => n2521_port, B2 => 
                           n1372, ZN => n1373);
   U759 : OAI211_X1 port map( C1 => n1482, C2 => n2293, A => n1374, B => n1373,
                           ZN => n1483);
   U760 : INV_X1 port map( A => n1483, ZN => n1995);
   U761 : OAI22_X1 port map( A1 => n1448, A2 => n2153, B1 => n1995, B2 => n2420
                           , ZN => n1375);
   U762 : AOI211_X1 port map( C1 => n2532_port, C2 => n2429, A => n1376, B => 
                           n1375, ZN => n1452);
   U763 : OAI22_X1 port map( A1 => n1413, A2 => n2100, B1 => n1452, B2 => n1999
                           , ZN => n1380);
   U764 : OAI22_X1 port map( A1 => n1378, A2 => n1969, B1 => n1377, B2 => n2461
                           , ZN => n1379);
   U765 : AOI22_X1 port map( A1 => n2736, A2 => n1380, B1 => n1383, B2 => n1379
                           , ZN => n1381);
   U766 : OAI211_X1 port map( C1 => n1384, C2 => n1383, A => n1382, B => n1381,
                           ZN => OUTALU(6));
   U767 : OAI21_X1 port map( B1 => n2600, B2 => n2458, A => n2437, ZN => n1387)
                           ;
   U768 : OAI22_X1 port map( A1 => n1385, A2 => n2083, B1 => n1424, B2 => n2081
                           , ZN => n1386);
   U769 : AOI22_X1 port map( A1 => DATA2(5), A2 => n1387, B1 => n2441, B2 => 
                           n1386, ZN => n1423);
   U770 : AOI22_X1 port map( A1 => DATA2(5), A2 => DATA1(5), B1 => n2600, B2 =>
                           n2773, ZN => n2564);
   U771 : AOI22_X1 port map( A1 => n2449, A2 => dataout_mul_5_port, B1 => n2438
                           , B2 => n2564, ZN => n1422);
   U772 : OAI22_X1 port map( A1 => n1969, A2 => n1389, B1 => n2461, B2 => n1388
                           , ZN => n1419);
   U773 : AOI22_X1 port map( A1 => n1389, A2 => n2466, B1 => n1388, B2 => n2004
                           , ZN => n1390);
   U774 : INV_X1 port map( A => n1390, ZN => n1417);
   U775 : OAI22_X1 port map( A1 => n1448, A2 => n2147, B1 => n1995, B2 => 
                           n2537_port, ZN => n1412);
   U776 : INV_X1 port map( A => n1978, ZN => n1434);
   U777 : NOR2_X1 port map( A1 => n1392, A2 => n1391, ZN => n1395);
   U778 : NAND2_X1 port map( A1 => DATA1(9), A2 => n1829, ZN => n1394);
   U779 : NAND2_X1 port map( A1 => n2039, A2 => n3096, ZN => n1674);
   U780 : NAND4_X1 port map( A1 => n1395, A2 => n1394, A3 => n1674, A4 => n1393
                           , ZN => n1470);
   U781 : AOI222_X1 port map( A1 => n1396, A2 => n2480, B1 => n1470, B2 => 
                           n2483, C1 => n1433, C2 => n1626, ZN => n2215);
   U782 : OAI22_X1 port map( A1 => n2213, A2 => n2215, B1 => n1471, B2 => n2487
                           , ZN => n1399);
   U783 : OAI22_X1 port map( A1 => n1631, A2 => n1397, B1 => n1435, B2 => n2491
                           , ZN => n1398);
   U784 : AOI211_X1 port map( C1 => n2494, C2 => n1434, A => n1399, B => n1398,
                           ZN => n2220);
   U785 : OAI22_X1 port map( A1 => n1474, A2 => n2497, B1 => n2220, B2 => n2499
                           , ZN => n1402);
   U786 : OAI22_X1 port map( A1 => n2501, A2 => n1400, B1 => n1982, B2 => n1779
                           , ZN => n1401);
   U787 : AOI211_X1 port map( C1 => n2373, C2 => n1403, A => n1402, B => n1401,
                           ZN => n1478);
   U788 : OAI222_X1 port map( A1 => n2510, A2 => n1443, B1 => n2508, B2 => 
                           n1478, C1 => n1404, C2 => n2512, ZN => n2225);
   U789 : AOI22_X1 port map( A1 => n2388, A2 => n1405, B1 => n2391, B2 => n2225
                           , ZN => n1408);
   U790 : AOI22_X1 port map( A1 => n2518_port, A2 => n1479, B1 => n2521_port, 
                           B2 => n1406, ZN => n1407);
   U791 : OAI211_X1 port map( C1 => n1482, C2 => n2268, A => n1408, B => n1407,
                           ZN => n2229);
   U792 : INV_X1 port map( A => n2229, ZN => n1410);
   U793 : OAI22_X1 port map( A1 => n1410, A2 => n2420, B1 => n1409, B2 => n1994
                           , ZN => n1411);
   U794 : AOI211_X1 port map( C1 => n2528_port, C2 => n1484, A => n1412, B => 
                           n1411, ZN => n1487);
   U795 : OAI222_X1 port map( A1 => n2100, A2 => n1452, B1 => n2113, B2 => 
                           n1487, C1 => n1413, C2 => n1996, ZN => n2236);
   U796 : INV_X1 port map( A => n2236, ZN => n1489);
   U797 : NOR2_X1 port map( A1 => n1414, A2 => n2775, ZN => n1826);
   U798 : AOI21_X1 port map( B1 => DATA2(4), B2 => n1415, A => n1826, ZN => 
                           n2548_port);
   U799 : INV_X1 port map( A => n2548_port, ZN => n1948);
   U800 : NOR3_X1 port map( A1 => n1489, A2 => n2455, A3 => n1948, ZN => n1416)
                           ;
   U801 : AOI221_X1 port map( B1 => n1420, B2 => n1419, C1 => n1418, C2 => 
                           n1417, A => n1416, ZN => n1421);
   U802 : NAND3_X1 port map( A1 => n1423, A2 => n1422, A3 => n1421, ZN => 
                           OUTALU(5));
   U803 : AOI22_X1 port map( A1 => n2466, A2 => n1454, B1 => n2004, B2 => n1453
                           , ZN => n1460);
   U804 : NOR3_X1 port map( A1 => n1424, A2 => n2083, A3 => n2427, ZN => n1427)
                           ;
   U805 : AOI22_X1 port map( A1 => DATA2(4), A2 => n2660, B1 => DATA1(4), B2 =>
                           n2774, ZN => n2597);
   U806 : AOI21_X1 port map( B1 => DATA1(4), B2 => n2412, A => n2410, ZN => 
                           n1425);
   U807 : OAI22_X1 port map( A1 => n2597, A2 => n2462, B1 => n1425, B2 => n2774
                           , ZN => n1426);
   U808 : AOI211_X1 port map( C1 => dataout_mul_4_port, C2 => n2449, A => n1427
                           , B => n1426, ZN => n1458);
   U809 : NOR2_X1 port map( A1 => n1826, A2 => n2548_port, ZN => n2235);
   U810 : INV_X1 port map( A => n2235, ZN => n2555);
   U811 : INV_X1 port map( A => n2537_port, ZN => n2431);
   U812 : INV_X1 port map( A => n2220, ZN => n1442);
   U813 : OAI211_X1 port map( C1 => n1548, C2 => n2609, A => n1429, B => n1428,
                           ZN => n1430);
   U814 : AOI211_X1 port map( C1 => DATA1(7), C2 => n2039, A => n1431, B => 
                           n1430, ZN => n1432);
   U815 : INV_X1 port map( A => n1432, ZN => n1976);
   U816 : AOI222_X1 port map( A1 => n2211, A2 => n1976, B1 => n1626, B2 => 
                           n1470, C1 => n2480, C2 => n1433, ZN => n2488);
   U817 : INV_X1 port map( A => n2488, ZN => n2218);
   U818 : AOI22_X1 port map( A1 => n2160, A2 => n1434, B1 => n1651, B2 => n2218
                           , ZN => n1438);
   U819 : OAI22_X1 port map( A1 => n1977, A2 => n2215, B1 => n2489, B2 => n1435
                           , ZN => n1436);
   U820 : INV_X1 port map( A => n1436, ZN => n1437);
   U821 : OAI211_X1 port map( C1 => n1471, C2 => n2491, A => n1438, B => n1437,
                           ZN => n1477);
   U822 : INV_X1 port map( A => n1477, ZN => n2500);
   U823 : OAI22_X1 port map( A1 => n2499, A2 => n2500, B1 => n2497, B2 => n1982
                           , ZN => n1441);
   U824 : OAI22_X1 port map( A1 => n2503, A2 => n1474, B1 => n2501, B2 => n1439
                           , ZN => n1440);
   U825 : AOI211_X1 port map( C1 => n1442, C2 => n2384, A => n1441, B => n1440,
                           ZN => n1986);
   U826 : OAI222_X1 port map( A1 => n1443, A2 => n2512, B1 => n1478, B2 => 
                           n2510, C1 => n1986, C2 => n2508, ZN => n2520_port);
   U827 : INV_X1 port map( A => n2520_port, ZN => n1444);
   U828 : INV_X1 port map( A => n1479, ZN => n1989);
   U829 : OAI22_X1 port map( A1 => n2323, A2 => n1444, B1 => n1989, B2 => n2268
                           , ZN => n1447);
   U830 : OAI22_X1 port map( A1 => n1990, A2 => n1445, B1 => n1482, B2 => 
                           n2525_port, ZN => n1446);
   U831 : AOI211_X1 port map( C1 => n2518_port, C2 => n2225, A => n1447, B => 
                           n1446, ZN => n1991);
   U832 : OAI22_X1 port map( A1 => n1995, A2 => n2153, B1 => n1991, B2 => n2420
                           , ZN => n1451);
   U833 : OAI22_X1 port map( A1 => n1449, A2 => n2147, B1 => n1448, B2 => n1994
                           , ZN => n1450);
   U834 : AOI211_X1 port map( C1 => n2431, C2 => n2229, A => n1451, B => n1450,
                           ZN => n1997);
   U835 : OAI222_X1 port map( A1 => n2100, A2 => n1487, B1 => n2113, B2 => 
                           n1997, C1 => n1452, C2 => n1996, ZN => n2551);
   U836 : INV_X1 port map( A => n2551, ZN => n1488);
   U837 : OAI22_X1 port map( A1 => n1489, A2 => n2555, B1 => n1488, B2 => n1948
                           , ZN => n1456);
   U838 : OAI22_X1 port map( A1 => n1454, A2 => n1969, B1 => n1453, B2 => n2461
                           , ZN => n1455);
   U839 : AOI22_X1 port map( A1 => n2736, A2 => n1456, B1 => n1459, B2 => n1455
                           , ZN => n1457);
   U840 : OAI211_X1 port map( C1 => n1460, C2 => n1459, A => n1458, B => n1457,
                           ZN => OUTALU(4));
   U841 : NOR2_X1 port map( A1 => n2474, A2 => n1463, ZN => n1466);
   U842 : NOR2_X1 port map( A1 => n1968, A2 => n2658, ZN => n2208);
   U843 : AOI211_X1 port map( C1 => DATA1(0), C2 => n2039, A => n1466, B => 
                           n2208, ZN => n1461);
   U844 : OAI21_X1 port map( B1 => n2025, B2 => n2651, A => n1461, ZN => n1462)
                           ;
   U845 : AOI22_X1 port map( A1 => DATA2(3), A2 => DATA1(3), B1 => n1463, B2 =>
                           n2775, ZN => n2570);
   U846 : AOI22_X1 port map( A1 => n2441, A2 => n1462, B1 => n2438, B2 => n2570
                           , ZN => n1499);
   U847 : OAI21_X1 port map( B1 => n1463, B2 => n2458, A => n2437, ZN => n1464)
                           ;
   U848 : AOI22_X1 port map( A1 => DATA2(3), A2 => n1464, B1 => n2354, B2 => 
                           dataout_mul_3_port, ZN => n1498);
   U849 : NAND2_X1 port map( A1 => n1826, A2 => n1465, ZN => n2239);
   U850 : AOI211_X1 port map( C1 => DATA1(6), C2 => n1830, A => n1467, B => 
                           n1466, ZN => n1469);
   U851 : NAND2_X1 port map( A1 => DATA1(7), A2 => n2477, ZN => n1468);
   U852 : OAI211_X1 port map( C1 => n2025, C2 => n2600, A => n1469, B => n1468,
                           ZN => n2212);
   U853 : AOI222_X1 port map( A1 => n1470, A2 => n2480, B1 => n2212, B2 => 
                           n2483, C1 => n1976, C2 => n1533, ZN => n2490);
   U854 : OAI22_X1 port map( A1 => n2213, A2 => n2490, B1 => n2215, B2 => n2487
                           , ZN => n1473);
   U855 : OAI22_X1 port map( A1 => n1631, A2 => n1471, B1 => n1978, B2 => n2491
                           , ZN => n1472);
   U856 : AOI211_X1 port map( C1 => n2494, C2 => n2218, A => n1473, B => n1472,
                           ZN => n2502);
   U857 : OAI22_X1 port map( A1 => n2220, A2 => n2497, B1 => n2502, B2 => n2499
                           , ZN => n1476);
   U858 : OAI22_X1 port map( A1 => n2501, A2 => n1474, B1 => n1982, B2 => n2503
                           , ZN => n1475);
   U859 : AOI211_X1 port map( C1 => n2506, C2 => n1477, A => n1476, B => n1475,
                           ZN => n2224);
   U860 : OAI222_X1 port map( A1 => n2510, A2 => n1986, B1 => n2508, B2 => 
                           n2224, C1 => n1478, C2 => n2512, ZN => n2206);
   U861 : AOI22_X1 port map( A1 => n2518_port, A2 => n2520_port, B1 => n2391, 
                           B2 => n2206, ZN => n1481);
   U862 : AOI22_X1 port map( A1 => n2514, A2 => n2225, B1 => n2388, B2 => n1479
                           , ZN => n1480);
   U863 : OAI211_X1 port map( C1 => n1990, C2 => n1482, A => n1481, B => n1480,
                           ZN => n2531_port);
   U864 : AOI22_X1 port map( A1 => n2526_port, A2 => n2531_port, B1 => 
                           n2528_port, B2 => n2229, ZN => n1486);
   U865 : INV_X1 port map( A => n2147, ZN => n2530_port);
   U866 : AOI22_X1 port map( A1 => n2532_port, A2 => n1484, B1 => n2530_port, 
                           B2 => n1483, ZN => n1485);
   U867 : OAI211_X1 port map( C1 => n1991, C2 => n2537_port, A => n1486, B => 
                           n1485, ZN => n2233);
   U868 : INV_X1 port map( A => n2233, ZN => n2000);
   U869 : OAI222_X1 port map( A1 => n2100, A2 => n1997, B1 => n1999, B2 => 
                           n2000, C1 => n1487, C2 => n1996, ZN => n2549);
   U870 : INV_X1 port map( A => n2549, ZN => n2240);
   U871 : OAI222_X1 port map( A1 => n2239, A2 => n1489, B1 => n2555, B2 => 
                           n1488, C1 => n1948, C2 => n2240, ZN => n1492);
   U872 : XOR2_X1 port map( A => n1495, B => n1490, Z => n1491);
   U873 : AOI22_X1 port map( A1 => n2736, A2 => n1492, B1 => n2466, B2 => n1491
                           , ZN => n1497);
   U874 : OAI211_X1 port map( C1 => n1495, C2 => n1494, A => n2004, B => n1493,
                           ZN => n1496);
   U875 : NAND4_X1 port map( A1 => n1499, A2 => n1498, A3 => n1497, A4 => n1496
                           , ZN => OUTALU(3));
   U876 : OAI211_X1 port map( C1 => n1710, C2 => n2578, A => n1501, B => n1500,
                           ZN => n1502);
   U877 : AOI211_X1 port map( C1 => DATA1(18), C2 => n2205, A => n1503, B => 
                           n1502, ZN => n1504);
   U878 : INV_X1 port map( A => n1504, ZN => n1535);
   U879 : OAI211_X1 port map( C1 => n1710, C2 => n2649, A => n1506, B => n1505,
                           ZN => n1507);
   U880 : AOI211_X1 port map( C1 => DATA1(17), C2 => n2205, A => n1508, B => 
                           n1507, ZN => n1509);
   U881 : INV_X1 port map( A => n1509, ZN => n1523);
   U882 : INV_X1 port map( A => n2397, ZN => n2681);
   U883 : OAI211_X1 port map( C1 => n1548, C2 => n2681, A => n1511, B => n1510,
                           ZN => n1512);
   U884 : AOI211_X1 port map( C1 => DATA1(16), C2 => n2205, A => n1513, B => 
                           n1512, ZN => n1514);
   U885 : INV_X1 port map( A => n1514, ZN => n1603);
   U886 : AOI222_X1 port map( A1 => n2211, A2 => n1535, B1 => n1626, B2 => 
                           n1523, C1 => n2480, C2 => n1603, ZN => n1647);
   U887 : INV_X1 port map( A => n1647, ZN => n1668);
   U888 : AOI22_X1 port map( A1 => DATA1(14), A2 => n2242, B1 => n2678, B2 => 
                           n2477, ZN => n1518);
   U889 : NAND4_X1 port map( A1 => n1518, A2 => n1517, A3 => n1516, A4 => n1515
                           , ZN => n1646);
   U890 : AOI222_X1 port map( A1 => n1646, A2 => n1975, B1 => n1523, B2 => 
                           n2483, C1 => n1603, C2 => n1533, ZN => n1679);
   U891 : AOI22_X1 port map( A1 => DATA1(16), A2 => n1830, B1 => n3098, B2 => 
                           n1829, ZN => n1522);
   U892 : NAND4_X1 port map( A1 => n1522, A2 => n1521, A3 => n1520, A4 => n1519
                           , ZN => n1534);
   U893 : AOI222_X1 port map( A1 => n1523, A2 => n2480, B1 => n1534, B2 => 
                           n2483, C1 => n1535, C2 => n1626, ZN => n1604);
   U894 : OAI22_X1 port map( A1 => n1631, A2 => n1679, B1 => n1604, B2 => n2487
                           , ZN => n1537);
   U895 : AOI22_X1 port map( A1 => DATA1(18), A2 => n1830, B1 => DATA1(17), B2 
                           => n2477, ZN => n1528);
   U896 : INV_X1 port map( A => n1524, ZN => n1525);
   U897 : NAND4_X1 port map( A1 => n1528, A2 => n1527, A3 => n1526, A4 => n1525
                           , ZN => n1560);
   U898 : AOI22_X1 port map( A1 => n1830, A2 => DATA1(17), B1 => n2315, B2 => 
                           n1829, ZN => n1532);
   U899 : NAND4_X1 port map( A1 => n1532, A2 => n1531, A3 => n1530, A4 => n1529
                           , ZN => n1558);
   U900 : AOI222_X1 port map( A1 => n1534, A2 => n1975, B1 => n1560, B2 => 
                           n2483, C1 => n1558, C2 => n1533, ZN => n1573);
   U901 : AOI222_X1 port map( A1 => n1535, A2 => n1975, B1 => n1558, B2 => 
                           n2483, C1 => n1534, C2 => n1626, ZN => n1598);
   U902 : OAI22_X1 port map( A1 => n1573, A2 => n2213, B1 => n1598, B2 => n2214
                           , ZN => n1536);
   U903 : AOI211_X1 port map( C1 => n1790, C2 => n1668, A => n1537, B => n1536,
                           ZN => n1682);
   U904 : AOI22_X1 port map( A1 => n1830, A2 => DATA1(20), B1 => n2256, B2 => 
                           n1829, ZN => n1541);
   U905 : NAND4_X1 port map( A1 => n1541, A2 => n1540, A3 => n1539, A4 => n1538
                           , ZN => n1551);
   U906 : AOI22_X1 port map( A1 => n1830, A2 => DATA1(19), B1 => n2284, B2 => 
                           n1829, ZN => n1545);
   U907 : NAND4_X1 port map( A1 => n1545, A2 => n1544, A3 => n1543, A4 => n1542
                           , ZN => n1559);
   U908 : AOI222_X1 port map( A1 => n1560, A2 => n1975, B1 => n1551, B2 => 
                           n2483, C1 => n1559, C2 => n1626, ZN => n1563);
   U909 : OAI211_X1 port map( C1 => n1548, C2 => n2701, A => n1547, B => n1546,
                           ZN => n1549);
   U910 : AOI211_X1 port map( C1 => n1145, C2 => DATA1(24), A => n1550, B => 
                           n1549, ZN => n1580);
   U911 : INV_X1 port map( A => n1551, ZN => n1557);
   U912 : INV_X1 port map( A => n1559, ZN => n1552);
   U913 : OAI222_X1 port map( A1 => n1174, A2 => n1580, B1 => n1754, B2 => 
                           n1557, C1 => n1752, C2 => n1552, ZN => n1615);
   U914 : OAI211_X1 port map( C1 => n1710, C2 => n2700, A => n1554, B => n1553,
                           ZN => n1555);
   U915 : AOI211_X1 port map( C1 => n1145, C2 => DATA1(25), A => n1556, B => 
                           n1555, ZN => n1590);
   U916 : OAI222_X1 port map( A1 => n1174, A2 => n1590, B1 => n1754, B2 => 
                           n1580, C1 => n1694, C2 => n1557, ZN => n1591);
   U917 : AOI22_X1 port map( A1 => n2494, A2 => n1615, B1 => n2156, B2 => n1591
                           , ZN => n1562);
   U918 : AOI222_X1 port map( A1 => n1626, A2 => n1560, B1 => n2483, B2 => 
                           n1559, C1 => n2480, C2 => n1558, ZN => n1569);
   U919 : INV_X1 port map( A => n1569, ZN => n1581);
   U920 : INV_X1 port map( A => n1573, ZN => n1566);
   U921 : AOI22_X1 port map( A1 => n1790, A2 => n1581, B1 => n1843, B2 => n1566
                           , ZN => n1561);
   U922 : OAI211_X1 port map( C1 => n1563, C2 => n2487, A => n1562, B => n1561,
                           ZN => n1618);
   U923 : INV_X1 port map( A => n1563, ZN => n1592);
   U924 : INV_X1 port map( A => n1604, ZN => n1650);
   U925 : AOI22_X1 port map( A1 => n1592, A2 => n1651, B1 => n1843, B2 => n1650
                           , ZN => n1565);
   U926 : INV_X1 port map( A => n1598, ZN => n1570);
   U927 : AOI22_X1 port map( A1 => n1790, A2 => n1570, B1 => n2494, B2 => n1581
                           , ZN => n1564);
   U928 : OAI211_X1 port map( C1 => n1573, C2 => n2487, A => n1565, B => n1564,
                           ZN => n1652);
   U929 : AOI22_X1 port map( A1 => n2442, A2 => n1618, B1 => n2383, B2 => n1652
                           , ZN => n1575);
   U930 : AOI22_X1 port map( A1 => n2494, A2 => n1592, B1 => n2156, B2 => n1615
                           , ZN => n1568);
   U931 : AOI22_X1 port map( A1 => n2219, A2 => n1566, B1 => n1925, B2 => n1570
                           , ZN => n1567);
   U932 : OAI211_X1 port map( C1 => n1569, C2 => n2487, A => n1568, B => n1567,
                           ZN => n1619);
   U933 : AOI22_X1 port map( A1 => n2160, A2 => n1570, B1 => n1581, B2 => n1651
                           , ZN => n1572);
   U934 : AOI22_X1 port map( A1 => n1790, A2 => n1650, B1 => n1843, B2 => n1668
                           , ZN => n1571);
   U935 : OAI211_X1 port map( C1 => n1573, C2 => n2214, A => n1572, B => n1571,
                           ZN => n1672);
   U936 : AOI22_X1 port map( A1 => n2506, A2 => n1619, B1 => n1932, B2 => n1672
                           , ZN => n1574);
   U937 : OAI211_X1 port map( C1 => n2501, C2 => n1682, A => n1575, B => n1574,
                           ZN => n1657);
   U938 : INV_X1 port map( A => n1618, ZN => n1636);
   U939 : INV_X1 port map( A => n1591, ZN => n1630);
   U940 : OAI211_X1 port map( C1 => n1710, C2 => n2161, A => n1577, B => n1576,
                           ZN => n1578);
   U941 : AOI211_X1 port map( C1 => n1145, C2 => DATA1(26), A => n1579, B => 
                           n1578, ZN => n1614);
   U942 : OAI222_X1 port map( A1 => n2083, A2 => n1614, B1 => n2081, B2 => 
                           n1590, C1 => n1694, C2 => n1580, ZN => n1716);
   U943 : AOI22_X1 port map( A1 => n2219, A2 => n1592, B1 => n2156, B2 => n1716
                           , ZN => n1583);
   U944 : AOI22_X1 port map( A1 => n2160, A2 => n1615, B1 => n1925, B2 => n1581
                           , ZN => n1582);
   U945 : OAI211_X1 port map( C1 => n1630, C2 => n2214, A => n1583, B => n1582,
                           ZN => n1719);
   U946 : AOI22_X1 port map( A1 => n2442, A2 => n1719, B1 => n2373, B2 => n1652
                           , ZN => n1585);
   U947 : AOI22_X1 port map( A1 => n2383, A2 => n1619, B1 => n1931, B2 => n1672
                           , ZN => n1584);
   U948 : OAI211_X1 port map( C1 => n1636, C2 => n1779, A => n1585, B => n1584,
                           ZN => n1640);
   U949 : INV_X1 port map( A => n1719, ZN => n1635);
   U950 : INV_X1 port map( A => n1716, ZN => n1595);
   U951 : OAI211_X1 port map( C1 => n1710, C2 => n2128, A => n1587, B => n1586,
                           ZN => n1588);
   U952 : AOI211_X1 port map( C1 => n1145, C2 => DATA1(27), A => n1589, B => 
                           n1588, ZN => n1622);
   U953 : OAI222_X1 port map( A1 => n1174, A2 => n1622, B1 => n1754, B2 => 
                           n1614, C1 => n1752, C2 => n1590, ZN => n1842);
   U954 : AOI22_X1 port map( A1 => n2160, A2 => n1591, B1 => n1651, B2 => n1842
                           , ZN => n1594);
   U955 : AOI22_X1 port map( A1 => n1790, A2 => n1615, B1 => n1592, B2 => n1925
                           , ZN => n1593);
   U956 : OAI211_X1 port map( C1 => n1595, C2 => n1977, A => n1594, B => n1593,
                           ZN => n1847);
   U957 : AOI22_X1 port map( A1 => n2442, A2 => n1847, B1 => n2383, B2 => n1618
                           , ZN => n1597);
   U958 : AOI22_X1 port map( A1 => n1932, A2 => n1619, B1 => n1931, B2 => n1652
                           , ZN => n1596);
   U959 : OAI211_X1 port map( C1 => n1635, C2 => n1779, A => n1597, B => n1596,
                           ZN => n1641);
   U960 : AOI222_X1 port map( A1 => n1657, A2 => n1938, B1 => n1640, B2 => 
                           n2321, C1 => n1641, C2 => n2357, ZN => n1858);
   U961 : INV_X1 port map( A => n1619, ZN => n1609);
   U962 : INV_X1 port map( A => n1682, ZN => n1653);
   U963 : AOI22_X1 port map( A1 => n1652, A2 => n2506, B1 => n1653, B2 => n1932
                           , ZN => n1608);
   U964 : OAI22_X1 port map( A1 => n2213, A2 => n1598, B1 => n1679, B2 => n2491
                           , ZN => n1606);
   U965 : AOI22_X1 port map( A1 => DATA1(14), A2 => n2205, B1 => DATA1(10), B2 
                           => n1829, ZN => n1602);
   U966 : NAND4_X1 port map( A1 => n1602, A2 => n1601, A3 => n1600, A4 => n1599
                           , ZN => n1665);
   U967 : AOI222_X1 port map( A1 => n1665, A2 => n1975, B1 => n1603, B2 => 
                           n2483, C1 => n1646, C2 => n1626, ZN => n1699);
   U968 : OAI22_X1 port map( A1 => n1631, A2 => n1699, B1 => n1604, B2 => n1977
                           , ZN => n1605);
   U969 : AOI211_X1 port map( C1 => n2127, C2 => n1668, A => n1606, B => n1605,
                           ZN => n1669);
   U970 : INV_X1 port map( A => n1669, ZN => n1701);
   U971 : AOI22_X1 port map( A1 => n1848, A2 => n1701, B1 => n1672, B2 => n2383
                           , ZN => n1607);
   U972 : OAI211_X1 port map( C1 => n2499, C2 => n1609, A => n1608, B => n1607,
                           ZN => n1704);
   U973 : AOI222_X1 port map( A1 => n2321, A2 => n1657, B1 => n1936, B2 => 
                           n1640, C1 => n1704, C2 => n1938, ZN => n1726);
   U974 : INV_X1 port map( A => n1726, ZN => n1732);
   U975 : INV_X1 port map( A => n1847, ZN => n1634);
   U976 : AOI22_X1 port map( A1 => DATA1(25), A2 => n1830, B1 => DATA1(24), B2 
                           => n1829, ZN => n1612);
   U977 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(28), ZN => n2042);
   U978 : NAND4_X1 port map( A1 => n1612, A2 => n1611, A3 => n1610, A4 => n2042
                           , ZN => n1714);
   U979 : INV_X1 port map( A => n1714, ZN => n1613);
   U980 : OAI222_X1 port map( A1 => n1614, A2 => n1694, B1 => n1613, B2 => 
                           n2083, C1 => n1622, C2 => n1754, ZN => n1629);
   U981 : AOI22_X1 port map( A1 => n2156, A2 => n1629, B1 => n1716, B2 => n2160
                           , ZN => n1617);
   U982 : AOI22_X1 port map( A1 => n1843, A2 => n1615, B1 => n1842, B2 => n2494
                           , ZN => n1616);
   U983 : OAI211_X1 port map( C1 => n2491, C2 => n1630, A => n1617, B => n1616,
                           ZN => n1852);
   U984 : AOI22_X1 port map( A1 => n1719, A2 => n2383, B1 => n1852, B2 => n2442
                           , ZN => n1621);
   U985 : AOI22_X1 port map( A1 => n1848, A2 => n1619, B1 => n1618, B2 => n2373
                           , ZN => n1620);
   U986 : OAI211_X1 port map( C1 => n1779, C2 => n1634, A => n1621, B => n1620,
                           ZN => n1723);
   U987 : INV_X1 port map( A => n1622, ZN => n1627);
   U988 : AOI22_X1 port map( A1 => DATA1(26), A2 => n1830, B1 => DATA1(25), B2 
                           => n1829, ZN => n1625);
   U989 : NAND2_X1 port map( A1 => n1145, A2 => DATA1(29), ZN => n2023);
   U990 : NAND4_X1 port map( A1 => n1625, A2 => n1624, A3 => n1623, A4 => n2023
                           , ZN => n1835);
   U991 : AOI222_X1 port map( A1 => n1627, A2 => n1975, B1 => n1835, B2 => 
                           n2483, C1 => n1714, C2 => n1626, ZN => n1836);
   U992 : INV_X1 port map( A => n1842, ZN => n1628);
   U993 : OAI22_X1 port map( A1 => n2213, A2 => n1836, B1 => n1628, B2 => n2487
                           , ZN => n1633);
   U994 : INV_X1 port map( A => n1629, ZN => n1839);
   U995 : OAI22_X1 port map( A1 => n1631, A2 => n1630, B1 => n1839, B2 => n2214
                           , ZN => n1632);
   U996 : AOI211_X1 port map( C1 => n2219, C2 => n1716, A => n1633, B => n1632,
                           ZN => n1845);
   U997 : OAI22_X1 port map( A1 => n1634, A2 => n2497, B1 => n1845, B2 => n2499
                           , ZN => n1638);
   U998 : OAI22_X1 port map( A1 => n1636, A2 => n2501, B1 => n1635, B2 => n2503
                           , ZN => n1637);
   U999 : AOI211_X1 port map( C1 => n2384, C2 => n1852, A => n1638, B => n1637,
                           ZN => n1853);
   U1000 : INV_X1 port map( A => n1853, ZN => n1722);
   U1001 : AOI222_X1 port map( A1 => n2321, A2 => n1723, B1 => n1936, B2 => 
                           n1722, C1 => n1641, C2 => n1938, ZN => n1639);
   U1002 : INV_X1 port map( A => n1639, ZN => n1857);
   U1003 : AOI22_X1 port map( A1 => n2388, A2 => n1732, B1 => n2391, B2 => 
                           n1857, ZN => n1660);
   U1004 : AOI222_X1 port map( A1 => n2321, A2 => n1641, B1 => n1936, B2 => 
                           n1723, C1 => n1640, C2 => n1938, ZN => n1859);
   U1005 : INV_X1 port map( A => n1672, ZN => n1656);
   U1006 : AOI22_X1 port map( A1 => DATA1(13), A2 => n2205, B1 => n3097, B2 => 
                           n1829, ZN => n1645);
   U1007 : NAND4_X1 port map( A1 => n1645, A2 => n1644, A3 => n1643, A4 => 
                           n1642, ZN => n1678);
   U1008 : AOI222_X1 port map( A1 => n1678, A2 => n1975, B1 => n1646, B2 => 
                           n2211, C1 => n1665, C2 => n1626, ZN => n1739);
   U1009 : OAI22_X1 port map( A1 => n2489, A2 => n1739, B1 => n1679, B2 => 
                           n2487, ZN => n1649);
   U1010 : OAI22_X1 port map( A1 => n1647, A2 => n1977, B1 => n1699, B2 => 
                           n2491, ZN => n1648);
   U1011 : AOI211_X1 port map( C1 => n1651, C2 => n1650, A => n1649, B => n1648
                           , ZN => n1741);
   U1012 : INV_X1 port map( A => n1741, ZN => n1700);
   U1013 : AOI22_X1 port map( A1 => n1848, A2 => n1700, B1 => n1652, B2 => 
                           n2442, ZN => n1655);
   U1014 : AOI22_X1 port map( A1 => n1653, A2 => n2383, B1 => n1701, B2 => 
                           n2373, ZN => n1654);
   U1015 : OAI211_X1 port map( C1 => n1779, C2 => n1656, A => n1655, B => n1654
                           , ZN => n1705);
   U1016 : AOI222_X1 port map( A1 => n2321, A2 => n1704, B1 => n1936, B2 => 
                           n1657, C1 => n1705, C2 => n1938, ZN => n1746);
   U1017 : OAI22_X1 port map( A1 => n2293, A2 => n1859, B1 => n1990, B2 => 
                           n1746, ZN => n1658);
   U1018 : INV_X1 port map( A => n1658, ZN => n1659);
   U1019 : OAI211_X1 port map( C1 => n1858, C2 => n2268, A => n1660, B => n1659
                           , ZN => n1864);
   U1020 : OAI22_X1 port map( A1 => n1682, A2 => n1779, B1 => n1741, B2 => 
                           n2503, ZN => n1671);
   U1021 : AOI22_X1 port map( A1 => n2397, A2 => n2205, B1 => n3096, B2 => 
                           n1829, ZN => n1664);
   U1022 : NAND4_X1 port map( A1 => n1664, A2 => n1663, A3 => n1662, A4 => 
                           n1661, ZN => n1687);
   U1023 : AOI222_X1 port map( A1 => n1687, A2 => n1975, B1 => n1665, B2 => 
                           n2211, C1 => n1678, C2 => n1626, ZN => n1758);
   U1024 : OAI22_X1 port map( A1 => n2489, A2 => n1758, B1 => n1699, B2 => 
                           n2487, ZN => n1667);
   U1025 : OAI22_X1 port map( A1 => n1679, A2 => n2214, B1 => n1739, B2 => 
                           n2491, ZN => n1666);
   U1026 : AOI211_X1 port map( C1 => n2156, C2 => n1668, A => n1667, B => n1666
                           , ZN => n1761);
   U1027 : OAI22_X1 port map( A1 => n2501, A2 => n1761, B1 => n1669, B2 => 
                           n2497, ZN => n1670);
   U1028 : AOI211_X1 port map( C1 => n2385, C2 => n1672, A => n1671, B => n1670
                           , ZN => n1673);
   U1029 : INV_X1 port map( A => n1673, ZN => n1706);
   U1030 : INV_X1 port map( A => n1758, ZN => n1736);
   U1031 : AOI22_X1 port map( A1 => DATA1(11), A2 => n2205, B1 => DATA1(7), B2 
                           => n1829, ZN => n1677);
   U1032 : NAND4_X1 port map( A1 => n1677, A2 => n1676, A3 => n1675, A4 => 
                           n1674, ZN => n1688);
   U1033 : AOI222_X1 port map( A1 => n1688, A2 => n1975, B1 => n1678, B2 => 
                           n2483, C1 => n1687, C2 => n1626, ZN => n1686);
   U1034 : OAI22_X1 port map( A1 => n2489, A2 => n1686, B1 => n1739, B2 => 
                           n2487, ZN => n1681);
   U1035 : OAI22_X1 port map( A1 => n2213, A2 => n1679, B1 => n1699, B2 => 
                           n1977, ZN => n1680);
   U1036 : AOI211_X1 port map( C1 => n1790, C2 => n1736, A => n1681, B => n1680
                           , ZN => n1740);
   U1037 : OAI22_X1 port map( A1 => n2501, A2 => n1740, B1 => n1682, B2 => 
                           n2499, ZN => n1684);
   U1038 : OAI22_X1 port map( A1 => n1741, A2 => n2497, B1 => n1761, B2 => 
                           n2503, ZN => n1683);
   U1039 : AOI211_X1 port map( C1 => n2384, C2 => n1701, A => n1684, B => n1683
                           , ZN => n1685);
   U1040 : INV_X1 port map( A => n1685, ZN => n1745);
   U1041 : AOI222_X1 port map( A1 => n2321, A2 => n1706, B1 => n1936, B2 => 
                           n1705, C1 => n1745, C2 => n1938, ZN => n1763);
   U1042 : INV_X1 port map( A => n1763, ZN => n1808);
   U1043 : INV_X1 port map( A => n1686, ZN => n1774);
   U1044 : AOI22_X1 port map( A1 => n2160, A2 => n1736, B1 => n2219, B2 => 
                           n1774, ZN => n1698);
   U1045 : INV_X1 port map( A => n1739, ZN => n1696);
   U1046 : INV_X1 port map( A => n1687, ZN => n1695);
   U1047 : INV_X1 port map( A => n1688, ZN => n1735);
   U1048 : OAI211_X1 port map( C1 => n2667, C2 => n1691, A => n1690, B => n1689
                           , ZN => n1692);
   U1049 : AOI211_X1 port map( C1 => DATA1(6), C2 => n2477, A => n1693, B => 
                           n1692, ZN => n1755);
   U1050 : OAI222_X1 port map( A1 => n2083, A2 => n1695, B1 => n1754, B2 => 
                           n1735, C1 => n1694, C2 => n1755, ZN => n1773);
   U1051 : AOI22_X1 port map( A1 => n2494, A2 => n1696, B1 => n1925, B2 => 
                           n1773, ZN => n1697);
   U1052 : OAI211_X1 port map( C1 => n2485, C2 => n1699, A => n1698, B => n1697
                           , ZN => n1781);
   U1053 : AOI22_X1 port map( A1 => n2506, A2 => n1700, B1 => n1931, B2 => 
                           n1781, ZN => n1703);
   U1054 : INV_X1 port map( A => n1740, ZN => n1782);
   U1055 : AOI22_X1 port map( A1 => n2442, A2 => n1701, B1 => n1932, B2 => 
                           n1782, ZN => n1702);
   U1056 : OAI211_X1 port map( C1 => n1761, C2 => n2497, A => n1703, B => n1702
                           , ZN => n1762);
   U1057 : AOI222_X1 port map( A1 => n1762, A2 => n1938, B1 => n1745, B2 => 
                           n2321, C1 => n1706, C2 => n2357, ZN => n1805);
   U1058 : AOI222_X1 port map( A1 => n1706, A2 => n1938, B1 => n1705, B2 => 
                           n2321, C1 => n1704, C2 => n2357, ZN => n1764);
   U1059 : OAI22_X1 port map( A1 => n1990, A2 => n1805, B1 => n1764, B2 => 
                           n2268, ZN => n1708);
   U1060 : OAI22_X1 port map( A1 => n2323, A2 => n1726, B1 => n1746, B2 => 
                           n2293, ZN => n1707);
   U1061 : AOI211_X1 port map( C1 => n2388, C2 => n1808, A => n1708, B => n1707
                           , ZN => n1818);
   U1062 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(29), ZN => n2041);
   U1063 : OAI211_X1 port map( C1 => n1710, C2 => n2557, A => n1709, B => n2041
                           , ZN => n1711);
   U1064 : AOI211_X1 port map( C1 => n1145, C2 => DATA1(30), A => n1712, B => 
                           n1711, ZN => n1713);
   U1065 : INV_X1 port map( A => n1713, ZN => n1833);
   U1066 : AOI222_X1 port map( A1 => n2211, A2 => n1833, B1 => n1626, B2 => 
                           n1835, C1 => n2480, C2 => n1714, ZN => n1838);
   U1067 : OAI22_X1 port map( A1 => n2487, A2 => n1839, B1 => n2485, B2 => 
                           n1838, ZN => n1715);
   U1068 : INV_X1 port map( A => n1715, ZN => n1718);
   U1069 : AOI22_X1 port map( A1 => n2219, A2 => n1842, B1 => n1843, B2 => 
                           n1716, ZN => n1717);
   U1070 : OAI211_X1 port map( C1 => n1836, C2 => n1977, A => n1718, B => n1717
                           , ZN => n1846);
   U1071 : AOI22_X1 port map( A1 => n2442, A2 => n1846, B1 => n2383, B2 => 
                           n1852, ZN => n1721);
   U1072 : AOI22_X1 port map( A1 => n2373, A2 => n1847, B1 => n1931, B2 => 
                           n1719, ZN => n1720);
   U1073 : OAI211_X1 port map( C1 => n1845, C2 => n1779, A => n1721, B => n1720
                           , ZN => n1828);
   U1074 : AOI222_X1 port map( A1 => n1723, A2 => n1938, B1 => n1722, B2 => 
                           n2321, C1 => n1828, C2 => n2357, ZN => n1863);
   U1075 : OAI22_X1 port map( A1 => n1858, A2 => n2525_port, B1 => n2323, B2 =>
                           n1863, ZN => n1725);
   U1076 : OAI22_X1 port map( A1 => n1726, A2 => n1990, B1 => n1859, B2 => 
                           n2268, ZN => n1724);
   U1077 : AOI211_X1 port map( C1 => n2518_port, C2 => n1857, A => n1725, B => 
                           n1724, ZN => n1867);
   U1078 : OAI22_X1 port map( A1 => n1818, A2 => n1994, B1 => n1867, B2 => 
                           n2420, ZN => n1734);
   U1079 : INV_X1 port map( A => n1859, ZN => n1729);
   U1080 : OAI22_X1 port map( A1 => n1726, A2 => n2268, B1 => n1858, B2 => 
                           n2293, ZN => n1728);
   U1081 : OAI22_X1 port map( A1 => n1746, A2 => n2525_port, B1 => n1990, B2 =>
                           n1764, ZN => n1727);
   U1082 : AOI211_X1 port map( C1 => n2517_port, C2 => n1729, A => n1728, B => 
                           n1727, ZN => n1866);
   U1083 : OAI22_X1 port map( A1 => n1990, A2 => n1763, B1 => n1764, B2 => 
                           n2525_port, ZN => n1731);
   U1084 : OAI22_X1 port map( A1 => n2323, A2 => n1858, B1 => n1746, B2 => 
                           n2268, ZN => n1730);
   U1085 : AOI211_X1 port map( C1 => n2518_port, C2 => n1732, A => n1731, B => 
                           n1730, ZN => n1871);
   U1086 : OAI22_X1 port map( A1 => n1866, A2 => n2153, B1 => n1871, B2 => 
                           n2147, ZN => n1733);
   U1087 : AOI211_X1 port map( C1 => n2431, C2 => n1864, A => n1734, B => n1733
                           , ZN => n1827);
   U1088 : INV_X1 port map( A => n1871, ZN => n1769);
   U1089 : AOI22_X1 port map( A1 => n1769, A2 => n2528_port, B1 => n1864, B2 =>
                           n2526_port, ZN => n1750);
   U1090 : INV_X1 port map( A => n1805, ZN => n1789);
   U1091 : OAI222_X1 port map( A1 => n1174, A2 => n1735, B1 => n2081, B2 => 
                           n1755, C1 => n1752, C2 => n1753, ZN => n1770);
   U1092 : AOI22_X1 port map( A1 => n2160, A2 => n1774, B1 => n1925, B2 => 
                           n1770, ZN => n1738);
   U1093 : AOI22_X1 port map( A1 => n1790, A2 => n1773, B1 => n2494, B2 => 
                           n1736, ZN => n1737);
   U1094 : OAI211_X1 port map( C1 => n2485, C2 => n1739, A => n1738, B => n1737
                           , ZN => n1796);
   U1095 : INV_X1 port map( A => n1796, ZN => n1780);
   U1096 : OAI22_X1 port map( A1 => n1779, A2 => n1761, B1 => n2501, B2 => 
                           n1780, ZN => n1743);
   U1097 : OAI22_X1 port map( A1 => n2499, A2 => n1741, B1 => n2497, B2 => 
                           n1740, ZN => n1742);
   U1098 : AOI211_X1 port map( C1 => n1781, C2 => n1932, A => n1743, B => n1742
                           , ZN => n1744);
   U1099 : INV_X1 port map( A => n1744, ZN => n1785);
   U1100 : AOI222_X1 port map( A1 => n1785, A2 => n1938, B1 => n1762, B2 => 
                           n2321, C1 => n1745, C2 => n1936, ZN => n1804);
   U1101 : OAI22_X1 port map( A1 => n1990, A2 => n1804, B1 => n1763, B2 => 
                           n2268, ZN => n1748);
   U1102 : OAI22_X1 port map( A1 => n2323, A2 => n1746, B1 => n1764, B2 => 
                           n2293, ZN => n1747);
   U1103 : AOI211_X1 port map( C1 => n2388, C2 => n1789, A => n1748, B => n1747
                           , ZN => n1819);
   U1104 : INV_X1 port map( A => n1819, ZN => n1814);
   U1105 : INV_X1 port map( A => n1818, ZN => n1811);
   U1106 : AOI22_X1 port map( A1 => n1814, A2 => n2532_port, B1 => n1811, B2 =>
                           n2530_port, ZN => n1749);
   U1107 : OAI211_X1 port map( C1 => n2537_port, C2 => n1866, A => n1750, B => 
                           n1749, ZN => n1874);
   U1108 : INV_X1 port map( A => n1874, ZN => n1822);
   U1109 : OAI22_X1 port map( A1 => n1819, A2 => n2147, B1 => n1818, B2 => 
                           n2153, ZN => n1768);
   U1110 : INV_X1 port map( A => n1804, ZN => n1803);
   U1111 : AOI22_X1 port map( A1 => n2160, A2 => n1773, B1 => n2219, B2 => 
                           n1770, ZN => n1757);
   U1112 : OAI222_X1 port map( A1 => n2083, A2 => n1755, B1 => n1754, B2 => 
                           n1753, C1 => n1752, C2 => n1751, ZN => n1923);
   U1113 : AOI22_X1 port map( A1 => n2494, A2 => n1774, B1 => n1843, B2 => 
                           n1923, ZN => n1756);
   U1114 : OAI211_X1 port map( C1 => n2213, C2 => n1758, A => n1757, B => n1756
                           , ZN => n1795);
   U1115 : AOI22_X1 port map( A1 => n2506, A2 => n1782, B1 => n1931, B2 => 
                           n1795, ZN => n1760);
   U1116 : AOI22_X1 port map( A1 => n2383, A2 => n1781, B1 => n2373, B2 => 
                           n1796, ZN => n1759);
   U1117 : OAI211_X1 port map( C1 => n1761, C2 => n2499, A => n1760, B => n1759
                           , ZN => n1786);
   U1118 : AOI222_X1 port map( A1 => n1786, A2 => n1938, B1 => n1785, B2 => 
                           n2321, C1 => n1762, C2 => n1936, ZN => n1922);
   U1119 : OAI22_X1 port map( A1 => n1990, A2 => n1922, B1 => n1805, B2 => 
                           n2268, ZN => n1766);
   U1120 : OAI22_X1 port map( A1 => n2323, A2 => n1764, B1 => n1763, B2 => 
                           n2293, ZN => n1765);
   U1121 : AOI211_X1 port map( C1 => n2388, C2 => n1803, A => n1766, B => n1765
                           , ZN => n1813);
   U1122 : OAI22_X1 port map( A1 => n1813, A2 => n1994, B1 => n1866, B2 => 
                           n2420, ZN => n1767);
   U1123 : AOI211_X1 port map( C1 => n2431, C2 => n1769, A => n1768, B => n1767
                           , ZN => n1825);
   U1124 : OAI222_X1 port map( A1 => n2113, A2 => n1827, B1 => n2100, B2 => 
                           n1822, C1 => n1825, C2 => n1996, ZN => n1920);
   U1125 : INV_X1 port map( A => n1770, ZN => n1794);
   U1126 : AOI22_X1 port map( A1 => n2160, A2 => n1923, B1 => n2156, B2 => 
                           n1773, ZN => n1772);
   U1127 : AOI22_X1 port map( A1 => n2219, A2 => n1791, B1 => n1843, B2 => 
                           n1927, ZN => n1771);
   U1128 : OAI211_X1 port map( C1 => n1794, C2 => n2214, A => n1772, B => n1771
                           , ZN => n2386);
   U1129 : AOI22_X1 port map( A1 => n2383, A2 => n1795, B1 => n1931, B2 => 
                           n2386, ZN => n1778);
   U1130 : AOI22_X1 port map( A1 => n1790, A2 => n1923, B1 => n2494, B2 => 
                           n1773, ZN => n1776);
   U1131 : AOI22_X1 port map( A1 => n1843, A2 => n1791, B1 => n2156, B2 => 
                           n1774, ZN => n1775);
   U1132 : OAI211_X1 port map( C1 => n1794, C2 => n2487, A => n1776, B => n1775
                           , ZN => n2372);
   U1133 : AOI22_X1 port map( A1 => n2385, A2 => n1781, B1 => n2373, B2 => 
                           n2372, ZN => n1777);
   U1134 : OAI211_X1 port map( C1 => n1780, C2 => n1779, A => n1778, B => n1777
                           , ZN => n1937);
   U1135 : INV_X1 port map( A => n1795, ZN => n1935);
   U1136 : AOI22_X1 port map( A1 => n2383, A2 => n1796, B1 => n1931, B2 => 
                           n2372, ZN => n1784);
   U1137 : AOI22_X1 port map( A1 => n2385, A2 => n1782, B1 => n2384, B2 => 
                           n1781, ZN => n1783);
   U1138 : OAI211_X1 port map( C1 => n1935, C2 => n2503, A => n1784, B => n1783
                           , ZN => n1800);
   U1139 : AOI222_X1 port map( A1 => n1937, A2 => n1938, B1 => n1800, B2 => 
                           n2321, C1 => n1786, C2 => n1936, ZN => n2269);
   U1140 : OAI22_X1 port map( A1 => n1990, A2 => n2269, B1 => n1922, B2 => 
                           n2268, ZN => n1788);
   U1141 : AOI222_X1 port map( A1 => n1800, A2 => n1938, B1 => n1786, B2 => 
                           n2321, C1 => n1785, C2 => n1936, ZN => n2254);
   U1142 : OAI22_X1 port map( A1 => n1804, A2 => n2293, B1 => n2254, B2 => 
                           n2525_port, ZN => n1787);
   U1143 : AOI211_X1 port map( C1 => n2517_port, C2 => n1789, A => n1788, B => 
                           n1787, ZN => n2154);
   U1144 : INV_X1 port map( A => n2154, ZN => n1812);
   U1145 : INV_X1 port map( A => n2386, ZN => n1799);
   U1146 : AOI22_X1 port map( A1 => n1925, A2 => n1926, B1 => n1923, B2 => 
                           n2494, ZN => n1793);
   U1147 : AOI22_X1 port map( A1 => n1791, A2 => n2160, B1 => n1927, B2 => 
                           n1790, ZN => n1792);
   U1148 : OAI211_X1 port map( C1 => n2213, C2 => n1794, A => n1793, B => n1792
                           , ZN => n2409);
   U1149 : AOI22_X1 port map( A1 => n1848, A2 => n2409, B1 => n2372, B2 => 
                           n2383, ZN => n1798);
   U1150 : AOI22_X1 port map( A1 => n1796, A2 => n2442, B1 => n1795, B2 => 
                           n2384, ZN => n1797);
   U1151 : OAI211_X1 port map( C1 => n2503, C2 => n1799, A => n1798, B => n1797
                           , ZN => n2322);
   U1152 : AOI222_X1 port map( A1 => n2321, A2 => n1937, B1 => n1936, B2 => 
                           n1800, C1 => n2322, C2 => n1938, ZN => n2294);
   U1153 : OAI22_X1 port map( A1 => n2268, A2 => n2254, B1 => n1990, B2 => 
                           n2294, ZN => n1802);
   U1154 : OAI22_X1 port map( A1 => n2293, A2 => n1922, B1 => n2525_port, B2 =>
                           n2269, ZN => n1801);
   U1155 : AOI211_X1 port map( C1 => n2517_port, C2 => n1803, A => n1802, B => 
                           n1801, ZN => n2176);
   U1156 : OAI22_X1 port map( A1 => n2268, A2 => n1804, B1 => n1990, B2 => 
                           n2254, ZN => n1807);
   U1157 : OAI22_X1 port map( A1 => n2293, A2 => n1805, B1 => n2525_port, B2 =>
                           n1922, ZN => n1806);
   U1158 : AOI211_X1 port map( C1 => n2517_port, C2 => n1808, A => n1807, B => 
                           n1806, ZN => n2146);
   U1159 : OAI22_X1 port map( A1 => n1994, A2 => n2176, B1 => n2153, B2 => 
                           n2146, ZN => n1810);
   U1160 : OAI22_X1 port map( A1 => n2537_port, A2 => n1813, B1 => n2420, B2 =>
                           n1819, ZN => n1809);
   U1161 : AOI211_X1 port map( C1 => n1812, C2 => n2530_port, A => n1810, B => 
                           n1809, ZN => n2099);
   U1162 : AOI22_X1 port map( A1 => n2532_port, A2 => n1812, B1 => n2526_port, 
                           B2 => n1811, ZN => n1816);
   U1163 : INV_X1 port map( A => n1813, ZN => n1944);
   U1164 : AOI22_X1 port map( A1 => n2431, A2 => n1814, B1 => n2228, B2 => 
                           n1944, ZN => n1815);
   U1165 : OAI211_X1 port map( C1 => n2146, C2 => n2147, A => n1816, B => n1815
                           , ZN => n1817);
   U1166 : INV_X1 port map( A => n1817, ZN => n1945);
   U1167 : OAI22_X1 port map( A1 => n1994, A2 => n2146, B1 => n2537_port, B2 =>
                           n1818, ZN => n1821);
   U1168 : OAI22_X1 port map( A1 => n2153, A2 => n1819, B1 => n2420, B2 => 
                           n1871, ZN => n1820);
   U1169 : AOI211_X1 port map( C1 => n1944, C2 => n2530_port, A => n1821, B => 
                           n1820, ZN => n1824);
   U1170 : OAI222_X1 port map( A1 => n2099, A2 => n1996, B1 => n1945, B2 => 
                           n2100, C1 => n1824, C2 => n1999, ZN => n2063);
   U1171 : OAI222_X1 port map( A1 => n1824, A2 => n1996, B1 => n1825, B2 => 
                           n2100, C1 => n1822, C2 => n1999, ZN => n2014);
   U1172 : INV_X1 port map( A => n2239, ZN => n2546_port);
   U1173 : AOI22_X1 port map( A1 => n2063, A2 => n2552, B1 => n2014, B2 => 
                           n2546_port, ZN => n1823);
   U1174 : INV_X1 port map( A => n1823, ZN => n1878);
   U1175 : OAI222_X1 port map( A1 => n1945, A2 => n1996, B1 => n1825, B2 => 
                           n2113, C1 => n1824, C2 => n2100, ZN => n2036);
   U1176 : INV_X1 port map( A => n2036, ZN => n1876);
   U1177 : INV_X1 port map( A => n2552, ZN => n1917);
   U1178 : NAND3_X1 port map( A1 => DATA2(0), A2 => n1826, A3 => n1917, ZN => 
                           n1921);
   U1179 : INV_X1 port map( A => n1827, ZN => n1873);
   U1180 : INV_X1 port map( A => n1828, ZN => n1855);
   U1181 : AOI22_X1 port map( A1 => DATA1(28), A2 => n1830, B1 => DATA1(27), B2
                           => n1829, ZN => n1832);
   U1182 : NAND2_X1 port map( A1 => n2242, A2 => DATA1(30), ZN => n2024);
   U1183 : NAND2_X1 port map( A1 => n2205, A2 => DATA1(31), ZN => n1909);
   U1184 : NAND4_X1 port map( A1 => n1832, A2 => n1831, A3 => n2024, A4 => 
                           n1909, ZN => n1834);
   U1185 : AOI222_X1 port map( A1 => n1835, A2 => n1975, B1 => n1834, B2 => 
                           n2211, C1 => n1833, C2 => n1626, ZN => n1837);
   U1186 : OAI22_X1 port map( A1 => n2213, A2 => n1837, B1 => n1836, B2 => 
                           n2487, ZN => n1841);
   U1187 : OAI22_X1 port map( A1 => n1839, A2 => n2491, B1 => n1838, B2 => 
                           n2214, ZN => n1840);
   U1188 : AOI211_X1 port map( C1 => n1843, C2 => n1842, A => n1841, B => n1840
                           , ZN => n1844);
   U1189 : OAI22_X1 port map( A1 => n1845, A2 => n2497, B1 => n1844, B2 => 
                           n2499, ZN => n1851);
   U1190 : AOI22_X1 port map( A1 => n1848, A2 => n1847, B1 => n1846, B2 => 
                           n2384, ZN => n1849);
   U1191 : INV_X1 port map( A => n1849, ZN => n1850);
   U1192 : AOI211_X1 port map( C1 => n2373, C2 => n1852, A => n1851, B => n1850
                           , ZN => n1854);
   U1193 : OAI222_X1 port map( A1 => n2510, A2 => n1855, B1 => n2508, B2 => 
                           n1854, C1 => n1853, C2 => n2512, ZN => n1856);
   U1194 : AOI22_X1 port map( A1 => n2366, A2 => n1857, B1 => n2391, B2 => 
                           n1856, ZN => n1862);
   U1195 : OAI22_X1 port map( A1 => n2525_port, A2 => n1859, B1 => n1858, B2 =>
                           n1990, ZN => n1860);
   U1196 : INV_X1 port map( A => n1860, ZN => n1861);
   U1197 : OAI211_X1 port map( C1 => n1863, C2 => n2293, A => n1862, B => n1861
                           , ZN => n1865);
   U1198 : AOI22_X1 port map( A1 => n2526_port, A2 => n1865, B1 => n2228, B2 =>
                           n1864, ZN => n1870);
   U1199 : OAI22_X1 port map( A1 => n2537_port, A2 => n1867, B1 => n2147, B2 =>
                           n1866, ZN => n1868);
   U1200 : INV_X1 port map( A => n1868, ZN => n1869);
   U1201 : OAI211_X1 port map( C1 => n1871, C2 => n1994, A => n1870, B => n1869
                           , ZN => n1872);
   U1202 : AOI222_X1 port map( A1 => n1874, A2 => n2538_port, B1 => n1873, B2 
                           => n2543_port, C1 => n1872, C2 => n2541_port, ZN => 
                           n1875);
   U1203 : OAI22_X1 port map( A1 => n1876, A2 => n1921, B1 => n1875, B2 => 
                           n1948, ZN => n1877);
   U1204 : AOI211_X1 port map( C1 => n2235, C2 => n1920, A => n1878, B => n1877
                           , ZN => n1952);
   U1205 : NAND2_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, ZN => 
                           n1895);
   U1206 : OAI21_X1 port map( B1 => DATA1(23), B2 => DATA2_I_23_port, A => 
                           n1895, ZN => n2143);
   U1207 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n2144);
   U1208 : NAND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n1892);
   U1209 : INV_X1 port map( A => n1892, ZN => n2138);
   U1210 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n2134);
   U1211 : OAI21_X1 port map( B1 => DATA1(17), B2 => DATA2_I_17_port, A => 
                           n2134, ZN => n2298);
   U1212 : NAND2_X1 port map( A1 => n2284, A2 => DATA2_I_18_port, ZN => n2135);
   U1213 : OAI21_X1 port map( B1 => n2284, B2 => DATA2_I_18_port, A => n2135, 
                           ZN => n2272);
   U1214 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n2136);
   U1215 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => 
                           n2136, ZN => n2265);
   U1216 : NAND2_X1 port map( A1 => n2315, A2 => DATA2_I_16_port, ZN => n2299);
   U1217 : OAI21_X1 port map( B1 => n2315, B2 => DATA2_I_16_port, A => n2299, 
                           ZN => n2318);
   U1218 : NOR4_X1 port map( A1 => n2298, A2 => n2272, A3 => n2265, A4 => n2318
                           , ZN => n1891);
   U1219 : NAND2_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, ZN => 
                           n2329);
   U1220 : OAI21_X1 port map( B1 => DATA1(14), B2 => DATA2_I_14_port, A => 
                           n2329, ZN => n2363);
   U1221 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n1882);
   U1222 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => 
                           n1882, ZN => n2371);
   U1223 : NAND2_X1 port map( A1 => n2397, A2 => DATA2_I_12_port, ZN => n2370);
   U1224 : OAI21_X1 port map( B1 => n2397, B2 => DATA2_I_12_port, A => n2370, 
                           ZN => n1883);
   U1225 : NAND2_X1 port map( A1 => n2678, A2 => DATA2_I_11_port, ZN => n2327);
   U1226 : OAI21_X1 port map( B1 => n2678, B2 => DATA2_I_11_port, A => n2327, 
                           ZN => n2418);
   U1227 : NOR4_X1 port map( A1 => n2363, A2 => n2371, A3 => n1883, A4 => n2418
                           , ZN => n1887);
   U1228 : NAND2_X1 port map( A1 => n2576, A2 => DATA2_I_10_port, ZN => n2326);
   U1229 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => 
                           n2326, ZN => n2450);
   U1230 : NOR4_X1 port map( A1 => n1881, A2 => n1880, A3 => n2450, A4 => n1879
                           , ZN => n1886);
   U1231 : INV_X1 port map( A => n1882, ZN => n2351);
   U1232 : INV_X1 port map( A => n1883, ZN => n2405);
   U1233 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n1885);
   U1234 : INV_X1 port map( A => n1884, ZN => n2445);
   U1235 : AOI21_X1 port map( B1 => n2436, B2 => n2445, A => n2450, ZN => n2434
                           );
   U1236 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => n2576, A => n2434, 
                           ZN => n2419);
   U1237 : OAI21_X1 port map( B1 => n1885, B2 => n2419, A => n2327, ZN => n2404
                           );
   U1238 : NAND2_X1 port map( A1 => n2405, A2 => n2404, ZN => n2402);
   U1239 : AOI21_X1 port map( B1 => n2370, B2 => n2402, A => n2371, ZN => n2346
                           );
   U1240 : NOR2_X1 port map( A1 => n2351, A2 => n2346, ZN => n2345);
   U1241 : OAI21_X1 port map( B1 => n2345, B2 => n2363, A => n2329, ZN => n2338
                           );
   U1242 : AOI21_X1 port map( B1 => n1887, B2 => n1886, A => n2338, ZN => n1889
                           );
   U1243 : NAND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n1888);
   U1244 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => 
                           n1888, ZN => n2337);
   U1245 : OAI21_X1 port map( B1 => n1889, B2 => n2337, A => n1888, ZN => n2133
                           );
   U1246 : NOR2_X1 port map( A1 => n2299, A2 => n2298, ZN => n2297);
   U1247 : AOI21_X1 port map( B1 => DATA2_I_17_port, B2 => DATA1(17), A => 
                           n2297, ZN => n2273);
   U1248 : NOR2_X1 port map( A1 => n2273, A2 => n2272, ZN => n2271);
   U1249 : AOI21_X1 port map( B1 => DATA2_I_18_port, B2 => DATA1(18), A => 
                           n2271, ZN => n2253);
   U1250 : NOR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n1890);
   U1251 : OAI21_X1 port map( B1 => n2253, B2 => n1890, A => n2136, ZN => n2187
                           );
   U1252 : AOI21_X1 port map( B1 => n1891, B2 => n2133, A => n2187, ZN => n1893
                           );
   U1253 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n2137);
   U1254 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => 
                           n2137, ZN => n2199);
   U1255 : OAI21_X1 port map( B1 => DATA1(21), B2 => DATA2_I_21_port, A => 
                           n1892, ZN => n2184);
   U1256 : AOI221_X1 port map( B1 => n1893, B2 => n2137, C1 => n2199, C2 => 
                           n2137, A => n2184, ZN => n1894);
   U1257 : XOR2_X1 port map( A => n2161, B => DATA2_I_22_port, Z => n2170);
   U1258 : INV_X1 port map( A => n2170, ZN => n2172);
   U1259 : OAI21_X1 port map( B1 => n2138, B2 => n1894, A => n2172, ZN => n1896
                           );
   U1260 : OAI221_X1 port map( B1 => n2143, B2 => n2144, C1 => n2143, C2 => 
                           n1896, A => n1895, ZN => n1901);
   U1261 : NAND2_X1 port map( A1 => n2744, A2 => n1901, ZN => n2103);
   U1262 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n1906);
   U1263 : NAND2_X1 port map( A1 => DATA1(29), A2 => DATA2_I_29_port, ZN => 
                           n1899);
   U1264 : INV_X1 port map( A => n1899, ZN => n1963);
   U1265 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n2020);
   U1266 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n1898);
   U1267 : INV_X1 port map( A => n1898, ZN => n2053);
   U1268 : NAND2_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, ZN => 
                           n2068);
   U1269 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n1897);
   U1270 : INV_X1 port map( A => n1897, ZN => n2093);
   U1271 : NOR2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n2124);
   U1272 : OAI21_X1 port map( B1 => DATA1(25), B2 => DATA2_I_25_port, A => 
                           n1897, ZN => n2105);
   U1273 : NOR2_X1 port map( A1 => n2124, A2 => n2105, ZN => n2104);
   U1274 : XOR2_X1 port map( A => DATA1(26), B => DATA2_I_26_port, Z => n2092);
   U1275 : OAI21_X1 port map( B1 => n2093, B2 => n2104, A => n2092, ZN => n2057
                           );
   U1276 : OAI21_X1 port map( B1 => DATA1(27), B2 => DATA2_I_27_port, A => 
                           n1898, ZN => n2069);
   U1277 : AOI21_X1 port map( B1 => n2068, B2 => n2057, A => n2069, ZN => n2058
                           );
   U1278 : XNOR2_X1 port map( A => n2723, B => DATA2_I_28_port, ZN => n2052);
   U1279 : OAI21_X1 port map( B1 => n2053, B2 => n2058, A => n2052, ZN => n2037
                           );
   U1280 : OAI21_X1 port map( B1 => DATA1(29), B2 => DATA2_I_29_port, A => 
                           n1899, ZN => n2019);
   U1281 : AOI21_X1 port map( B1 => n2020, B2 => n2037, A => n2019, ZN => n1955
                           );
   U1282 : XOR2_X1 port map( A => DATA1(30), B => DATA2_I_30_port, Z => n1964);
   U1283 : OAI21_X1 port map( B1 => n1963, B2 => n1955, A => n1964, ZN => n1904
                           );
   U1284 : INV_X1 port map( A => n2105, ZN => n1900);
   U1285 : NAND3_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, A3 => 
                           n1900, ZN => n2096);
   U1286 : INV_X1 port map( A => n2096, ZN => n2102);
   U1287 : OAI21_X1 port map( B1 => n2093, B2 => n2102, A => n2092, ZN => n2065
                           );
   U1288 : AOI21_X1 port map( B1 => n2068, B2 => n2065, A => n2069, ZN => n2066
                           );
   U1289 : OAI21_X1 port map( B1 => n2053, B2 => n2066, A => n2052, ZN => n2016
                           );
   U1290 : AOI21_X1 port map( B1 => n2020, B2 => n2016, A => n2019, ZN => n1953
                           );
   U1291 : OAI21_X1 port map( B1 => n1963, B2 => n1953, A => n1964, ZN => n1905
                           );
   U1292 : NOR2_X1 port map( A1 => n3099, A2 => n1901, ZN => n2117);
   U1293 : INV_X1 port map( A => n2117, ZN => n2101);
   U1294 : AOI21_X1 port map( B1 => n1906, B2 => n1905, A => n2101, ZN => n1902
                           );
   U1295 : INV_X1 port map( A => n1902, ZN => n1903);
   U1296 : OAI221_X1 port map( B1 => n2103, B2 => n1906, C1 => n2103, C2 => 
                           n1904, A => n1903, ZN => n1915);
   U1297 : INV_X1 port map( A => DATA1(31), ZN => n2646);
   U1298 : XOR2_X1 port map( A => n2646, B => DATA2_I_31_port, Z => n1914);
   U1299 : INV_X1 port map( A => n2103, ZN => n2123);
   U1300 : NAND2_X1 port map( A1 => n2123, A2 => n1904, ZN => n1958);
   U1301 : NAND2_X1 port map( A1 => n2117, A2 => n1905, ZN => n1967);
   U1302 : NAND2_X1 port map( A1 => n1958, A2 => n1967, ZN => n1962);
   U1303 : NAND2_X1 port map( A1 => n1906, A2 => n1962, ZN => n1912);
   U1304 : OAI221_X1 port map( B1 => DATA1(31), B2 => n2462, C1 => n2646, C2 =>
                           n2458, A => n2437, ZN => n1907);
   U1305 : NOR2_X1 port map( A1 => DATA2(31), A2 => n2646, ZN => n2727);
   U1306 : AOI22_X1 port map( A1 => DATA2(31), A2 => n1907, B1 => n2727, B2 => 
                           n2438, ZN => n1908);
   U1307 : OAI21_X1 port map( B1 => n1909, B2 => n2455, A => n1908, ZN => n1910
                           );
   U1308 : AOI21_X1 port map( B1 => n2449, B2 => dataout_mul_31_port, A => 
                           n1910, ZN => n1911);
   U1309 : OAI21_X1 port map( B1 => n1912, B2 => n1914, A => n1911, ZN => n1913
                           );
   U1310 : AOI21_X1 port map( B1 => n1915, B2 => n1914, A => n1913, ZN => n1951
                           );
   U1311 : OR3_X1 port map( A1 => n2778, A2 => n1917, A3 => n1916, ZN => n1918)
                           ;
   U1312 : NOR2_X1 port map( A1 => n1919, A2 => n1918, ZN => n2738);
   U1313 : INV_X1 port map( A => n1920, ZN => n1949);
   U1314 : INV_X1 port map( A => n1921, ZN => n2550);
   U1315 : AOI22_X1 port map( A1 => n2550, A2 => n2063, B1 => n2235, B2 => 
                           n2014, ZN => n1947);
   U1316 : INV_X1 port map( A => n1922, ZN => n1941);
   U1317 : AOI22_X1 port map( A1 => n1925, A2 => n1924, B1 => n2156, B2 => 
                           n1923, ZN => n1929);
   U1318 : AOI22_X1 port map( A1 => n2160, A2 => n1927, B1 => n2219, B2 => 
                           n1926, ZN => n1928);
   U1319 : OAI211_X1 port map( C1 => n1930, C2 => n2214, A => n1929, B => n1928
                           , ZN => n2440);
   U1320 : AOI22_X1 port map( A1 => n2383, A2 => n2386, B1 => n1931, B2 => 
                           n2440, ZN => n1934);
   U1321 : AOI22_X1 port map( A1 => n2506, A2 => n2372, B1 => n1932, B2 => 
                           n2409, ZN => n1933);
   U1322 : OAI211_X1 port map( C1 => n1935, C2 => n2499, A => n1934, B => n1933
                           , ZN => n2356);
   U1323 : AOI222_X1 port map( A1 => n2356, A2 => n1938, B1 => n2322, B2 => 
                           n2321, C1 => n1937, C2 => n1936, ZN => n2307);
   U1324 : OAI22_X1 port map( A1 => n1990, A2 => n2307, B1 => n2269, B2 => 
                           n2268, ZN => n1940);
   U1325 : OAI22_X1 port map( A1 => n2254, A2 => n2293, B1 => n2294, B2 => 
                           n2525_port, ZN => n1939);
   U1326 : AOI211_X1 port map( C1 => n2517_port, C2 => n1941, A => n1940, B => 
                           n1939, ZN => n2191);
   U1327 : OAI22_X1 port map( A1 => n2154, A2 => n2153, B1 => n2191, B2 => 
                           n1994, ZN => n1943);
   U1328 : OAI22_X1 port map( A1 => n2146, A2 => n2537_port, B1 => n2176, B2 =>
                           n2147, ZN => n1942);
   U1329 : AOI211_X1 port map( C1 => n2526_port, C2 => n1944, A => n1943, B => 
                           n1942, ZN => n2114);
   U1330 : OAI222_X1 port map( A1 => n2100, A2 => n2099, B1 => n1999, B2 => 
                           n1945, C1 => n2114, C2 => n1996, ZN => n2080);
   U1331 : AOI22_X1 port map( A1 => n2552, A2 => n2080, B1 => n2546_port, B2 =>
                           n2036, ZN => n1946);
   U1332 : OAI211_X1 port map( C1 => n1949, C2 => n1948, A => n1947, B => n1946
                           , ZN => n1961);
   U1333 : NAND3_X1 port map( A1 => n2738, A2 => n2743, A3 => n1961, ZN => 
                           n1950);
   U1334 : OAI211_X1 port map( C1 => n1952, C2 => n2427, A => n1951, B => n1950
                           , ZN => OUTALU(31));
   U1335 : INV_X1 port map( A => n1953, ZN => n2015);
   U1336 : INV_X1 port map( A => DATA2(30), ZN => n2746);
   U1337 : AOI22_X1 port map( A1 => DATA1(30), A2 => n2746, B1 => DATA2(30), B2
                           => n2581, ZN => n2726);
   U1338 : AOI21_X1 port map( B1 => DATA1(30), B2 => n2412, A => n2410, ZN => 
                           n1954);
   U1339 : OAI22_X1 port map( A1 => n2726, A2 => n2462, B1 => n1954, B2 => 
                           n2746, ZN => n1960);
   U1340 : INV_X1 port map( A => n1955, ZN => n2017);
   U1341 : OAI22_X1 port map( A1 => n1968, A2 => n2646, B1 => n2474, B2 => 
                           n2581, ZN => n1956);
   U1342 : AOI22_X1 port map( A1 => n2736, A2 => n1956, B1 => n2468, B2 => 
                           dataout_mul_30_port, ZN => n1957);
   U1343 : OAI21_X1 port map( B1 => n2017, B2 => n1958, A => n1957, ZN => n1959
                           );
   U1344 : AOI211_X1 port map( C1 => n2441, C2 => n1961, A => n1960, B => n1959
                           , ZN => n1966);
   U1345 : OAI21_X1 port map( B1 => n1964, B2 => n1963, A => n1962, ZN => n1965
                           );
   U1346 : OAI211_X1 port map( C1 => n1967, C2 => n2015, A => n1966, B => n1965
                           , ZN => OUTALU(30));
   U1347 : NOR2_X1 port map( A1 => n2474, A2 => n2658, ZN => n1972);
   U1348 : NOR2_X1 port map( A1 => n1968, A2 => n2651, ZN => n2476);
   U1349 : AOI211_X1 port map( C1 => DATA1(0), C2 => n2040, A => n1972, B => 
                           n2476, ZN => n2013);
   U1350 : OAI22_X1 port map( A1 => n2003, A2 => n2461, B1 => n2005, B2 => 
                           n1969, ZN => n1970);
   U1351 : AOI22_X1 port map( A1 => dataout_mul_2_port, A2 => n2468, B1 => 
                           n2006, B2 => n1970, ZN => n2012);
   U1352 : OAI21_X1 port map( B1 => n2658, B2 => n2458, A => n2437, ZN => n2010
                           );
   U1353 : AOI22_X1 port map( A1 => n2546_port, A2 => n2551, B1 => n2235, B2 =>
                           n2549, ZN => n2002);
   U1354 : AOI22_X1 port map( A1 => n2431, A2 => n2531_port, B1 => n2530_port, 
                           B2 => n2229, ZN => n1993);
   U1355 : INV_X1 port map( A => n2502, ZN => n1985);
   U1356 : INV_X1 port map( A => n2215, ZN => n1981);
   U1357 : AOI211_X1 port map( C1 => DATA1(6), C2 => n2477, A => n1972, B => 
                           n1971, ZN => n1974);
   U1358 : OAI211_X1 port map( C1 => n2025, C2 => n2660, A => n1974, B => n1973
                           , ZN => n2479);
   U1359 : AOI222_X1 port map( A1 => n1976, A2 => n1975, B1 => n2479, B2 => 
                           n2483, C1 => n2212, C2 => n1626, ZN => n2486);
   U1360 : OAI22_X1 port map( A1 => n2213, A2 => n2486, B1 => n2488, B2 => 
                           n2487, ZN => n1980);
   U1361 : OAI22_X1 port map( A1 => n2489, A2 => n1978, B1 => n2490, B2 => 
                           n1977, ZN => n1979);
   U1362 : AOI211_X1 port map( C1 => n2219, C2 => n1981, A => n1980, B => n1979
                           , ZN => n2496);
   U1363 : OAI22_X1 port map( A1 => n2500, A2 => n2497, B1 => n2496, B2 => 
                           n2499, ZN => n1984);
   U1364 : OAI22_X1 port map( A1 => n2501, A2 => n1982, B1 => n2220, B2 => 
                           n2503, ZN => n1983);
   U1365 : AOI211_X1 port map( C1 => n2384, C2 => n1985, A => n1984, B => n1983
                           , ZN => n2513);
   U1366 : OAI222_X1 port map( A1 => n2510, A2 => n2224, B1 => n2508, B2 => 
                           n2513, C1 => n1986, C2 => n2512, ZN => n2515);
   U1367 : AOI22_X1 port map( A1 => n2388, A2 => n2225, B1 => n2391, B2 => 
                           n2515, ZN => n1988);
   U1368 : AOI22_X1 port map( A1 => n2518_port, A2 => n2206, B1 => n2366, B2 =>
                           n2520_port, ZN => n1987);
   U1369 : OAI211_X1 port map( C1 => n1990, C2 => n1989, A => n1988, B => n1987
                           , ZN => n2529_port);
   U1370 : INV_X1 port map( A => n1991, ZN => n2533_port);
   U1371 : AOI22_X1 port map( A1 => n2526_port, A2 => n2529_port, B1 => n2228, 
                           B2 => n2533_port, ZN => n1992);
   U1372 : OAI211_X1 port map( C1 => n1995, C2 => n1994, A => n1993, B => n1992
                           , ZN => n2539_port);
   U1373 : INV_X1 port map( A => n2539_port, ZN => n1998);
   U1374 : OAI222_X1 port map( A1 => n2100, A2 => n2000, B1 => n1999, B2 => 
                           n1998, C1 => n1997, C2 => n1996, ZN => n2545_port);
   U1375 : AOI22_X1 port map( A1 => n2548_port, A2 => n2545_port, B1 => n2550, 
                           B2 => n2236, ZN => n2001);
   U1376 : AOI21_X1 port map( B1 => n2002, B2 => n2001, A => n2455, ZN => n2009
                           );
   U1377 : AOI22_X1 port map( A1 => DATA2(2), A2 => n2658, B1 => DATA1(2), B2 
                           => n2776, ZN => n2653);
   U1378 : AOI22_X1 port map( A1 => n2466, A2 => n2005, B1 => n2004, B2 => 
                           n2003, ZN => n2007);
   U1379 : OAI22_X1 port map( A1 => n2653, A2 => n2462, B1 => n2007, B2 => 
                           n2006, ZN => n2008);
   U1380 : AOI211_X1 port map( C1 => DATA2(2), C2 => n2010, A => n2009, B => 
                           n2008, ZN => n2011);
   U1381 : OAI211_X1 port map( C1 => n2013, C2 => n2427, A => n2012, B => n2011
                           , ZN => OUTALU(2));
   U1382 : AOI22_X1 port map( A1 => n2548_port, A2 => n2014, B1 => n2546_port, 
                           B2 => n2063, ZN => n2035);
   U1383 : AOI22_X1 port map( A1 => n2235, A2 => n2036, B1 => n2550, B2 => 
                           n2080, ZN => n2034);
   U1384 : NAND2_X1 port map( A1 => n2015, A2 => n2117, ZN => n2018);
   U1385 : INV_X1 port map( A => n2018, ZN => n2032);
   U1386 : INV_X1 port map( A => n2016, ZN => n2049);
   U1387 : NAND2_X1 port map( A1 => n2123, A2 => n2017, ZN => n2029);
   U1388 : AOI22_X1 port map( A1 => n2020, A2 => n2019, B1 => n2018, B2 => 
                           n2029, ZN => n2031);
   U1389 : INV_X1 port map( A => DATA1(29), ZN => n2021);
   U1390 : NAND2_X1 port map( A1 => DATA2(29), A2 => n2021, ZN => n2725);
   U1391 : INV_X1 port map( A => DATA2(29), ZN => n2747);
   U1392 : NAND2_X1 port map( A1 => DATA1(29), A2 => n2747, ZN => n2722);
   U1393 : NAND2_X1 port map( A1 => n2725, A2 => n2722, ZN => n2567);
   U1394 : OAI21_X1 port map( B1 => n2021, B2 => n2458, A => n2437, ZN => n2022
                           );
   U1395 : AOI22_X1 port map( A1 => n2438, A2 => n2567, B1 => DATA2(29), B2 => 
                           n2022, ZN => n2028);
   U1396 : OAI211_X1 port map( C1 => n2025, C2 => n2646, A => n2024, B => n2023
                           , ZN => n2026);
   U1397 : AOI22_X1 port map( A1 => n2736, A2 => n2026, B1 => n2354, B2 => 
                           dataout_mul_29_port, ZN => n2027);
   U1398 : OAI211_X1 port map( C1 => n2037, C2 => n2029, A => n2028, B => n2027
                           , ZN => n2030);
   U1399 : AOI211_X1 port map( C1 => n2032, C2 => n2049, A => n2031, B => n2030
                           , ZN => n2033);
   U1400 : OAI221_X1 port map( B1 => n2427, B2 => n2035, C1 => n2427, C2 => 
                           n2034, A => n2033, ZN => OUTALU(29));
   U1401 : AOI222_X1 port map( A1 => n2036, A2 => n2548_port, B1 => n2080, B2 
                           => n2546_port, C1 => n2063, C2 => n2235, ZN => n2056
                           );
   U1402 : AND2_X1 port map( A1 => n2037, A2 => n2123, ZN => n2050);
   U1403 : INV_X1 port map( A => n2066, ZN => n2038);
   U1404 : NOR3_X1 port map( A1 => n2052, A2 => n2038, A3 => n2101, ZN => n2048
                           );
   U1405 : INV_X1 port map( A => DATA2(28), ZN => n2748);
   U1406 : AOI22_X1 port map( A1 => DATA1(28), A2 => n2748, B1 => DATA2(28), B2
                           => n2723, ZN => n2718);
   U1407 : AOI22_X1 port map( A1 => n2040, A2 => DATA1(30), B1 => n2039, B2 => 
                           DATA1(31), ZN => n2043);
   U1408 : NAND3_X1 port map( A1 => n2043, A2 => n2042, A3 => n2041, ZN => 
                           n2044);
   U1409 : AOI22_X1 port map( A1 => n2736, A2 => n2044, B1 => n2449, B2 => 
                           dataout_mul_28_port, ZN => n2046);
   U1410 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => DATA2(28), B => 
                           DATA1(28), ZN => n2045);
   U1411 : OAI211_X1 port map( C1 => n2718, C2 => n2462, A => n2046, B => n2045
                           , ZN => n2047);
   U1412 : AOI211_X1 port map( C1 => n2050, C2 => n2058, A => n2048, B => n2047
                           , ZN => n2055);
   U1413 : NOR2_X1 port map( A1 => n2049, A2 => n2101, ZN => n2051);
   U1414 : OAI22_X1 port map( A1 => n2053, A2 => n2052, B1 => n2051, B2 => 
                           n2050, ZN => n2054);
   U1415 : OAI211_X1 port map( C1 => n2056, C2 => n2427, A => n2055, B => n2054
                           , ZN => OUTALU(28));
   U1416 : INV_X1 port map( A => n2057, ZN => n2079);
   U1417 : NOR2_X1 port map( A1 => n2058, A2 => n2103, ZN => n2070);
   U1418 : AOI22_X1 port map( A1 => n2079, A2 => n2070, B1 => n2468, B2 => 
                           dataout_mul_27_port, ZN => n2077);
   U1419 : INV_X1 port map( A => DATA2(27), ZN => n2749);
   U1420 : OAI21_X1 port map( B1 => n2458, B2 => n2749, A => n2437, ZN => n2062
                           );
   U1421 : NOR3_X1 port map( A1 => n2082, A2 => n2455, A3 => n2083, ZN => n2061
                           );
   U1422 : NAND2_X1 port map( A1 => n2059, A2 => DATA2(27), ZN => n2717);
   U1423 : NAND2_X1 port map( A1 => DATA1(27), A2 => n2749, ZN => n2641);
   U1424 : AOI21_X1 port map( B1 => n2717, B2 => n2641, A => n2462, ZN => n2060
                           );
   U1425 : AOI211_X1 port map( C1 => DATA1(27), C2 => n2062, A => n2061, B => 
                           n2060, ZN => n2076);
   U1426 : AOI22_X1 port map( A1 => n2080, A2 => n2235, B1 => n2063, B2 => 
                           n2548_port, ZN => n2064);
   U1427 : INV_X1 port map( A => n2064, ZN => n2067);
   U1428 : INV_X1 port map( A => n2065, ZN => n2078);
   U1429 : NOR2_X1 port map( A1 => n2066, A2 => n2101, ZN => n2071);
   U1430 : AOI22_X1 port map( A1 => n2441, A2 => n2067, B1 => n2078, B2 => 
                           n2071, ZN => n2075);
   U1431 : INV_X1 port map( A => n2068, ZN => n2073);
   U1432 : INV_X1 port map( A => n2069, ZN => n2072);
   U1433 : OAI22_X1 port map( A1 => n2073, A2 => n2072, B1 => n2071, B2 => 
                           n2070, ZN => n2074);
   U1434 : NAND4_X1 port map( A1 => n2077, A2 => n2076, A3 => n2075, A4 => 
                           n2074, ZN => OUTALU(27));
   U1435 : NOR2_X1 port map( A1 => n2101, A2 => n2078, ZN => n2091);
   U1436 : INV_X1 port map( A => n2091, ZN => n2097);
   U1437 : NOR2_X1 port map( A1 => n2079, A2 => n2103, ZN => n2090);
   U1438 : AND3_X1 port map( A1 => n2080, A2 => n2548_port, A3 => n2441, ZN => 
                           n2089);
   U1439 : INV_X1 port map( A => DATA2(26), ZN => n2750);
   U1440 : OAI22_X1 port map( A1 => n2557, A2 => n2750, B1 => DATA2(26), B2 => 
                           DATA1(26), ZN => n2638);
   U1441 : OAI22_X1 port map( A1 => n2084, A2 => n2083, B1 => n2082, B2 => 
                           n2081, ZN => n2085);
   U1442 : AOI22_X1 port map( A1 => n2736, A2 => n2085, B1 => n2354, B2 => 
                           dataout_mul_26_port, ZN => n2087);
   U1443 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => DATA2(26), B => 
                           DATA1(26), ZN => n2086);
   U1444 : OAI211_X1 port map( C1 => n2638, C2 => n2462, A => n2087, B => n2086
                           , ZN => n2088);
   U1445 : AOI211_X1 port map( C1 => n2090, C2 => n2104, A => n2089, B => n2088
                           , ZN => n2095);
   U1446 : OAI22_X1 port map( A1 => n2093, A2 => n2092, B1 => n2091, B2 => 
                           n2090, ZN => n2094);
   U1447 : OAI211_X1 port map( C1 => n2097, C2 => n2096, A => n2095, B => n2094
                           , ZN => OUTALU(26));
   U1448 : NAND2_X1 port map( A1 => DATA2(25), A2 => n2716, ZN => n2098);
   U1449 : OAI21_X1 port map( B1 => DATA2(25), B2 => n2716, A => n2098, ZN => 
                           n2566);
   U1450 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_25_port, B1 => 
                           n2438, B2 => n2566, ZN => n2112);
   U1451 : OAI22_X1 port map( A1 => n2114, A2 => n2100, B1 => n2099, B2 => 
                           n2113, ZN => n2108);
   U1452 : NAND2_X1 port map( A1 => DATA1(24), A2 => DATA2_I_24_port, ZN => 
                           n2116);
   U1453 : AOI211_X1 port map( C1 => n2116, C2 => n2105, A => n2102, B => n2101
                           , ZN => n2107);
   U1454 : AOI211_X1 port map( C1 => n2124, C2 => n2105, A => n2104, B => n2103
                           , ZN => n2106);
   U1455 : AOI211_X1 port map( C1 => n2441, C2 => n2108, A => n2107, B => n2106
                           , ZN => n2111);
   U1456 : NAND3_X1 port map( A1 => n2736, A2 => n2156, A3 => n2158, ZN => 
                           n2110);
   U1457 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => DATA2(25), B => 
                           DATA1(25), ZN => n2109);
   U1458 : NAND4_X1 port map( A1 => n2112, A2 => n2111, A3 => n2110, A4 => 
                           n2109, ZN => OUTALU(25));
   U1459 : AOI22_X1 port map( A1 => DATA2_I_24_port, A2 => n2123, B1 => n2412, 
                           B2 => DATA2(24), ZN => n2126);
   U1460 : NOR3_X1 port map( A1 => n2114, A2 => n2113, A3 => n2427, ZN => n2122
                           );
   U1461 : AOI22_X1 port map( A1 => n2494, A2 => n2158, B1 => n2156, B2 => 
                           n2159, ZN => n2120);
   U1462 : INV_X1 port map( A => DATA2(24), ZN => n2752);
   U1463 : OAI22_X1 port map( A1 => n2709, A2 => DATA2(24), B1 => n2752, B2 => 
                           DATA1(24), ZN => n2706);
   U1464 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_24_port, B1 => 
                           n2438, B2 => n2706, ZN => n2119);
   U1465 : INV_X1 port map( A => n2124, ZN => n2115);
   U1466 : NAND3_X1 port map( A1 => n2117, A2 => n2116, A3 => n2115, ZN => 
                           n2118);
   U1467 : OAI211_X1 port map( C1 => n2120, C2 => n2455, A => n2119, B => n2118
                           , ZN => n2121);
   U1468 : AOI211_X1 port map( C1 => n2124, C2 => n2123, A => n2122, B => n2121
                           , ZN => n2125);
   U1469 : OAI221_X1 port map( B1 => n2709, B2 => n2126, C1 => n2709, C2 => 
                           n2437, A => n2125, ZN => OUTALU(24));
   U1470 : NAND2_X1 port map( A1 => DATA2(23), A2 => n2128, ZN => n2712);
   U1471 : INV_X1 port map( A => DATA2(23), ZN => n2753);
   U1472 : NAND2_X1 port map( A1 => DATA1(23), A2 => n2753, ZN => n2634);
   U1473 : AOI21_X1 port map( B1 => n2712, B2 => n2634, A => n2462, ZN => n2132
                           );
   U1474 : AOI222_X1 port map( A1 => n2157, A2 => n2156, B1 => n2159, B2 => 
                           n2494, C1 => n2158, C2 => n2127, ZN => n2130);
   U1475 : AOI21_X1 port map( B1 => n2412, B2 => DATA2(23), A => n2410, ZN => 
                           n2129);
   U1476 : OAI22_X1 port map( A1 => n2130, A2 => n2455, B1 => n2129, B2 => 
                           n2128, ZN => n2131);
   U1477 : AOI211_X1 port map( C1 => n2449, C2 => dataout_mul_23_port, A => 
                           n2132, B => n2131, ZN => n2152);
   U1478 : NOR2_X1 port map( A1 => n3099, A2 => n2133, ZN => n2252);
   U1479 : INV_X1 port map( A => n2184, ZN => n2186);
   U1480 : INV_X1 port map( A => n2187, ZN => n2190);
   U1481 : OAI21_X1 port map( B1 => n2190, B2 => n2199, A => n2137, ZN => n2174
                           );
   U1482 : AOI21_X1 port map( B1 => n2186, B2 => n2174, A => n2138, ZN => n2140
                           );
   U1483 : NAND2_X1 port map( A1 => n2133, A2 => n2744, ZN => n2319);
   U1484 : INV_X1 port map( A => n2319, ZN => n2286);
   U1485 : INV_X1 port map( A => n2272, ZN => n2288);
   U1486 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n2296);
   U1487 : OAI21_X1 port map( B1 => n2296, B2 => n2298, A => n2134, ZN => n2287
                           );
   U1488 : NAND2_X1 port map( A1 => n2288, A2 => n2287, ZN => n2285);
   U1489 : AND2_X1 port map( A1 => n2135, A2 => n2285, ZN => n2251);
   U1490 : OAI21_X1 port map( B1 => n2265, B2 => n2251, A => n2136, ZN => n2188
                           );
   U1491 : INV_X1 port map( A => n2188, ZN => n2189);
   U1492 : OAI21_X1 port map( B1 => n2189, B2 => n2199, A => n2137, ZN => n2173
                           );
   U1493 : AOI21_X1 port map( B1 => n2186, B2 => n2173, A => n2138, ZN => n2139
                           );
   U1494 : AOI22_X1 port map( A1 => n2252, A2 => n2140, B1 => n2286, B2 => 
                           n2139, ZN => n2169);
   U1495 : AOI211_X1 port map( C1 => n2169, C2 => n2172, A => n2143, B => n3099
                           , ZN => n2145);
   U1496 : INV_X1 port map( A => n2252, ZN => n2317);
   U1497 : OAI22_X1 port map( A1 => n2317, A2 => n2140, B1 => n2319, B2 => 
                           n2139, ZN => n2141);
   U1498 : INV_X1 port map( A => n2141, ZN => n2171);
   U1499 : OAI22_X1 port map( A1 => n2171, A2 => n2170, B1 => n3099, B2 => 
                           n2144, ZN => n2142);
   U1500 : AOI22_X1 port map( A1 => n2145, A2 => n2144, B1 => n2143, B2 => 
                           n2142, ZN => n2151);
   U1501 : OAI22_X1 port map( A1 => n2146, A2 => n2420, B1 => n2154, B2 => 
                           n2537_port, ZN => n2149);
   U1502 : OAI22_X1 port map( A1 => n2176, A2 => n2153, B1 => n2191, B2 => 
                           n2147, ZN => n2148);
   U1503 : OAI21_X1 port map( B1 => n2149, B2 => n2148, A => n2441, ZN => n2150
                           );
   U1504 : NAND3_X1 port map( A1 => n2152, A2 => n2151, A3 => n2150, ZN => 
                           OUTALU(23));
   U1505 : OAI222_X1 port map( A1 => n2420, A2 => n2154, B1 => n2153, B2 => 
                           n2191, C1 => n2537_port, C2 => n2176, ZN => n2167);
   U1506 : INV_X1 port map( A => DATA2(22), ZN => n2754);
   U1507 : AOI211_X1 port map( C1 => n2437, C2 => n2458, A => n2161, B => n2754
                           , ZN => n2166);
   U1508 : AOI22_X1 port map( A1 => n2494, A2 => n2157, B1 => n2156, B2 => 
                           n2155, ZN => n2164);
   U1509 : AOI22_X1 port map( A1 => n2160, A2 => n2159, B1 => n2219, B2 => 
                           n2158, ZN => n2163);
   U1510 : OAI22_X1 port map( A1 => n2161, A2 => n2754, B1 => DATA2(22), B2 => 
                           DATA1(22), ZN => n2703);
   U1511 : INV_X1 port map( A => n2703, ZN => n2630);
   U1512 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_22_port, B1 => 
                           n2438, B2 => n2630, ZN => n2162);
   U1513 : OAI221_X1 port map( B1 => n2455, B2 => n2164, C1 => n2455, C2 => 
                           n2163, A => n2162, ZN => n2165);
   U1514 : AOI211_X1 port map( C1 => n2441, C2 => n2167, A => n2166, B => n2165
                           , ZN => n2168);
   U1515 : OAI221_X1 port map( B1 => n2172, B2 => n2171, C1 => n2170, C2 => 
                           n2169, A => n2168, ZN => OUTALU(22));
   U1516 : AOI22_X1 port map( A1 => n2252, A2 => n2174, B1 => n2286, B2 => 
                           n2173, ZN => n2185);
   U1517 : OAI22_X1 port map( A1 => n2317, A2 => n2174, B1 => n2319, B2 => 
                           n2173, ZN => n2175);
   U1518 : INV_X1 port map( A => n2175, ZN => n2183);
   U1519 : OAI22_X1 port map( A1 => n2176, A2 => n2420, B1 => n2191, B2 => 
                           n2537_port, ZN => n2181);
   U1520 : AOI21_X1 port map( B1 => n2412, B2 => DATA2(21), A => n2410, ZN => 
                           n2179);
   U1521 : NAND2_X1 port map( A1 => DATA2(21), A2 => n2700, ZN => n2702);
   U1522 : OAI21_X1 port map( B1 => DATA2(21), B2 => n2700, A => n2702, ZN => 
                           n2569);
   U1523 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_21_port, B1 => 
                           n2438, B2 => n2569, ZN => n2178);
   U1524 : NAND3_X1 port map( A1 => n2736, A2 => n2442, A3 => n2276, ZN => 
                           n2177);
   U1525 : OAI211_X1 port map( C1 => n2179, C2 => n2700, A => n2178, B => n2177
                           , ZN => n2180);
   U1526 : AOI21_X1 port map( B1 => n2441, B2 => n2181, A => n2180, ZN => n2182
                           );
   U1527 : OAI221_X1 port map( B1 => n2186, B2 => n2185, C1 => n2184, C2 => 
                           n2183, A => n2182, ZN => OUTALU(21));
   U1528 : INV_X1 port map( A => n2199, ZN => n2201);
   U1529 : AOI22_X1 port map( A1 => n2286, A2 => n2188, B1 => n2252, B2 => 
                           n2187, ZN => n2200);
   U1530 : AOI22_X1 port map( A1 => n2190, A2 => n2252, B1 => n2286, B2 => 
                           n2189, ZN => n2198);
   U1531 : INV_X1 port map( A => DATA2(20), ZN => n2756);
   U1532 : OAI21_X1 port map( B1 => n2458, B2 => n2756, A => n2437, ZN => n2196
                           );
   U1533 : NOR3_X1 port map( A1 => n2191, A2 => n2420, A3 => n2427, ZN => n2195
                           );
   U1534 : AOI22_X1 port map( A1 => n2385, A2 => n2274, B1 => n2384, B2 => 
                           n2276, ZN => n2193);
   U1535 : OAI22_X1 port map( A1 => n2701, A2 => DATA2(20), B1 => n2756, B2 => 
                           DATA1(20), ZN => n2696);
   U1536 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_20_port, B1 => 
                           n2438, B2 => n2696, ZN => n2192);
   U1537 : OAI21_X1 port map( B1 => n2193, B2 => n2455, A => n2192, ZN => n2194
                           );
   U1538 : AOI211_X1 port map( C1 => DATA1(20), C2 => n2196, A => n2195, B => 
                           n2194, ZN => n2197);
   U1539 : OAI221_X1 port map( B1 => n2201, B2 => n2200, C1 => n2199, C2 => 
                           n2198, A => n2197, ZN => OUTALU(20));
   U1540 : AOI22_X1 port map( A1 => DATA2(1), A2 => DATA1(1), B1 => n2651, B2 
                           => n2777, ZN => n2558);
   U1541 : AND2_X1 port map( A1 => n2438, A2 => n2558, ZN => n2204);
   U1542 : AOI211_X1 port map( C1 => n2459, C2 => n2243, A => n2202, B => n2461
                           , ZN => n2203);
   U1543 : AOI211_X1 port map( C1 => n2449, C2 => dataout_mul_1_port, A => 
                           n2204, B => n2203, ZN => n2249);
   U1544 : AOI21_X1 port map( B1 => n2441, B2 => n2205, A => n2410, ZN => n2457
                           );
   U1545 : OAI21_X1 port map( B1 => n2777, B2 => n2458, A => n2457, ZN => n2241
                           );
   U1546 : INV_X1 port map( A => n2529_port, ZN => n2232);
   U1547 : INV_X1 port map( A => n2206, ZN => n2524_port);
   U1548 : INV_X1 port map( A => n2496, ZN => n2223);
   U1549 : AOI211_X1 port map( C1 => DATA1(5), C2 => n2477, A => n2208, B => 
                           n2207, ZN => n2210);
   U1550 : OAI211_X1 port map( C1 => n2474, C2 => n2651, A => n2210, B => n2209
                           , ZN => n2481);
   U1551 : AOI222_X1 port map( A1 => n2212, A2 => n2480, B1 => n2481, B2 => 
                           n2211, C1 => n2479, C2 => n1626, ZN => n2471);
   U1552 : OAI22_X1 port map( A1 => n2213, A2 => n2471, B1 => n2490, B2 => 
                           n2487, ZN => n2217);
   U1553 : OAI22_X1 port map( A1 => n2489, A2 => n2215, B1 => n2486, B2 => 
                           n2214, ZN => n2216);
   U1554 : AOI211_X1 port map( C1 => n2219, C2 => n2218, A => n2217, B => n2216
                           , ZN => n2470);
   U1555 : OAI22_X1 port map( A1 => n2502, A2 => n2497, B1 => n2470, B2 => 
                           n2499, ZN => n2222);
   U1556 : OAI22_X1 port map( A1 => n2501, A2 => n2220, B1 => n2500, B2 => 
                           n2503, ZN => n2221);
   U1557 : AOI211_X1 port map( C1 => n2384, C2 => n2223, A => n2222, B => n2221
                           , ZN => n2511);
   U1558 : OAI222_X1 port map( A1 => n2510, A2 => n2513, B1 => n2508, B2 => 
                           n2511, C1 => n2224, C2 => n2512, ZN => n2519_port);
   U1559 : AOI22_X1 port map( A1 => n2388, A2 => n2520_port, B1 => n2391, B2 =>
                           n2519_port, ZN => n2227);
   U1560 : AOI22_X1 port map( A1 => n2518_port, A2 => n2515, B1 => n2521_port, 
                           B2 => n2225, ZN => n2226);
   U1561 : OAI211_X1 port map( C1 => n2524_port, C2 => n2268, A => n2227, B => 
                           n2226, ZN => n2469);
   U1562 : AOI22_X1 port map( A1 => n2526_port, A2 => n2469, B1 => n2228, B2 =>
                           n2531_port, ZN => n2231);
   U1563 : AOI22_X1 port map( A1 => n2532_port, A2 => n2229, B1 => n2530_port, 
                           B2 => n2533_port, ZN => n2230);
   U1564 : OAI211_X1 port map( C1 => n2232, C2 => n2537_port, A => n2231, B => 
                           n2230, ZN => n2542_port);
   U1565 : AOI222_X1 port map( A1 => n2233, A2 => n2538_port, B1 => n2539_port,
                           B2 => n2543_port, C1 => n2542_port, C2 => n2541_port
                           , ZN => n2556);
   U1566 : INV_X1 port map( A => n2556, ZN => n2234);
   U1567 : AOI22_X1 port map( A1 => n2548_port, A2 => n2234, B1 => n2550, B2 =>
                           n2551, ZN => n2238);
   U1568 : AOI22_X1 port map( A1 => n2552, A2 => n2236, B1 => n2235, B2 => 
                           n2545_port, ZN => n2237);
   U1569 : OAI211_X1 port map( C1 => n2240, C2 => n2239, A => n2238, B => n2237
                           , ZN => n2737);
   U1570 : AOI22_X1 port map( A1 => DATA1(1), A2 => n2241, B1 => n2736, B2 => 
                           n2737, ZN => n2248);
   U1571 : NAND3_X1 port map( A1 => n2242, A2 => DATA1(0), A3 => n2441, ZN => 
                           n2247);
   U1572 : OAI221_X1 port map( B1 => n2460, B2 => n2245, C1 => n2244, C2 => 
                           n2243, A => n2466, ZN => n2246);
   U1573 : NAND4_X1 port map( A1 => n2249, A2 => n2248, A3 => n2247, A4 => 
                           n2246, ZN => OUTALU(1));
   U1574 : INV_X1 port map( A => n2265, ZN => n2267);
   U1575 : OAI22_X1 port map( A1 => n2319, A2 => n2251, B1 => n2317, B2 => 
                           n2253, ZN => n2250);
   U1576 : INV_X1 port map( A => n2250, ZN => n2266);
   U1577 : AOI22_X1 port map( A1 => n2253, A2 => n2252, B1 => n2286, B2 => 
                           n2251, ZN => n2264);
   U1578 : OAI22_X1 port map( A1 => n2323, A2 => n2254, B1 => n2269, B2 => 
                           n2293, ZN => n2262);
   U1579 : OAI22_X1 port map( A1 => n2294, A2 => n2268, B1 => n2307, B2 => 
                           n2525_port, ZN => n2261);
   U1580 : AOI222_X1 port map( A1 => n2275, A2 => n2442, B1 => n2274, B2 => 
                           n2384, C1 => n2276, C2 => n2383, ZN => n2259);
   U1581 : INV_X1 port map( A => DATA2(19), ZN => n2757);
   U1582 : OAI21_X1 port map( B1 => n2458, B2 => n2757, A => n2437, ZN => n2255
                           );
   U1583 : AOI22_X1 port map( A1 => n2256, A2 => n2255, B1 => n2449, B2 => 
                           dataout_mul_19_port, ZN => n2258);
   U1584 : NOR2_X1 port map( A1 => DATA1(19), A2 => n2757, ZN => n2697);
   U1585 : NAND2_X1 port map( A1 => n2256, A2 => n2757, ZN => n2626);
   U1586 : INV_X1 port map( A => n2626, ZN => n2562);
   U1587 : OAI21_X1 port map( B1 => n2697, B2 => n2562, A => n2438, ZN => n2257
                           );
   U1588 : OAI211_X1 port map( C1 => n2259, C2 => n2455, A => n2258, B => n2257
                           , ZN => n2260);
   U1589 : AOI221_X1 port map( B1 => n2262, B2 => n2441, C1 => n2261, C2 => 
                           n2441, A => n2260, ZN => n2263);
   U1590 : OAI221_X1 port map( B1 => n2267, B2 => n2266, C1 => n2265, C2 => 
                           n2264, A => n2263, ZN => OUTALU(19));
   U1591 : OAI222_X1 port map( A1 => n2269, A2 => n2323, B1 => n2307, B2 => 
                           n2268, C1 => n2294, C2 => n2293, ZN => n2270);
   U1592 : INV_X1 port map( A => n2270, ZN => n2291);
   U1593 : INV_X1 port map( A => DATA2(18), ZN => n2758);
   U1594 : OAI21_X1 port map( B1 => n2458, B2 => n2758, A => n2437, ZN => n2283
                           );
   U1595 : AOI211_X1 port map( C1 => n2273, C2 => n2272, A => n2271, B => n2317
                           , ZN => n2282);
   U1596 : AOI22_X1 port map( A1 => n2506, A2 => n2275, B1 => n2383, B2 => 
                           n2274, ZN => n2280);
   U1597 : AOI22_X1 port map( A1 => n2385, A2 => n2277, B1 => n2373, B2 => 
                           n2276, ZN => n2279);
   U1598 : INV_X1 port map( A => DATA1(18), ZN => n2584);
   U1599 : OAI22_X1 port map( A1 => n2584, A2 => n2758, B1 => DATA2(18), B2 => 
                           n2284, ZN => n2693);
   U1600 : INV_X1 port map( A => n2693, ZN => n2623);
   U1601 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_18_port, B1 => 
                           n2438, B2 => n2623, ZN => n2278);
   U1602 : OAI221_X1 port map( B1 => n2455, B2 => n2280, C1 => n2455, C2 => 
                           n2279, A => n2278, ZN => n2281);
   U1603 : AOI211_X1 port map( C1 => n2284, C2 => n2283, A => n2282, B => n2281
                           , ZN => n2290);
   U1604 : OAI211_X1 port map( C1 => n2288, C2 => n2287, A => n2286, B => n2285
                           , ZN => n2289);
   U1605 : OAI211_X1 port map( C1 => n2291, C2 => n2427, A => n2290, B => n2289
                           , ZN => OUTALU(18));
   U1606 : NAND2_X1 port map( A1 => DATA2(17), A2 => n2292, ZN => n2692);
   U1607 : NOR2_X1 port map( A1 => n2292, A2 => DATA2(17), ZN => n2624);
   U1608 : INV_X1 port map( A => n2624, ZN => n2690);
   U1609 : NAND2_X1 port map( A1 => n2692, A2 => n2690, ZN => n2568);
   U1610 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_17_port, B1 => 
                           n2438, B2 => n2568, ZN => n2306);
   U1611 : OAI22_X1 port map( A1 => n2323, A2 => n2294, B1 => n2307, B2 => 
                           n2293, ZN => n2302);
   U1612 : NOR2_X1 port map( A1 => n2296, A2 => n2298, ZN => n2295);
   U1613 : AOI211_X1 port map( C1 => n2296, C2 => n2298, A => n2295, B => n2319
                           , ZN => n2301);
   U1614 : AOI211_X1 port map( C1 => n2299, C2 => n2298, A => n2297, B => n2317
                           , ZN => n2300);
   U1615 : AOI211_X1 port map( C1 => n2441, C2 => n2302, A => n2301, B => n2300
                           , ZN => n2305);
   U1616 : NAND3_X1 port map( A1 => n2736, A2 => n2357, A3 => n2308, ZN => 
                           n2304);
   U1617 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => DATA1(17), B => 
                           DATA2(17), ZN => n2303);
   U1618 : NAND4_X1 port map( A1 => n2306, A2 => n2305, A3 => n2304, A4 => 
                           n2303, ZN => OUTALU(17));
   U1619 : INV_X1 port map( A => n2318, ZN => n2320);
   U1620 : INV_X1 port map( A => DATA2(16), ZN => n2760);
   U1621 : OAI21_X1 port map( B1 => n2458, B2 => n2760, A => n2437, ZN => n2314
                           );
   U1622 : NOR3_X1 port map( A1 => n2323, A2 => n2307, A3 => n2427, ZN => n2313
                           );
   U1623 : AOI22_X1 port map( A1 => n2357, A2 => n2309, B1 => n2321, B2 => 
                           n2308, ZN => n2311);
   U1624 : OAI22_X1 port map( A1 => n2691, A2 => DATA2(16), B1 => n2760, B2 => 
                           n2315, ZN => n2686);
   U1625 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_16_port, B1 => 
                           n2438, B2 => n2686, ZN => n2310);
   U1626 : OAI21_X1 port map( B1 => n2311, B2 => n2455, A => n2310, ZN => n2312
                           );
   U1627 : AOI211_X1 port map( C1 => n2315, C2 => n2314, A => n2313, B => n2312
                           , ZN => n2316);
   U1628 : OAI221_X1 port map( B1 => n2320, B2 => n2319, C1 => n2318, C2 => 
                           n2317, A => n2316, ZN => OUTALU(16));
   U1629 : AOI22_X1 port map( A1 => n2357, A2 => n2322, B1 => n2321, B2 => 
                           n2356, ZN => n2342);
   U1630 : NOR3_X1 port map( A1 => n2323, A2 => n2343, A3 => n2455, ZN => n2335
                           );
   U1631 : INV_X1 port map( A => n2337, ZN => n2339);
   U1632 : INV_X1 port map( A => n2452, ZN => n2324);
   U1633 : AOI21_X1 port map( B1 => n2436, B2 => n2324, A => n2450, ZN => n2325
                           );
   U1634 : INV_X1 port map( A => n2325, ZN => n2432);
   U1635 : NAND2_X1 port map( A1 => n2326, A2 => n2432, ZN => n2415);
   U1636 : INV_X1 port map( A => n2415, ZN => n2328);
   U1637 : OAI21_X1 port map( B1 => n2418, B2 => n2328, A => n2327, ZN => n2396
                           );
   U1638 : NAND2_X1 port map( A1 => n2396, A2 => n2405, ZN => n2395);
   U1639 : AOI21_X1 port map( B1 => n2370, B2 => n2395, A => n2371, ZN => n2348
                           );
   U1640 : NOR2_X1 port map( A1 => n2351, A2 => n2348, ZN => n2344);
   U1641 : OAI21_X1 port map( B1 => n2344, B2 => n2363, A => n2329, ZN => n2330
                           );
   U1642 : XNOR2_X1 port map( A => n2339, B => n2330, ZN => n2333);
   U1643 : INV_X1 port map( A => DATA2(15), ZN => n2761);
   U1644 : NOR2_X1 port map( A1 => DATA1(15), A2 => n2761, ZN => n2687);
   U1645 : NOR2_X1 port map( A1 => DATA2(15), A2 => n2577, ZN => n2619);
   U1646 : OAI21_X1 port map( B1 => n2687, B2 => n2619, A => n2438, ZN => n2332
                           );
   U1647 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => DATA2(15), B => 
                           n3098, ZN => n2331);
   U1648 : OAI211_X1 port map( C1 => n2333, C2 => n2347, A => n2332, B => n2331
                           , ZN => n2334);
   U1649 : AOI211_X1 port map( C1 => n2449, C2 => dataout_mul_15_port, A => 
                           n2335, B => n2334, ZN => n2341);
   U1650 : INV_X1 port map( A => n2338, ZN => n2336);
   U1651 : INV_X1 port map( A => n2433, ZN => n2403);
   U1652 : OAI221_X1 port map( B1 => n2339, B2 => n2338, C1 => n2337, C2 => 
                           n2336, A => n2403, ZN => n2340);
   U1653 : OAI211_X1 port map( C1 => n2342, C2 => n2427, A => n2341, B => n2340
                           , ZN => OUTALU(15));
   U1654 : INV_X1 port map( A => n2343, ZN => n2387);
   U1655 : AOI22_X1 port map( A1 => n2518_port, A2 => n2387, B1 => n2391, B2 =>
                           n2389, ZN => n2365);
   U1656 : OAI22_X1 port map( A1 => n2345, A2 => n2433, B1 => n2344, B2 => 
                           n2347, ZN => n2362);
   U1657 : INV_X1 port map( A => n2346, ZN => n2350);
   U1658 : NOR2_X1 port map( A1 => n2348, A2 => n2347, ZN => n2349);
   U1659 : AOI21_X1 port map( B1 => n2403, B2 => n2350, A => n2349, ZN => n2369
                           );
   U1660 : NOR3_X1 port map( A1 => n2351, A2 => n2369, A3 => n2363, ZN => n2361
                           );
   U1661 : INV_X1 port map( A => DATA2(14), ZN => n2762);
   U1662 : AOI22_X1 port map( A1 => DATA1(14), A2 => n2762, B1 => DATA2(14), B2
                           => n2578, ZN => n2683);
   U1663 : OAI21_X1 port map( B1 => n2578, B2 => n2458, A => n2437, ZN => n2355
                           );
   U1664 : XOR2_X1 port map( A => boothmul_pipelined_i_sum_B_in_7_14_port, B =>
                           n2352, Z => n2353);
   U1665 : AOI22_X1 port map( A1 => DATA2(14), A2 => n2355, B1 => n2354, B2 => 
                           n2353, ZN => n2359);
   U1666 : NAND3_X1 port map( A1 => n2357, A2 => n2441, A3 => n2356, ZN => 
                           n2358);
   U1667 : OAI211_X1 port map( C1 => n2683, C2 => n2462, A => n2359, B => n2358
                           , ZN => n2360);
   U1668 : AOI211_X1 port map( C1 => n2363, C2 => n2362, A => n2361, B => n2360
                           , ZN => n2364);
   U1669 : OAI21_X1 port map( B1 => n2365, B2 => n2455, A => n2364, ZN => 
                           OUTALU(14));
   U1670 : AOI222_X1 port map( A1 => n2392, A2 => n2517_port, B1 => n2387, B2 
                           => n2366, C1 => n2389, C2 => n2518_port, ZN => n2382
                           );
   U1671 : NOR2_X1 port map( A1 => n2402, A2 => n2433, ZN => n2368);
   U1672 : INV_X1 port map( A => n2395, ZN => n2367);
   U1673 : OAI211_X1 port map( C1 => n2368, C2 => n2451, A => n2367, B => n2371
                           , ZN => n2381);
   U1674 : OAI21_X1 port map( B1 => n2763, B2 => n2458, A => n2437, ZN => n2379
                           );
   U1675 : AOI21_X1 port map( B1 => n2371, B2 => n2370, A => n2369, ZN => n2378
                           );
   U1676 : AOI22_X1 port map( A1 => n2442, A2 => n2372, B1 => n2506, B2 => 
                           n2386, ZN => n2376);
   U1677 : AOI22_X1 port map( A1 => n2383, A2 => n2409, B1 => n2373, B2 => 
                           n2440, ZN => n2375);
   U1678 : NAND2_X1 port map( A1 => DATA2(13), A2 => n2649, ZN => n2682);
   U1679 : OAI21_X1 port map( B1 => DATA2(13), B2 => n2649, A => n2682, ZN => 
                           n2571);
   U1680 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_13_port, B1 => 
                           n2438, B2 => n2571, ZN => n2374);
   U1681 : OAI221_X1 port map( B1 => n2427, B2 => n2376, C1 => n2427, C2 => 
                           n2375, A => n2374, ZN => n2377);
   U1682 : AOI211_X1 port map( C1 => DATA1(13), C2 => n2379, A => n2378, B => 
                           n2377, ZN => n2380);
   U1683 : OAI211_X1 port map( C1 => n2382, C2 => n2455, A => n2381, B => n2380
                           , ZN => OUTALU(13));
   U1684 : AOI222_X1 port map( A1 => n2386, A2 => n2385, B1 => n2409, B2 => 
                           n2384, C1 => n2440, C2 => n2383, ZN => n2408);
   U1685 : AOI22_X1 port map( A1 => n2514, A2 => n2389, B1 => n2388, B2 => 
                           n2387, ZN => n2394);
   U1686 : AOI22_X1 port map( A1 => n2518_port, A2 => n2392, B1 => n2391, B2 =>
                           n2390, ZN => n2393);
   U1687 : AOI21_X1 port map( B1 => n2394, B2 => n2393, A => n2455, ZN => n2401
                           );
   U1688 : OAI22_X1 port map( A1 => n2681, A2 => DATA2(12), B1 => n2764, B2 => 
                           DATA1(12), ZN => n2680);
   U1689 : INV_X1 port map( A => n2680, ZN => n2614);
   U1690 : OAI211_X1 port map( C1 => n2405, C2 => n2396, A => n2451, B => n2395
                           , ZN => n2399);
   U1691 : OAI211_X1 port map( C1 => n2410, C2 => n2412, A => n2397, B => 
                           DATA2(12), ZN => n2398);
   U1692 : OAI211_X1 port map( C1 => n2614, C2 => n2462, A => n2399, B => n2398
                           , ZN => n2400);
   U1693 : AOI211_X1 port map( C1 => n2449, C2 => dataout_mul_12_port, A => 
                           n2401, B => n2400, ZN => n2407);
   U1694 : OAI211_X1 port map( C1 => n2405, C2 => n2404, A => n2403, B => n2402
                           , ZN => n2406);
   U1695 : OAI211_X1 port map( C1 => n2408, C2 => n2427, A => n2407, B => n2406
                           , ZN => OUTALU(12));
   U1696 : AOI22_X1 port map( A1 => n2442, A2 => n2409, B1 => n2506, B2 => 
                           n2440, ZN => n2428);
   U1697 : AOI221_X1 port map( B1 => n2412, B2 => n2678, C1 => n2438, C2 => 
                           n2411, A => n2410, ZN => n2413);
   U1698 : NAND2_X1 port map( A1 => n2678, A2 => n2765, ZN => n2613);
   U1699 : OAI22_X1 port map( A1 => n2413, A2 => n2765, B1 => n2462, B2 => 
                           n2613, ZN => n2414);
   U1700 : AOI21_X1 port map( B1 => n2449, B2 => dataout_mul_11_port, A => 
                           n2414, ZN => n2426);
   U1701 : INV_X1 port map( A => n2418, ZN => n2416);
   U1702 : XOR2_X1 port map( A => n2416, B => n2415, Z => n2424);
   U1703 : INV_X1 port map( A => n2419, ZN => n2417);
   U1704 : AOI221_X1 port map( B1 => n2419, B2 => n2418, C1 => n2417, C2 => 
                           n2416, A => n2433, ZN => n2423);
   U1705 : NOR3_X1 port map( A1 => n2421, A2 => n2455, A3 => n2420, ZN => n2422
                           );
   U1706 : AOI211_X1 port map( C1 => n2451, C2 => n2424, A => n2423, B => n2422
                           , ZN => n2425);
   U1707 : OAI211_X1 port map( C1 => n2428, C2 => n2427, A => n2426, B => n2425
                           , ZN => OUTALU(11));
   U1708 : AOI22_X1 port map( A1 => n2431, A2 => n2430, B1 => n2526_port, B2 =>
                           n2429, ZN => n2456);
   U1709 : NAND2_X1 port map( A1 => n2451, A2 => n2432, ZN => n2435);
   U1710 : OR2_X1 port map( A1 => n2434, A2 => n2433, ZN => n2446);
   U1711 : AOI22_X1 port map( A1 => n2450, A2 => n2436, B1 => n2435, B2 => 
                           n2446, ZN => n2448);
   U1712 : OAI21_X1 port map( B1 => n2766, B2 => n2458, A => n2437, ZN => n2439
                           );
   U1713 : AOI22_X1 port map( A1 => n2576, A2 => DATA2(10), B1 => n2766, B2 => 
                           n2561, ZN => n2672);
   U1714 : AOI22_X1 port map( A1 => n2576, A2 => n2439, B1 => n2438, B2 => 
                           n2672, ZN => n2444);
   U1715 : NAND3_X1 port map( A1 => n2442, A2 => n2441, A3 => n2440, ZN => 
                           n2443);
   U1716 : OAI211_X1 port map( C1 => n2446, C2 => n2445, A => n2444, B => n2443
                           , ZN => n2447);
   U1717 : AOI211_X1 port map( C1 => n2449, C2 => dataout_mul_10_port, A => 
                           n2448, B => n2447, ZN => n2454);
   U1718 : NAND3_X1 port map( A1 => n2452, A2 => n2451, A3 => n2450, ZN => 
                           n2453);
   U1719 : OAI211_X1 port map( C1 => n2456, C2 => n2455, A => n2454, B => n2453
                           , ZN => OUTALU(10));
   U1720 : OAI21_X1 port map( B1 => n2778, B2 => n2458, A => n2457, ZN => n2465
                           );
   U1721 : OAI22_X1 port map( A1 => n2778, A2 => DATA1(0), B1 => n2650, B2 => 
                           DATA2(0), ZN => n2559);
   U1722 : INV_X1 port map( A => n2559, ZN => n2463);
   U1723 : NOR2_X1 port map( A1 => n2460, A2 => n2459, ZN => n2467);
   U1724 : OAI22_X1 port map( A1 => n2463, A2 => n2462, B1 => n2467, B2 => 
                           n2461, ZN => n2464);
   U1725 : AOI21_X1 port map( B1 => DATA1(0), B2 => n2465, A => n2464, ZN => 
                           n2742);
   U1726 : AOI22_X1 port map( A1 => n2468, A2 => dataout_mul_0_port, B1 => 
                           n2467, B2 => n2466, ZN => n2741);
   U1727 : INV_X1 port map( A => n2469, ZN => n2536_port);
   U1728 : INV_X1 port map( A => n2470, ZN => n2507);
   U1729 : INV_X1 port map( A => n2471, ZN => n2495);
   U1730 : OAI211_X1 port map( C1 => n2474, C2 => n2650, A => n2473, B => n2472
                           , ZN => n2475);
   U1731 : AOI211_X1 port map( C1 => DATA1(4), C2 => n2477, A => n2476, B => 
                           n2475, ZN => n2478);
   U1732 : INV_X1 port map( A => n2478, ZN => n2482);
   U1733 : AOI222_X1 port map( A1 => n2483, A2 => n2482, B1 => n1626, B2 => 
                           n2481, C1 => n2480, C2 => n2479, ZN => n2484);
   U1734 : OAI22_X1 port map( A1 => n2487, A2 => n2486, B1 => n2485, B2 => 
                           n2484, ZN => n2493);
   U1735 : OAI22_X1 port map( A1 => n2491, A2 => n2490, B1 => n2489, B2 => 
                           n2488, ZN => n2492);
   U1736 : AOI211_X1 port map( C1 => n2495, C2 => n2494, A => n2493, B => n2492
                           , ZN => n2498);
   U1737 : OAI22_X1 port map( A1 => n2499, A2 => n2498, B1 => n2497, B2 => 
                           n2496, ZN => n2505);
   U1738 : OAI22_X1 port map( A1 => n2503, A2 => n2502, B1 => n2501, B2 => 
                           n2500, ZN => n2504);
   U1739 : AOI211_X1 port map( C1 => n2507, C2 => n2506, A => n2505, B => n2504
                           , ZN => n2509);
   U1740 : OAI222_X1 port map( A1 => n2513, A2 => n2512, B1 => n2511, B2 => 
                           n2510, C1 => n2509, C2 => n2508, ZN => n2516);
   U1741 : AOI22_X1 port map( A1 => n2517_port, A2 => n2516, B1 => n2515, B2 =>
                           n2514, ZN => n2523_port);
   U1742 : AOI22_X1 port map( A1 => n2521_port, A2 => n2520_port, B1 => 
                           n2519_port, B2 => n2518_port, ZN => n2522_port);
   U1743 : OAI211_X1 port map( C1 => n2525_port, C2 => n2524_port, A => 
                           n2523_port, B => n2522_port, ZN => n2527_port);
   U1744 : AOI22_X1 port map( A1 => n2529_port, A2 => n2528_port, B1 => 
                           n2527_port, B2 => n2526_port, ZN => n2535_port);
   U1745 : AOI22_X1 port map( A1 => n2533_port, A2 => n2532_port, B1 => 
                           n2531_port, B2 => n2530_port, ZN => n2534_port);
   U1746 : OAI211_X1 port map( C1 => n2537_port, C2 => n2536_port, A => 
                           n2535_port, B => n2534_port, ZN => n2540_port);
   U1747 : AOI222_X1 port map( A1 => n2543_port, A2 => n2542_port, B1 => 
                           n2541_port, B2 => n2540_port, C1 => n2539_port, C2 
                           => n2538_port, ZN => n2544_port);
   U1748 : INV_X1 port map( A => n2544_port, ZN => n2547_port);
   U1749 : AOI22_X1 port map( A1 => n2548_port, A2 => n2547_port, B1 => 
                           n2546_port, B2 => n2545_port, ZN => n2554);
   U1750 : AOI22_X1 port map( A1 => n2552, A2 => n2551, B1 => n2550, B2 => 
                           n2549, ZN => n2553);
   U1751 : OAI211_X1 port map( C1 => n2556, C2 => n2555, A => n2554, B => n2553
                           , ZN => n2735);
   U1752 : OAI21_X1 port map( B1 => DATA2(26), B2 => n2557, A => n2641, ZN => 
                           n2719);
   U1753 : AOI22_X1 port map( A1 => n2646, A2 => DATA2(31), B1 => n2746, B2 => 
                           DATA1(30), ZN => n2729);
   U1754 : INV_X1 port map( A => n2729, ZN => n2560);
   U1755 : NOR4_X1 port map( A1 => n2719, A2 => n2560, A3 => n2559, A4 => n2558
                           , ZN => n2575);
   U1756 : OAI21_X1 port map( B1 => DATA2(10), B2 => n2561, A => n2613, ZN => 
                           n2676);
   U1757 : INV_X1 port map( A => n2676, ZN => n2563);
   U1758 : AOI22_X1 port map( A1 => n2762, A2 => DATA1(14), B1 => n2761, B2 => 
                           n3098, ZN => n2689);
   U1759 : AOI21_X1 port map( B1 => n2758, B2 => DATA1(18), A => n2562, ZN => 
                           n2699);
   U1760 : AOI22_X1 port map( A1 => n2754, A2 => DATA1(22), B1 => n2753, B2 => 
                           DATA1(23), ZN => n2708);
   U1761 : AND4_X1 port map( A1 => n2563, A2 => n2689, A3 => n2699, A4 => n2708
                           , ZN => n2574);
   U1762 : NOR4_X1 port map( A1 => n2567, A2 => n2566, A3 => n2565, A4 => n2564
                           , ZN => n2573);
   U1763 : NOR4_X1 port map( A1 => n2571, A2 => n2570, A3 => n2569, A4 => n2568
                           , ZN => n2572);
   U1764 : NAND4_X1 port map( A1 => n2575, A2 => n2574, A3 => n2573, A4 => 
                           n2572, ZN => n2591);
   U1765 : OAI22_X1 port map( A1 => n2766, A2 => n2576, B1 => n2765, B2 => 
                           DATA1(11), ZN => n2615);
   U1766 : AOI22_X1 port map( A1 => DATA2(14), A2 => n2578, B1 => DATA2(15), B2
                           => n2577, ZN => n2621);
   U1767 : INV_X1 port map( A => n2621, ZN => n2579);
   U1768 : OR4_X1 port map( A1 => n2615, A2 => n2680, A3 => n2579, A4 => n2686,
                           ZN => n2589);
   U1769 : AOI22_X1 port map( A1 => DATA2(6), A2 => n2580, B1 => DATA2(7), B2 
                           => n2667, ZN => n2607);
   U1770 : INV_X1 port map( A => n2604, ZN => n2671);
   U1771 : NAND4_X1 port map( A1 => n2653, A2 => n2597, A3 => n2607, A4 => 
                           n2671, ZN => n2588);
   U1772 : OAI21_X1 port map( B1 => n2750, B2 => DATA1(26), A => n2717, ZN => 
                           n2642);
   U1773 : INV_X1 port map( A => n2642, ZN => n2583);
   U1774 : AOI21_X1 port map( B1 => DATA2(30), B2 => n2581, A => n2727, ZN => 
                           n2648);
   U1775 : AOI21_X1 port map( B1 => n2582, B2 => n2772, A => n2605, ZN => n2669
                           );
   U1776 : NAND4_X1 port map( A1 => n2583, A2 => n2718, A3 => n2648, A4 => 
                           n2669, ZN => n2587);
   U1777 : AOI21_X1 port map( B1 => DATA2(18), B2 => n2584, A => n2697, ZN => 
                           n2585);
   U1778 : INV_X1 port map( A => n2585, ZN => n2628);
   U1779 : OAI22_X1 port map( A1 => n2753, A2 => DATA1(23), B1 => n2754, B2 => 
                           DATA1(22), ZN => n2636);
   U1780 : OR4_X1 port map( A1 => n2628, A2 => n2696, A3 => n2636, A4 => n2706,
                           ZN => n2586);
   U1781 : OR4_X1 port map( A1 => n2589, A2 => n2588, A3 => n2587, A4 => n2586,
                           ZN => n2590);
   U1782 : OAI21_X1 port map( B1 => n2591, B2 => n2590, A => n2743, ZN => n2593
                           );
   U1783 : INV_X1 port map( A => FUNC(0), ZN => n2592);
   U1784 : AOI211_X1 port map( C1 => FUNC(2), C2 => n2593, A => FUNC(1), B => 
                           n2592, ZN => n2734);
   U1785 : AOI22_X1 port map( A1 => DATA2(25), A2 => n2716, B1 => DATA2(24), B2
                           => n2709, ZN => n2640);
   U1786 : AOI22_X1 port map( A1 => DATA2(21), A2 => n2700, B1 => DATA2(20), B2
                           => n2701, ZN => n2633);
   U1787 : OAI21_X1 port map( B1 => DATA2(1), B2 => n2651, A => DATA2(0), ZN =>
                           n2594);
   U1788 : OAI22_X1 port map( A1 => DATA1(0), A2 => n2594, B1 => DATA1(1), B2 
                           => n2777, ZN => n2595);
   U1789 : AOI22_X1 port map( A1 => DATA2(2), A2 => n2658, B1 => n2653, B2 => 
                           n2595, ZN => n2596);
   U1790 : INV_X1 port map( A => n2596, ZN => n2598);
   U1791 : NOR2_X1 port map( A1 => n2775, A2 => DATA1(3), ZN => n2662);
   U1792 : NAND2_X1 port map( A1 => n2775, A2 => DATA1(3), ZN => n2656);
   U1793 : OAI211_X1 port map( C1 => n2598, C2 => n2662, A => n2656, B => n2597
                           , ZN => n2599);
   U1794 : INV_X1 port map( A => n2599, ZN => n2603);
   U1795 : NAND2_X1 port map( A1 => DATA2(5), A2 => n2600, ZN => n2663);
   U1796 : OAI21_X1 port map( B1 => DATA1(4), B2 => n2774, A => n2663, ZN => 
                           n2602);
   U1797 : NOR2_X1 port map( A1 => n2600, A2 => DATA2(5), ZN => n2666);
   U1798 : INV_X1 port map( A => n2666, ZN => n2601);
   U1799 : OAI211_X1 port map( C1 => n2603, C2 => n2602, A => n2664, B => n2601
                           , ZN => n2606);
   U1800 : AOI211_X1 port map( C1 => n2607, C2 => n2606, A => n2605, B => n2604
                           , ZN => n2608);
   U1801 : AOI21_X1 port map( B1 => DATA2(8), B2 => n2609, A => n2608, ZN => 
                           n2612);
   U1802 : INV_X1 port map( A => n2674, ZN => n2610);
   U1803 : AOI211_X1 port map( C1 => n2612, C2 => n2611, A => n2610, B => n2672
                           , ZN => n2616);
   U1804 : OAI211_X1 port map( C1 => n2616, C2 => n2615, A => n2614, B => n2613
                           , ZN => n2617);
   U1805 : OAI211_X1 port map( C1 => DATA1(12), C2 => n2764, A => n2617, B => 
                           n2682, ZN => n2618);
   U1806 : OAI211_X1 port map( C1 => DATA2(13), C2 => n2649, A => n2683, B => 
                           n2618, ZN => n2620);
   U1807 : AOI211_X1 port map( C1 => n2621, C2 => n2620, A => n2619, B => n2686
                           , ZN => n2622);
   U1808 : AOI21_X1 port map( B1 => DATA2(16), B2 => n2691, A => n2622, ZN => 
                           n2625);
   U1809 : AOI211_X1 port map( C1 => n2625, C2 => n2692, A => n2624, B => n2623
                           , ZN => n2629);
   U1810 : INV_X1 port map( A => n2696, ZN => n2627);
   U1811 : OAI211_X1 port map( C1 => n2629, C2 => n2628, A => n2627, B => n2626
                           , ZN => n2632);
   U1812 : NOR2_X1 port map( A1 => DATA2(21), A2 => n2700, ZN => n2631);
   U1813 : AOI211_X1 port map( C1 => n2633, C2 => n2632, A => n2631, B => n2630
                           , ZN => n2637);
   U1814 : INV_X1 port map( A => n2706, ZN => n2635);
   U1815 : OAI211_X1 port map( C1 => n2637, C2 => n2636, A => n2635, B => n2634
                           , ZN => n2639);
   U1816 : NOR2_X1 port map( A1 => DATA2(25), A2 => n2716, ZN => n2711);
   U1817 : INV_X1 port map( A => n2638, ZN => n2714);
   U1818 : AOI211_X1 port map( C1 => n2640, C2 => n2639, A => n2711, B => n2714
                           , ZN => n2643);
   U1819 : OAI211_X1 port map( C1 => n2643, C2 => n2642, A => n2718, B => n2641
                           , ZN => n2644);
   U1820 : OAI211_X1 port map( C1 => DATA1(28), C2 => n2748, A => n2644, B => 
                           n2725, ZN => n2645);
   U1821 : NAND3_X1 port map( A1 => n2726, A2 => n2722, A3 => n2645, ZN => 
                           n2647);
   U1822 : AOI22_X1 port map( A1 => n2648, A2 => n2647, B1 => DATA2(31), B2 => 
                           n2646, ZN => n2732);
   U1823 : NOR2_X1 port map( A1 => DATA2(13), A2 => n2649, ZN => n2685);
   U1824 : NOR2_X1 port map( A1 => DATA2(0), A2 => n2650, ZN => n2655);
   U1825 : NOR2_X1 port map( A1 => DATA2(1), A2 => n2651, ZN => n2654);
   U1826 : NAND2_X1 port map( A1 => DATA2(1), A2 => n2651, ZN => n2652);
   U1827 : OAI211_X1 port map( C1 => n2655, C2 => n2654, A => n2653, B => n2652
                           , ZN => n2657);
   U1828 : OAI211_X1 port map( C1 => DATA2(2), C2 => n2658, A => n2657, B => 
                           n2656, ZN => n2659);
   U1829 : OAI21_X1 port map( B1 => DATA1(4), B2 => n2774, A => n2659, ZN => 
                           n2661);
   U1830 : OAI22_X1 port map( A1 => n2662, A2 => n2661, B1 => DATA2(4), B2 => 
                           n2660, ZN => n2665);
   U1831 : OAI211_X1 port map( C1 => n2666, C2 => n2665, A => n2664, B => n2663
                           , ZN => n2668);
   U1832 : AOI22_X1 port map( A1 => n2669, A2 => n2668, B1 => DATA2(7), B2 => 
                           n2667, ZN => n2670);
   U1833 : AOI22_X1 port map( A1 => DATA1(8), A2 => n2768, B1 => n2671, B2 => 
                           n2670, ZN => n2675);
   U1834 : AOI211_X1 port map( C1 => n2675, C2 => n2674, A => n2673, B => n2672
                           , ZN => n2677);
   U1835 : OAI22_X1 port map( A1 => n2678, A2 => n2765, B1 => n2677, B2 => 
                           n2676, ZN => n2679);
   U1836 : OAI22_X1 port map( A1 => DATA2(12), A2 => n2681, B1 => n2680, B2 => 
                           n2679, ZN => n2684);
   U1837 : OAI211_X1 port map( C1 => n2685, C2 => n2684, A => n2683, B => n2682
                           , ZN => n2688);
   U1838 : AOI211_X1 port map( C1 => n2689, C2 => n2688, A => n2687, B => n2686
                           , ZN => n2695);
   U1839 : OAI21_X1 port map( B1 => DATA2(16), B2 => n2691, A => n2690, ZN => 
                           n2694);
   U1840 : OAI211_X1 port map( C1 => n2695, C2 => n2694, A => n2693, B => n2692
                           , ZN => n2698);
   U1841 : AOI211_X1 port map( C1 => n2699, C2 => n2698, A => n2697, B => n2696
                           , ZN => n2705);
   U1842 : OAI22_X1 port map( A1 => DATA2(20), A2 => n2701, B1 => DATA2(21), B2
                           => n2700, ZN => n2704);
   U1843 : OAI211_X1 port map( C1 => n2705, C2 => n2704, A => n2703, B => n2702
                           , ZN => n2707);
   U1844 : AOI21_X1 port map( B1 => n2708, B2 => n2707, A => n2706, ZN => n2713
                           );
   U1845 : NOR2_X1 port map( A1 => DATA2(24), A2 => n2709, ZN => n2710);
   U1846 : AOI211_X1 port map( C1 => n2713, C2 => n2712, A => n2711, B => n2710
                           , ZN => n2715);
   U1847 : AOI211_X1 port map( C1 => DATA2(25), C2 => n2716, A => n2715, B => 
                           n2714, ZN => n2720);
   U1848 : OAI211_X1 port map( C1 => n2720, C2 => n2719, A => n2718, B => n2717
                           , ZN => n2721);
   U1849 : OAI211_X1 port map( C1 => DATA2(28), C2 => n2723, A => n2722, B => 
                           n2721, ZN => n2724);
   U1850 : NAND3_X1 port map( A1 => n2726, A2 => n2725, A3 => n2724, ZN => 
                           n2728);
   U1851 : AOI21_X1 port map( B1 => n2729, B2 => n2728, A => n2727, ZN => n2731
                           );
   U1852 : OAI221_X1 port map( B1 => FUNC(3), B2 => n2732, C1 => n2743, C2 => 
                           n2731, A => n2730, ZN => n2733);
   U1853 : AOI22_X1 port map( A1 => n2736, A2 => n2735, B1 => n2734, B2 => 
                           n2733, ZN => n2740);
   U1854 : NAND3_X1 port map( A1 => n2738, A2 => FUNC(3), A3 => n2737, ZN => 
                           n2739);
   U1855 : NAND4_X1 port map( A1 => n2742, A2 => n2741, A3 => n2740, A4 => 
                           n2739, ZN => OUTALU(0));
   U1856 : NAND2_X1 port map( A1 => n2744, A2 => n2743, ZN => n2780);
   U1857 : CLKBUF_X1 port map( A => n2780, Z => n2770);
   U1858 : NAND2_X1 port map( A1 => FUNC(3), A2 => n2744, ZN => n2779);
   U1859 : INV_X1 port map( A => DATA2(31), ZN => n2745);
   U1860 : AOI22_X1 port map( A1 => DATA2(31), A2 => n2770, B1 => n2769, B2 => 
                           n2745, ZN => N2548);
   U1861 : AOI22_X1 port map( A1 => DATA2(30), A2 => n2780, B1 => n2779, B2 => 
                           n2746, ZN => N2547);
   U1862 : AOI22_X1 port map( A1 => DATA2(29), A2 => n2770, B1 => n2769, B2 => 
                           n2747, ZN => N2546);
   U1863 : AOI22_X1 port map( A1 => DATA2(28), A2 => n2780, B1 => n2779, B2 => 
                           n2748, ZN => N2545);
   U1864 : AOI22_X1 port map( A1 => DATA2(27), A2 => n2770, B1 => n2769, B2 => 
                           n2749, ZN => N2544);
   U1865 : AOI22_X1 port map( A1 => DATA2(26), A2 => n2780, B1 => n2779, B2 => 
                           n2750, ZN => N2543);
   U1866 : INV_X1 port map( A => DATA2(25), ZN => n2751);
   U1867 : AOI22_X1 port map( A1 => DATA2(25), A2 => n2770, B1 => n2769, B2 => 
                           n2751, ZN => N2542);
   U1868 : AOI22_X1 port map( A1 => DATA2(24), A2 => n2780, B1 => n2779, B2 => 
                           n2752, ZN => N2541);
   U1869 : AOI22_X1 port map( A1 => DATA2(23), A2 => n2770, B1 => n2769, B2 => 
                           n2753, ZN => N2540);
   U1870 : AOI22_X1 port map( A1 => DATA2(22), A2 => n2780, B1 => n2779, B2 => 
                           n2754, ZN => N2539);
   U1871 : INV_X1 port map( A => DATA2(21), ZN => n2755);
   U1872 : AOI22_X1 port map( A1 => DATA2(21), A2 => n2780, B1 => n2779, B2 => 
                           n2755, ZN => N2538);
   U1873 : AOI22_X1 port map( A1 => DATA2(20), A2 => n2780, B1 => n2779, B2 => 
                           n2756, ZN => N2537);
   U1874 : AOI22_X1 port map( A1 => DATA2(19), A2 => n2770, B1 => n2769, B2 => 
                           n2757, ZN => N2536);
   U1875 : AOI22_X1 port map( A1 => DATA2(18), A2 => n2770, B1 => n2769, B2 => 
                           n2758, ZN => N2535);
   U1876 : INV_X1 port map( A => DATA2(17), ZN => n2759);
   U1877 : AOI22_X1 port map( A1 => DATA2(17), A2 => n2770, B1 => n2769, B2 => 
                           n2759, ZN => N2534);
   U1878 : AOI22_X1 port map( A1 => DATA2(16), A2 => n2770, B1 => n2769, B2 => 
                           n2760, ZN => N2533);
   U1879 : AOI22_X1 port map( A1 => DATA2(15), A2 => n2770, B1 => n2769, B2 => 
                           n2761, ZN => N2532);
   U1880 : AOI22_X1 port map( A1 => DATA2(14), A2 => n2770, B1 => n2769, B2 => 
                           n2762, ZN => N2531);
   U1881 : AOI22_X1 port map( A1 => DATA2(13), A2 => n2770, B1 => n2769, B2 => 
                           n2763, ZN => N2530);
   U1882 : AOI22_X1 port map( A1 => DATA2(12), A2 => n2770, B1 => n2769, B2 => 
                           n2764, ZN => N2529);
   U1883 : AOI22_X1 port map( A1 => DATA2(11), A2 => n2770, B1 => n2769, B2 => 
                           n2765, ZN => N2528);
   U1884 : AOI22_X1 port map( A1 => DATA2(10), A2 => n2770, B1 => n2769, B2 => 
                           n2766, ZN => N2527);
   U1885 : AOI22_X1 port map( A1 => DATA2(9), A2 => n2770, B1 => n2769, B2 => 
                           n2767, ZN => N2526);
   U1886 : AOI22_X1 port map( A1 => DATA2(8), A2 => n2770, B1 => n2769, B2 => 
                           n2768, ZN => N2525);
   U1887 : INV_X1 port map( A => DATA2(7), ZN => n2771);
   U1888 : AOI22_X1 port map( A1 => DATA2(7), A2 => n2780, B1 => n2779, B2 => 
                           n2771, ZN => N2524);
   U1889 : AOI22_X1 port map( A1 => DATA2(6), A2 => n2780, B1 => n2779, B2 => 
                           n2772, ZN => N2523);
   U1890 : AOI22_X1 port map( A1 => DATA2(5), A2 => n2780, B1 => n2779, B2 => 
                           n2773, ZN => N2522);
   U1891 : AOI22_X1 port map( A1 => DATA2(4), A2 => n2780, B1 => n2779, B2 => 
                           n2774, ZN => N2521);
   U1892 : AOI22_X1 port map( A1 => DATA2(3), A2 => n2780, B1 => n2779, B2 => 
                           n2775, ZN => N2520);
   U1893 : AOI22_X1 port map( A1 => DATA2(2), A2 => n2780, B1 => n2779, B2 => 
                           n2776, ZN => N2519);
   U1894 : AOI22_X1 port map( A1 => DATA2(1), A2 => n2780, B1 => n2779, B2 => 
                           n2777, ZN => N2518);
   U1895 : AOI22_X1 port map( A1 => DATA2(0), A2 => n2780, B1 => n2779, B2 => 
                           n2778, ZN => N2517);
   U1896 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           A2 => n2781, ZN => 
                           boothmul_pipelined_i_sum_out_1_0_port);
   U1897 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN
                           => n2783);
   U1898 : NAND2_X1 port map( A1 => data2_mul_3_port, A2 => n2783, ZN => n2819)
                           ;
   U1899 : INV_X1 port map( A => data2_mul_3_port, ZN => n2817);
   U1900 : NAND3_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, 
                           A3 => n2817, ZN => n2816);
   U1901 : NOR2_X1 port map( A1 => n2817, A2 => n2782, ZN => n2818);
   U1902 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2818, B1 => data1_mul_1_port, B2 => n2811, ZN
                           => n2784);
   U1903 : OAI221_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           B2 => n2819, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           C2 => n2816, A => n2784, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1904 : CLKBUF_X1 port map( A => n2818, Z => n2812);
   U1905 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           n2811, B2 => data1_mul_2_port, ZN => n2786);
   U1906 : INV_X1 port map( A => n2819, ZN => n2813);
   U1907 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2813, ZN => n2785);
   U1908 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, 
                           C2 => n2816, A => n2786, B => n2785, ZN => 
                           boothmul_pipelined_i_mux_out_1_4_port);
   U1909 : AOI22_X1 port map( A1 => n2818, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B1 => 
                           n2811, B2 => data1_mul_3_port, ZN => n2788);
   U1910 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, ZN => 
                           n2787);
   U1911 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, 
                           C2 => n2816, A => n2788, B => n2787, ZN => 
                           boothmul_pipelined_i_mux_out_1_5_port);
   U1912 : AOI22_X1 port map( A1 => n2818, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n2811, B2 => data1_mul_4_port, ZN => n2790);
   U1913 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n2789);
   U1914 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, 
                           C2 => n2816, A => n2790, B => n2789, ZN => 
                           boothmul_pipelined_i_mux_out_1_6_port);
   U1915 : AOI22_X1 port map( A1 => n2818, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n2811, B2 => data1_mul_5_port, ZN => n2792);
   U1916 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n2791);
   U1917 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, 
                           C2 => n2816, A => n2792, B => n2791, ZN => 
                           boothmul_pipelined_i_mux_out_1_7_port);
   U1918 : AOI22_X1 port map( A1 => n2818, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n2811, B2 => data1_mul_6_port, ZN => n2794);
   U1919 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n2793);
   U1920 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, 
                           C2 => n2816, A => n2794, B => n2793, ZN => 
                           boothmul_pipelined_i_mux_out_1_8_port);
   U1921 : AOI22_X1 port map( A1 => n2818, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n2811, B2 => data1_mul_7_port, ZN => n2796);
   U1922 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n2795);
   U1923 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, 
                           C2 => n2816, A => n2796, B => n2795, ZN => 
                           boothmul_pipelined_i_mux_out_1_9_port);
   U1924 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n2811, B2 => data1_mul_8_port, ZN => n2798);
   U1925 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n2797);
   U1926 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, 
                           C2 => n2816, A => n2798, B => n2797, ZN => 
                           boothmul_pipelined_i_mux_out_1_10_port);
   U1927 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n2811, B2 => data1_mul_9_port, ZN => n2800);
   U1928 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n2799);
   U1929 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, 
                           C2 => n2816, A => n2800, B => n2799, ZN => 
                           boothmul_pipelined_i_mux_out_1_11_port);
   U1930 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n2811, B2 => data1_mul_10_port, ZN => n2802);
   U1931 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n2801);
   U1932 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, 
                           C2 => n2816, A => n2802, B => n2801, ZN => 
                           boothmul_pipelined_i_mux_out_1_12_port);
   U1933 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n2811, B2 => data1_mul_11_port, ZN => n2804);
   U1934 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n2803);
   U1935 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, 
                           C2 => n2816, A => n2804, B => n2803, ZN => 
                           boothmul_pipelined_i_mux_out_1_13_port);
   U1936 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n2811, B2 => data1_mul_12_port, ZN => n2806);
   U1937 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n2805);
   U1938 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, 
                           C2 => n2816, A => n2806, B => n2805, ZN => 
                           boothmul_pipelined_i_mux_out_1_14_port);
   U1939 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n2811, B2 => data1_mul_13_port, ZN => n2808);
   U1940 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n2807);
   U1941 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, 
                           C2 => n2816, A => n2808, B => n2807, ZN => 
                           boothmul_pipelined_i_mux_out_1_15_port);
   U1942 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n2811, B2 => data1_mul_14_port, ZN => n2810);
   U1943 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n2809);
   U1944 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, 
                           C2 => n2816, A => n2810, B => n2809, ZN => 
                           boothmul_pipelined_i_mux_out_1_16_port);
   U1945 : AOI22_X1 port map( A1 => n2812, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n2811, B2 => data1_mul_15_port, ZN => n2815);
   U1946 : NAND2_X1 port map( A1 => n2813, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n2814);
   U1947 : OAI211_X1 port map( C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, 
                           C2 => n2816, A => n2815, B => n2814, ZN => 
                           boothmul_pipelined_i_mux_out_1_17_port);
   U1948 : OAI21_X1 port map( B1 => data2_mul_1_port, B2 => data2_mul_2_port, A
                           => n2817, ZN => n2821);
   U1949 : INV_X1 port map( A => n2818, ZN => n2820);
   U1950 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_119_port, ZN 
                           => n2859);
   U1951 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_102_port, ZN 
                           => n2861);
   U1952 : OAI222_X1 port map( A1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           A2 => n2821, B1 => n2820, B2 => n2859, C1 => n2819, 
                           C2 => n2861, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1953 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n2823);
   U1954 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n2823, ZN => n2862);
   U1955 : NAND3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           A3 => n3076, ZN => n2856);
   U1956 : NOR2_X1 port map( A1 => n3076, A2 => n2822, ZN => n2857);
   U1957 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2857, B1 => data1_mul_1_port, B2 => n2852, ZN
                           => n2824);
   U1958 : OAI221_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           B2 => n2862, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           C2 => n2856, A => n2824, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1959 : CLKBUF_X1 port map( A => n2857, Z => n2851);
   U1960 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B2 => 
                           n2851, ZN => n2826);
   U1961 : INV_X1 port map( A => n2862, ZN => n2853);
   U1962 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n2853, ZN => n2825);
   U1963 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, A 
                           => n2826, B => n2825, ZN => 
                           boothmul_pipelined_i_mux_out_2_6_port);
   U1964 : AOI22_X1 port map( A1 => data1_mul_3_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n2857, ZN => n2828);
   U1965 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n2853, ZN => n2827);
   U1966 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_2_port, A 
                           => n2828, B => n2827, ZN => 
                           boothmul_pipelined_i_mux_out_2_7_port);
   U1967 : AOI22_X1 port map( A1 => data1_mul_4_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n2857, ZN => n2830);
   U1968 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n2853, ZN => n2829);
   U1969 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, A 
                           => n2830, B => n2829, ZN => 
                           boothmul_pipelined_i_mux_out_2_8_port);
   U1970 : AOI22_X1 port map( A1 => data1_mul_5_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n2857, ZN => n2832);
   U1971 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n2853, ZN => n2831);
   U1972 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, A 
                           => n2832, B => n2831, ZN => 
                           boothmul_pipelined_i_mux_out_2_9_port);
   U1973 : AOI22_X1 port map( A1 => data1_mul_6_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n2857, ZN => n2834);
   U1974 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n2853, ZN => n2833);
   U1975 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, A 
                           => n2834, B => n2833, ZN => 
                           boothmul_pipelined_i_mux_out_2_10_port);
   U1976 : AOI22_X1 port map( A1 => data1_mul_7_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n2857, ZN => n2836);
   U1977 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n2853, ZN => n2835);
   U1978 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, A 
                           => n2836, B => n2835, ZN => 
                           boothmul_pipelined_i_mux_out_2_11_port);
   U1979 : AOI22_X1 port map( A1 => data1_mul_8_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n2851, ZN => n2838);
   U1980 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n2853, ZN => n2837);
   U1981 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, A 
                           => n2838, B => n2837, ZN => 
                           boothmul_pipelined_i_mux_out_2_12_port);
   U1982 : AOI22_X1 port map( A1 => data1_mul_9_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n2851, ZN => n2840);
   U1983 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n2853, ZN => n2839);
   U1984 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, A 
                           => n2840, B => n2839, ZN => 
                           boothmul_pipelined_i_mux_out_2_13_port);
   U1985 : AOI22_X1 port map( A1 => data1_mul_10_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n2851, ZN => n2842);
   U1986 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n2853, ZN => n2841);
   U1987 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, A 
                           => n2842, B => n2841, ZN => 
                           boothmul_pipelined_i_mux_out_2_14_port);
   U1988 : AOI22_X1 port map( A1 => data1_mul_11_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n2851, ZN => n2844);
   U1989 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n2853, ZN => n2843);
   U1990 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, A 
                           => n2844, B => n2843, ZN => 
                           boothmul_pipelined_i_mux_out_2_15_port);
   U1991 : AOI22_X1 port map( A1 => data1_mul_12_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n2851, ZN => n2846);
   U1992 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n2853, ZN => n2845);
   U1993 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, A 
                           => n2846, B => n2845, ZN => 
                           boothmul_pipelined_i_mux_out_2_16_port);
   U1994 : AOI22_X1 port map( A1 => data1_mul_13_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n2851, ZN => n2848);
   U1995 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n2853, ZN => n2847);
   U1996 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, A 
                           => n2848, B => n2847, ZN => 
                           boothmul_pipelined_i_mux_out_2_17_port);
   U1997 : AOI22_X1 port map( A1 => data1_mul_14_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n2851, ZN => n2850);
   U1998 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n2853, ZN => n2849);
   U1999 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, A 
                           => n2850, B => n2849, ZN => 
                           boothmul_pipelined_i_mux_out_2_18_port);
   U2000 : AOI22_X1 port map( A1 => data1_mul_15_port, A2 => n2852, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n2851, ZN => n2855);
   U2001 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n2853, ZN => n2854);
   U2002 : OAI211_X1 port map( C1 => n2856, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, A 
                           => n2855, B => n2854, ZN => 
                           boothmul_pipelined_i_mux_out_2_19_port);
   U2003 : INV_X1 port map( A => n2857, ZN => n2860);
   U2004 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n3076, ZN => n2858);
   U2005 : OAI222_X1 port map( A1 => n2862, A2 => n2861, B1 => n2860, B2 => 
                           n2859, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           C2 => n2858, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U2006 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_60_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_176_port, ZN
                           => n2863);
   U2007 : OAI221_X1 port map( B1 => n3077, B2 => n2865, C1 => n3077, C2 => 
                           n2864, A => n2863, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U2008 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_3_60_port, A2
                           => n2895, B1 => n2894, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n2867);
   U2009 : AOI22_X1 port map( A1 => n2879, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n2878
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n2866);
   U2010 : NAND2_X1 port map( A1 => n2867, A2 => n2866, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U2011 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n2869);
   U2012 : AOI22_X1 port map( A1 => n2879, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n2878
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n2868);
   U2013 : NAND2_X1 port map( A1 => n2869, A2 => n2868, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U2014 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n2871);
   U2015 : AOI22_X1 port map( A1 => n2879, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n2878
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n2870);
   U2016 : NAND2_X1 port map( A1 => n2871, A2 => n2870, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U2017 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n2873);
   U2018 : AOI22_X1 port map( A1 => n2879, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n2878
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n2872);
   U2019 : NAND2_X1 port map( A1 => n2873, A2 => n2872, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U2020 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n2875);
   U2021 : AOI22_X1 port map( A1 => n2879, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n2878
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n2874);
   U2022 : NAND2_X1 port map( A1 => n2875, A2 => n2874, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U2023 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n2877);
   U2024 : AOI22_X1 port map( A1 => n2879, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n2878
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n2876);
   U2025 : NAND2_X1 port map( A1 => n2877, A2 => n2876, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U2026 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n2881);
   U2027 : AOI22_X1 port map( A1 => n2879, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n2878
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n2880);
   U2028 : NAND2_X1 port map( A1 => n2881, A2 => n2880, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U2029 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n2883);
   U2030 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n2882);
   U2031 : NAND2_X1 port map( A1 => n2883, A2 => n2882, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U2032 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n2885);
   U2033 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n2884);
   U2034 : NAND2_X1 port map( A1 => n2885, A2 => n2884, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U2035 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n2887);
   U2036 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n2886);
   U2037 : NAND2_X1 port map( A1 => n2887, A2 => n2886, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U2038 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n2889);
   U2039 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n2888);
   U2040 : NAND2_X1 port map( A1 => n2889, A2 => n2888, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U2041 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n2891);
   U2042 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n2890);
   U2043 : NAND2_X1 port map( A1 => n2891, A2 => n2890, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U2044 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n2893);
   U2045 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n2892);
   U2046 : NAND2_X1 port map( A1 => n2893, A2 => n2892, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U2047 : AOI22_X1 port map( A1 => n2895, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n2894
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n2899);
   U2048 : AOI22_X1 port map( A1 => n2897, A2 => 
                           boothmul_pipelined_i_muxes_in_3_46_port, B1 => n2896
                           , B2 => boothmul_pipelined_i_muxes_in_3_162_port, ZN
                           => n2898);
   U2049 : NAND2_X1 port map( A1 => n2899, A2 => n2898, ZN => 
                           boothmul_pipelined_i_mux_out_3_21_port);
   U2050 : CLKBUF_X1 port map( A => n2912, Z => n2933);
   U2051 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_65_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_65_port, ZN 
                           => n2901);
   U2052 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_190_port, ZN
                           => n2900);
   U2053 : NAND2_X1 port map( A1 => n2901, A2 => n2900, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U2054 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_64_port, A2
                           => n2912, B1 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, B2 => 
                           n2932, ZN => n2903);
   U2055 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n2902);
   U2056 : NAND2_X1 port map( A1 => n2903, A2 => n2902, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U2057 : AOI22_X1 port map( A1 => n2912, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n2932
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n2905);
   U2058 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n2904);
   U2059 : NAND2_X1 port map( A1 => n2905, A2 => n2904, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U2060 : AOI22_X1 port map( A1 => n2912, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n2932
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n2907);
   U2061 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n2906);
   U2062 : NAND2_X1 port map( A1 => n2907, A2 => n2906, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U2063 : AOI22_X1 port map( A1 => n2912, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n2932
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n2909);
   U2064 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n2908);
   U2065 : NAND2_X1 port map( A1 => n2909, A2 => n2908, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U2066 : AOI22_X1 port map( A1 => n2912, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n2911);
   U2067 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n2910);
   U2068 : NAND2_X1 port map( A1 => n2911, A2 => n2910, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U2069 : AOI22_X1 port map( A1 => n2912, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n2914);
   U2070 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n2913);
   U2071 : NAND2_X1 port map( A1 => n2914, A2 => n2913, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U2072 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n2916);
   U2073 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n2915);
   U2074 : NAND2_X1 port map( A1 => n2916, A2 => n2915, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U2075 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n2918);
   U2076 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n2917);
   U2077 : NAND2_X1 port map( A1 => n2918, A2 => n2917, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U2078 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n2920);
   U2079 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n2919);
   U2080 : NAND2_X1 port map( A1 => n2920, A2 => n2919, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U2081 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n2932
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n2922);
   U2082 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n2921);
   U2083 : NAND2_X1 port map( A1 => n2922, A2 => n2921, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U2084 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n2925);
   U2085 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n2923
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n2924);
   U2086 : NAND2_X1 port map( A1 => n2925, A2 => n2924, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U2087 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n2927);
   U2088 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n2926);
   U2089 : NAND2_X1 port map( A1 => n2927, A2 => n2926, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U2090 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n2928
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n2931);
   U2091 : AOI22_X1 port map( A1 => n2929, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n2930);
   U2092 : NAND2_X1 port map( A1 => n2931, A2 => n2930, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U2093 : AOI22_X1 port map( A1 => n2933, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n2932
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n2937);
   U2094 : AOI22_X1 port map( A1 => n2935, A2 => 
                           boothmul_pipelined_i_muxes_in_4_50_port, B1 => n2934
                           , B2 => boothmul_pipelined_i_muxes_in_4_176_port, ZN
                           => n2936);
   U2095 : NAND2_X1 port map( A1 => n2937, A2 => n2936, ZN => 
                           boothmul_pipelined_i_mux_out_4_23_port);
   U2096 : CLKBUF_X1 port map( A => n2950, Z => n2971);
   U2097 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_205_port, B1 => 
                           n2966, B2 => 
                           boothmul_pipelined_i_muxes_in_5_205_port, ZN => 
                           n2939);
   U2098 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_68_port, B1 => n2961
                           , B2 => boothmul_pipelined_i_muxes_in_5_204_port, ZN
                           => n2938);
   U2099 : NAND2_X1 port map( A1 => n2939, A2 => n2938, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2100 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_5_68_port, A2
                           => n2950, B1 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, B2 => 
                           n2970, ZN => n2941);
   U2101 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n2961
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n2940);
   U2102 : NAND2_X1 port map( A1 => n2941, A2 => n2940, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2103 : AOI22_X1 port map( A1 => n2950, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n2970
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n2943);
   U2104 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n2961
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n2942);
   U2105 : NAND2_X1 port map( A1 => n2943, A2 => n2942, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2106 : AOI22_X1 port map( A1 => n2950, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n2970
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n2945);
   U2107 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n2961
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n2944);
   U2108 : NAND2_X1 port map( A1 => n2945, A2 => n2944, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2109 : AOI22_X1 port map( A1 => n2950, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n2970
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n2947);
   U2110 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n2946);
   U2111 : NAND2_X1 port map( A1 => n2947, A2 => n2946, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2112 : AOI22_X1 port map( A1 => n2950, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n2949);
   U2113 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n2948);
   U2114 : NAND2_X1 port map( A1 => n2949, A2 => n2948, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2115 : AOI22_X1 port map( A1 => n2950, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n2952);
   U2116 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n2961
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n2951);
   U2117 : NAND2_X1 port map( A1 => n2952, A2 => n2951, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2118 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n2954);
   U2119 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n2961
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n2953);
   U2120 : NAND2_X1 port map( A1 => n2954, A2 => n2953, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2121 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n2956);
   U2122 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n2955);
   U2123 : NAND2_X1 port map( A1 => n2956, A2 => n2955, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2124 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n2958);
   U2125 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n2957);
   U2126 : NAND2_X1 port map( A1 => n2958, A2 => n2957, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2127 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n2970
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n2960);
   U2128 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n2959);
   U2129 : NAND2_X1 port map( A1 => n2960, A2 => n2959, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2130 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n2963);
   U2131 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n2961
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n2962);
   U2132 : NAND2_X1 port map( A1 => n2963, A2 => n2962, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2133 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n2965);
   U2134 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n2964);
   U2135 : NAND2_X1 port map( A1 => n2965, A2 => n2964, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2136 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n2966
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n2969);
   U2137 : AOI22_X1 port map( A1 => n2967, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n2968);
   U2138 : NAND2_X1 port map( A1 => n2969, A2 => n2968, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2139 : AOI22_X1 port map( A1 => n2971, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n2970
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n2975);
   U2140 : AOI22_X1 port map( A1 => n2973, A2 => 
                           boothmul_pipelined_i_muxes_in_5_54_port, B1 => n2972
                           , B2 => boothmul_pipelined_i_muxes_in_5_190_port, ZN
                           => n2974);
   U2141 : NAND2_X1 port map( A1 => n2975, A2 => n2974, ZN => 
                           boothmul_pipelined_i_mux_out_5_25_port);
   U2142 : CLKBUF_X1 port map( A => n2988, Z => n3009);
   U2143 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_73_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_73_port, ZN 
                           => n2977);
   U2144 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_72_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_218_port, ZN
                           => n2976);
   U2145 : NAND2_X1 port map( A1 => n2977, A2 => n2976, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2146 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_6_72_port, A2
                           => n2988, B1 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, B2 => 
                           n3008, ZN => n2979);
   U2147 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n2978);
   U2148 : NAND2_X1 port map( A1 => n2979, A2 => n2978, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2149 : AOI22_X1 port map( A1 => n2988, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n3008
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n2981);
   U2150 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n2980);
   U2151 : NAND2_X1 port map( A1 => n2981, A2 => n2980, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2152 : AOI22_X1 port map( A1 => n2988, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n3008
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n2983);
   U2153 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n2982);
   U2154 : NAND2_X1 port map( A1 => n2983, A2 => n2982, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2155 : AOI22_X1 port map( A1 => n2988, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n3008
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n2985);
   U2156 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n2984);
   U2157 : NAND2_X1 port map( A1 => n2985, A2 => n2984, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2158 : AOI22_X1 port map( A1 => n2988, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n2987);
   U2159 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n2986);
   U2160 : NAND2_X1 port map( A1 => n2987, A2 => n2986, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2161 : AOI22_X1 port map( A1 => n2988, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n2990);
   U2162 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n2989);
   U2163 : NAND2_X1 port map( A1 => n2990, A2 => n2989, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2164 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n2992);
   U2165 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n2991);
   U2166 : NAND2_X1 port map( A1 => n2992, A2 => n2991, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2167 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n2994);
   U2168 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n2993);
   U2169 : NAND2_X1 port map( A1 => n2994, A2 => n2993, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2170 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n2996);
   U2171 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n2995);
   U2172 : NAND2_X1 port map( A1 => n2996, A2 => n2995, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2173 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n3008
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n2998);
   U2174 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n2997);
   U2175 : NAND2_X1 port map( A1 => n2998, A2 => n2997, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2176 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n3001);
   U2177 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n2999
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n3000);
   U2178 : NAND2_X1 port map( A1 => n3001, A2 => n3000, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2179 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n3003);
   U2180 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n3002);
   U2181 : NAND2_X1 port map( A1 => n3003, A2 => n3002, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2182 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n3004
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n3007);
   U2183 : AOI22_X1 port map( A1 => n3005, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n3006);
   U2184 : NAND2_X1 port map( A1 => n3007, A2 => n3006, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2185 : AOI22_X1 port map( A1 => n3009, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n3008
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n3013);
   U2186 : AOI22_X1 port map( A1 => n3011, A2 => 
                           boothmul_pipelined_i_muxes_in_6_58_port, B1 => n3010
                           , B2 => boothmul_pipelined_i_muxes_in_6_204_port, ZN
                           => n3012);
   U2187 : NAND2_X1 port map( A1 => n3013, A2 => n3012, ZN => 
                           boothmul_pipelined_i_mux_out_6_27_port);
   U2188 : CLKBUF_X1 port map( A => n3043, Z => n3049);
   U2189 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_76_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_232_port, ZN
                           => n3016);
   U2190 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_13_port, 
                           A3 => n3081, ZN => n3052);
   U2191 : CLKBUF_X1 port map( A => n3052, Z => n3040);
   U2192 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, A2 
                           => n3014, ZN => n3050);
   U2193 : CLKBUF_X1 port map( A => n3050, Z => n3046);
   U2194 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_233_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_77_port
                           , ZN => n3015);
   U2195 : NAND2_X1 port map( A1 => n3016, A2 => n3015, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2196 : AOI22_X1 port map( A1 => n3043, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_231_port, ZN
                           => n3018);
   U2197 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, B1 => 
                           n3050, B2 => boothmul_pipelined_i_muxes_in_7_76_port
                           , ZN => n3017);
   U2198 : NAND2_X1 port map( A1 => n3018, A2 => n3017, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2199 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_230_port, ZN
                           => n3020);
   U2200 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_231_port, B1 => 
                           n3050, B2 => boothmul_pipelined_i_muxes_in_7_75_port
                           , ZN => n3019);
   U2201 : NAND2_X1 port map( A1 => n3020, A2 => n3019, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2202 : AOI22_X1 port map( A1 => n3043, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_229_port, ZN
                           => n3022);
   U2203 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_230_port, B1 => 
                           n3050, B2 => boothmul_pipelined_i_muxes_in_7_74_port
                           , ZN => n3021);
   U2204 : NAND2_X1 port map( A1 => n3022, A2 => n3021, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2205 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_228_port, ZN
                           => n3024);
   U2206 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_229_port, B1 => 
                           n3050, B2 => boothmul_pipelined_i_muxes_in_7_73_port
                           , ZN => n3023);
   U2207 : NAND2_X1 port map( A1 => n3024, A2 => n3023, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2208 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => n3051
                           , B2 => boothmul_pipelined_i_muxes_in_7_227_port, ZN
                           => n3026);
   U2209 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_228_port, B1 => 
                           n3050, B2 => boothmul_pipelined_i_muxes_in_7_72_port
                           , ZN => n3025);
   U2210 : NAND2_X1 port map( A1 => n3026, A2 => n3025, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2211 : AOI22_X1 port map( A1 => n3043, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => n3051
                           , B2 => boothmul_pipelined_i_muxes_in_7_226_port, ZN
                           => n3028);
   U2212 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_227_port, B1 => 
                           n3050, B2 => boothmul_pipelined_i_muxes_in_7_71_port
                           , ZN => n3027);
   U2213 : NAND2_X1 port map( A1 => n3028, A2 => n3027, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2214 : AOI22_X1 port map( A1 => n3043, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_225_port, ZN
                           => n3030);
   U2215 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_226_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_70_port
                           , ZN => n3029);
   U2216 : NAND2_X1 port map( A1 => n3030, A2 => n3029, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2217 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_224_port, ZN
                           => n3032);
   U2218 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_225_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_69_port
                           , ZN => n3031);
   U2219 : NAND2_X1 port map( A1 => n3032, A2 => n3031, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2220 : AOI22_X1 port map( A1 => n3043, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => n3051
                           , B2 => boothmul_pipelined_i_muxes_in_7_223_port, ZN
                           => n3034);
   U2221 : AOI22_X1 port map( A1 => n3052, A2 => 
                           boothmul_pipelined_i_muxes_in_7_224_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_68_port
                           , ZN => n3033);
   U2222 : NAND2_X1 port map( A1 => n3034, A2 => n3033, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2223 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => n3051
                           , B2 => boothmul_pipelined_i_muxes_in_7_222_port, ZN
                           => n3036);
   U2224 : AOI22_X1 port map( A1 => n3052, A2 => 
                           boothmul_pipelined_i_muxes_in_7_223_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_67_port
                           , ZN => n3035);
   U2225 : NAND2_X1 port map( A1 => n3036, A2 => n3035, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2226 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => n3051
                           , B2 => boothmul_pipelined_i_muxes_in_7_221_port, ZN
                           => n3038);
   U2227 : AOI22_X1 port map( A1 => n3052, A2 => 
                           boothmul_pipelined_i_muxes_in_7_222_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_66_port
                           , ZN => n3037);
   U2228 : NAND2_X1 port map( A1 => n3038, A2 => n3037, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2229 : AOI22_X1 port map( A1 => n3043, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => n3039
                           , B2 => boothmul_pipelined_i_muxes_in_7_220_port, ZN
                           => n3042);
   U2230 : AOI22_X1 port map( A1 => n3040, A2 => 
                           boothmul_pipelined_i_muxes_in_7_221_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_65_port
                           , ZN => n3041);
   U2231 : NAND2_X1 port map( A1 => n3042, A2 => n3041, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2232 : AOI22_X1 port map( A1 => n3043, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => n3051
                           , B2 => boothmul_pipelined_i_muxes_in_7_219_port, ZN
                           => n3045);
   U2233 : AOI22_X1 port map( A1 => n3052, A2 => 
                           boothmul_pipelined_i_muxes_in_7_220_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_64_port
                           , ZN => n3044);
   U2234 : NAND2_X1 port map( A1 => n3045, A2 => n3044, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2235 : AOI22_X1 port map( A1 => n3049, A2 => 
                           boothmul_pipelined_i_muxes_in_7_62_port, B1 => n3051
                           , B2 => boothmul_pipelined_i_muxes_in_7_218_port, ZN
                           => n3048);
   U2236 : AOI22_X1 port map( A1 => n3052, A2 => 
                           boothmul_pipelined_i_muxes_in_7_219_port, B1 => 
                           n3046, B2 => boothmul_pipelined_i_muxes_in_7_63_port
                           , ZN => n3047);
   U2237 : NAND2_X1 port map( A1 => n3048, A2 => n3047, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2238 : OAI21_X1 port map( B1 => n3050, B2 => n3049, A => 
                           boothmul_pipelined_i_muxes_in_7_62_port, ZN => n3054
                           );
   U2239 : AOI22_X1 port map( A1 => n3052, A2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, B1 => 
                           n3051, B2 => 
                           boothmul_pipelined_i_muxes_in_7_217_port, ZN => 
                           n3053);
   U2240 : NAND2_X1 port map( A1 => n3054, A2 => n3053, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2241 : OAI222_X1 port map( A1 => n3075, A2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_1_port, 
                           B1 => n3070, B2 => n3055, C1 => n3069, C2 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_0_port, 
                           ZN => boothmul_pipelined_i_sum_out_1_1_port);
   U2242 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_114_port, ZN 
                           => n3057);
   U2243 : OAI222_X1 port map( A1 => n3070, A2 => n3057, B1 => n3069, B2 => 
                           n3056, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_3_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U2244 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_113_port, ZN 
                           => n3058);
   U2245 : OAI222_X1 port map( A1 => n3070, A2 => n3058, B1 => n3069, B2 => 
                           n3057, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_4_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U2246 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_112_port, ZN 
                           => n3059);
   U2247 : OAI222_X1 port map( A1 => n3070, A2 => n3059, B1 => n3069, B2 => 
                           n3058, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_5_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U2248 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_111_port, ZN 
                           => n3060);
   U2249 : OAI222_X1 port map( A1 => n3070, A2 => n3060, B1 => n3069, B2 => 
                           n3059, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_6_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U2250 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_110_port, ZN 
                           => n3061);
   U2251 : OAI222_X1 port map( A1 => n3070, A2 => n3061, B1 => n3069, B2 => 
                           n3060, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_7_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U2252 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_109_port, ZN 
                           => n3062);
   U2253 : OAI222_X1 port map( A1 => n3070, A2 => n3062, B1 => n3069, B2 => 
                           n3061, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_8_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U2254 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_108_port, ZN 
                           => n3063);
   U2255 : OAI222_X1 port map( A1 => n3070, A2 => n3063, B1 => n3069, B2 => 
                           n3062, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_9_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U2256 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_107_port, ZN 
                           => n3064);
   U2257 : OAI222_X1 port map( A1 => n3070, A2 => n3064, B1 => n3069, B2 => 
                           n3063, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_10_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U2258 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_106_port, ZN 
                           => n3065);
   U2259 : OAI222_X1 port map( A1 => n3070, A2 => n3065, B1 => n3069, B2 => 
                           n3064, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_11_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U2260 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_105_port, ZN 
                           => n3066);
   U2261 : OAI222_X1 port map( A1 => n3070, A2 => n3066, B1 => n3069, B2 => 
                           n3065, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_12_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U2262 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_104_port, ZN 
                           => n3067);
   U2263 : OAI222_X1 port map( A1 => n3070, A2 => n3067, B1 => n3069, B2 => 
                           n3066, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_13_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U2264 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_103_port, ZN 
                           => n3068);
   U2265 : OAI222_X1 port map( A1 => n3070, A2 => n3068, B1 => n3069, B2 => 
                           n3067, C1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_14_port, 
                           C2 => n3075, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U2266 : INV_X1 port map( A => n3069, ZN => n3073);
   U2267 : INV_X1 port map( A => n3070, ZN => n3072);
   U2268 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n3073, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n3072, ZN => n3071);
   U2269 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           B2 => n3075, A => n3071, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2270 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n3073, B1 => n3072, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n3074);
   U2271 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_A_15_port, 
                           B2 => n3075, A => n3074, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N385, N386, N387, N388, N389, N390, N391, N392, N393
      , N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, 
      n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, 
      n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, 
      n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, 
      n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, 
      n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, 
      n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, 
      n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, 
      n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, 
      n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, 
      n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, 
      n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, 
      n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, 
      n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, 
      n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, 
      n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
      n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, 
      n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, 
      n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, 
      n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, 
      n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, 
      n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, 
      n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
      n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, 
      n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, 
      n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, 
      n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, 
      n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, 
      n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
      n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, 
      n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, 
      n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
      n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, 
      n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, 
      n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, 
      n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, 
      n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, 
      n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, 
      n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, 
      n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
      n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, 
      n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, 
      n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, 
      n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, 
      n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, 
      n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, 
      n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, 
      n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, 
      n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, 
      n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, 
      n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, 
      n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, 
      n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, 
      n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, 
      n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, 
      n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, 
      n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, 
      n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, 
      n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, 
      n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, 
      n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, 
      n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, 
      n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, 
      n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, 
      n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, 
      n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, 
      n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, 
      n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, 
      n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, 
      n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, 
      n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, 
      n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, 
      n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, 
      n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, 
      n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, 
      n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, 
      n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, 
      n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, 
      n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, 
      n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, 
      n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, 
      n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, 
      n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, 
      n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, 
      n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, 
      n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, 
      n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, 
      n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, 
      n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, 
      n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, 
      n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, 
      n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, 
      n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, 
      n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, 
      n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, 
      n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, 
      n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, 
      n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, 
      n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, 
      n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, 
      n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, 
      n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, 
      n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, 
      n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, 
      n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, 
      n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, 
      n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, 
      n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, 
      n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, 
      n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, 
      n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, 
      n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, 
      n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, 
      n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, 
      n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, 
      n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, 
      n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, 
      n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, 
      n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, 
      n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, 
      n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, 
      n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, 
      n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, 
      n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, 
      n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, 
      n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, 
      n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, 
      n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, 
      n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, 
      n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, 
      n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, 
      n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, 
      n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, 
      n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
      n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, 
      n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, 
      n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, 
      n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
      n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, 
      n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, 
      n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, 
      n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, 
      n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, 
      n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, 
      n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, 
      n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, 
      n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, 
      n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, 
      n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
      n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
      n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, 
      n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, 
      n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, 
      n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, 
      n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, 
      n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, 
      n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, 
      n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, 
      n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, 
      n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, 
      n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, 
      n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
      n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, 
      n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, 
      n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, 
      n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, 
      n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, 
      n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, 
      n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, 
      n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, 
      n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, 
      n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, 
      n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, 
      n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, 
      n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, 
      n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, 
      n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, 
      n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, 
      n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, 
      n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, 
      n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, 
      n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, 
      n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, 
      n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, 
      n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, 
      n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, 
      n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, 
      n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, 
      n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, 
      n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, 
      n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, 
      n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, 
      n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, 
      n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, 
      n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, 
      n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, 
      n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, 
      n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, 
      n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, 
      n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, 
      n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, 
      n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, 
      n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, 
      n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, 
      n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, 
      n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, 
      n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, 
      n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, 
      n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, 
      n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, 
      n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, 
      n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, 
      n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, 
      n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, 
      n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, 
      n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, 
      n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, 
      n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, 
      n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, 
      n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, 
      n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, 
      n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, 
      n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, 
      n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, 
      n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, 
      n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, 
      n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, 
      n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, 
      n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, 
      n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, 
      n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, 
      n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, 
      n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, 
      n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, 
      n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, 
      n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, 
      n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, 
      n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, 
      n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, 
      n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, 
      n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, 
      n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, 
      n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, 
      n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, 
      n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, 
      n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, 
      n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, 
      n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, 
      n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, 
      n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, 
      n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, 
      n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, 
      n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, 
      n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, 
      n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, 
      n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, 
      n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, 
      n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, 
      n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, 
      n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, 
      n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, 
      n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, 
      n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, 
      n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, 
      n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, 
      n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, 
      n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, 
      n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, 
      n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, 
      n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, 
      n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, 
      n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, 
      n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, 
      n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, 
      n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, 
      n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, 
      n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, 
      n5665, n5666, n5667, n5668, n5669, n5670, n5671, n_1357, n_1358, n_1359, 
      n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, 
      n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, 
      n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, 
      n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, 
      n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, 
      n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, 
      n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n5168);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n5169);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n5408);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n5170);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n5409);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n5410);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n5171);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n5172);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n5173);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n5174);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n5411);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n5412);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n5413);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n5414);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n5175);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n5415);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n5176);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n5177);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n5416);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n5178);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n5417);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n5179);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n5180);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n5418);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n5419);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n5420);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n5181);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n5182);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n5421);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n5183);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n5422);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n5184);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n4924);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n5423);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n5185);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           REGISTERS_1_28_port, QN => n4652);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n4925);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n5424);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n5425);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n4926);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n5426);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n4927);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n5186);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n5427);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n5187);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n5428);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n5188);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n5429);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n4928);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n5430);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n5189);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n4929);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n4930);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n4653);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n5431);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n4654);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n4655);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n5190);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n5432);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n4656);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n5191);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n4657);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n5192);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n4658);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n4659);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n5433);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n4931);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n5193);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n5434);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n4660);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n4932);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n4661);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n4933);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n5194);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n4934);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n4662);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n4663);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n4664);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n4935);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n4665);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n4936);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n4937);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n4666);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n4938);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n5195);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n4939);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n4940);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n4667);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n4941);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n4942);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n5435);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n5436);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n4943);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n5437);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n4668);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n5438);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n5439);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n4669);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n4944);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n4945);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n4670);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n4946);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n4947);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n5440);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n4671);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n4948);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n4672);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n4673);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n4674);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n4675);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n4676);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n4949);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n5196);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n5441);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n4677);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n4678);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n4950);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n5197);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n4679);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n4680);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n5442);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n4681);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n4951);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n4682);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n4952);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n4953);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n4683);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n4684);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n5443);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n4685);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n5198);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n5444);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n5199);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n5200);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n5201);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n5445);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n5202);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n5446);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n4686);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n5203);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n5447);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n5204);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n5448);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n5205);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n5449);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n5206);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n5207);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n5450);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n4687);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n5451);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n5208);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n5209);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n5210);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n5211);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n4688);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n5452);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n5453);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n4954);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n4689);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n5212);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n4690);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n5454);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n4691);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n4955);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n5213);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n5214);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n4692);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n5215);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n5455);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n5216);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n5217);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n5218);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n5456);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n4956);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n5219);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           REGISTERS_5_16_port, QN => n5220);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n4957);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n4693);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n5457);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n5458);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n5221);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n5459);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n5222);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n5460);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n5461);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n4958);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n5223);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n5224);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n5225);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n5226);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n5462);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n5463);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n5227);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n4959);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n5464);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n5465);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n4694);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n4695);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n5466);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n4696);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n4697);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n4960);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n5467);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n4961);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n4698);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n5468);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n4962);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n4699);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n5228);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n4963);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n4964);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n5229);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n5469);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n4965);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n4966);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n5470);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n4700);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n5471);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n4701);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n4967);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n4702);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n5230);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n5472);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n4968);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n4969);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n4703);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n4704);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n4705);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n4970);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n4971);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n4706);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n4972);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n4973);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n4707);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n4974);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n4975);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n4976);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n4708);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n4977);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n4978);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n4709);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n4710);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n4979);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n4711);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n4712);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n4713);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n4980);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n4981);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n4714);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n4715);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n4982);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n4983);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n4716);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n4984);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n4985);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n4986);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n5473);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n5474);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n5231);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n5232);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n5475);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n5233);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n5476);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n5234);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n5235);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n5236);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n5477);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n5478);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n5237);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n5238);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n5239);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n5240);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n5479);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n5480);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n5481);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n5482);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n5241);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n5242);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n5243);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n5244);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n5483);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n5245);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n5484);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n5246);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n5485);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n5247);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n5248);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n5486);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n4717);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n5487);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n4718);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n4987);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n4988);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n4719);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n4720);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n4989);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n4990);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n5249);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n5488);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n5489);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n4721);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n5490);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n5250);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n4722);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n4991);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n4723);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n5251);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n4992);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n4724);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n5491);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n5492);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n5493);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n5494);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n5495);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n5252);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n5496);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n5253);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n5497);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n4725);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n4726);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n4727);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n4993);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n4728);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n4729);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n5254);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n4730);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n4731);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n4994);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n5255);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n4732);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n4995);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n4733);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n4734);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n4735);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n4996);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n4997);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n4736);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n4998);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           REGISTERS_10_13_port, QN => n4737);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n4738);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n4999);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n5000);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n5001);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           REGISTERS_10_8_port, QN => n4739);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n4740);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n4741);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n4742);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n4743);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n4744);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n5002);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n5498);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n4745);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n5256);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n4746);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n5003);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n5004);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n5005);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n5499);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n5006);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n5007);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n5008);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n5500);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n4747);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n5009);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n5501);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n4748);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n5010);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n5502);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n4749);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n5257);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n4750);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n5011);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n5258);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n4751);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n4752);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n4753);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n5012);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n5013);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n4754);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n5014);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n5015);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n4755);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n4756);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n5503);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n5504);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n4757);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n5505);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n5259);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n5260);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n5506);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n5261);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n5507);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n5262);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n5016);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n5263);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n4758);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n5017);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n4759);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n5018);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n5508);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n5264);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n4760);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n5265);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           REGISTERS_12_12_port, QN => n5266);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n5267);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n5019);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n4761);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n4762);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n5509);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n5268);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n5020);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n5510);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n5511);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n4763);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n5512);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n5513);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n5514);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n5269);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n5270);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n5515);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n5271);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n5516);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n5272);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n5273);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n5517);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n5518);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n5274);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n5275);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n5276);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n5519);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n5520);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n5277);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n5521);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n5522);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n5523);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n5278);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n5524);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n5279);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n5525);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n5526);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n5280);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n5527);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n5528);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n5281);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n5021);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n5282);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n5529);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n5022);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n4764);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n5530);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n5531);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n5283);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n5023);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n4765);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n5532);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n5284);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n5024);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n4766);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n5025);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n5285);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n5533);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n5534);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n5286);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n5026);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n5287);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n5535);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n5027);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n5536);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n5028);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n5537);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n5288);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n5538);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n4767);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n4768);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n5289);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n4769);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n5290);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n5539);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n4770);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n5291);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n5029);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n4771);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n5030);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n5031);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n4772);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n5032);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n5033);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n4773);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n4774);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n5034);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n4775);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n5035);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n5036);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n5037);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n4776);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n4777);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n5038);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n4778);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n5039);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n4779);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n5040);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n4780);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n5041);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n5042);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n4781);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n5043);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n5044);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n5045);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n4782);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n5046);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n5047);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n4783);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n5164);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n5292);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n5293);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n5540);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n5294);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n5295);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n5296);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n5541);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n4784);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n5542);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n5297);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n5298);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n4785);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n5543);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n5299);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n5544);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n5545);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n5300);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n5546);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n5301);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n5547);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n4786);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n5548);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n5549);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n5550);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n5302);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n5303);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n5551);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n5304);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n5552);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n4787);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n5048);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n4916);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n5553);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n5305);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n5049);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n4788);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           REGISTERS_17_26_port, QN => n5554);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n5555);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n5306);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n5556);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n4789);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n4790);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n4791);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n5050);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n5051);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n5307);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n5557);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n5308);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n5558);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n4792);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n5309);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n5310);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n5052);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n5311);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n4793);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n5559);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n5560);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n5312);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n5561);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n4794);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n5562);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n4795);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n4796);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n4917);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n5053);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n5054);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n5055);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n5056);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n4797);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n5057);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n5058);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n5059);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n4798);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n4799);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n5060);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n4800);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n4801);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n5061);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n5062);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n5063);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n5313);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n5064);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n4802);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n5065);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n4803);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n5066);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n4804);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n4805);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n5067);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n5068);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n4806);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n5069);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n4807);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           REGISTERS_18_1_port, QN => n5070);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n5071);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n4918);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n4808);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n5563);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n4809);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n4810);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n5564);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n5072);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n4811);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n5073);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n5074);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n5075);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n5565);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n5076);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n5566);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n5314);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n5567);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n5077);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n5078);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n4812);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n5079);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n5080);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n5568);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n4813);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n4814);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n4815);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n4816);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n5315);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n4817);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n5316);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n4818);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n5569);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n5570);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n4919);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n4819);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n4820);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n5571);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n5317);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n4821);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n4822);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n5081);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n5572);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n5573);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n4823);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n5082);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n4824);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n5318);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           REGISTERS_20_17_port, QN => n5083);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n4825);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n5574);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n5084);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n4826);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n4827);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n4828);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n5319);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n5320);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n5085);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n5575);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n4829);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n5576);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n4830);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n5577);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n4831);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n4832);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n5321);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n5165);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n5322);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n5323);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n5324);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n5578);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n5325);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n5579);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n5580);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n5581);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n5086);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n5582);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n4833);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n5583);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n4834);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n5584);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n5326);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n5087);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n4835);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n5585);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n5088);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n5586);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n4836);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n5587);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n5588);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n5089);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n5327);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n5589);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n5590);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n5328);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n5090);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n5591);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n5329);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n5166);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n5330);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n5592);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n5331);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n5593);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n5332);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n5333);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n5594);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n5091);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n5334);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n5092);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n5595);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n5596);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n4837);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n5597);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n5093);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n5335);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n5598);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n5336);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n5094);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n5599);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n5337);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n5600);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n5338);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n5601);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n5602);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n4838);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n5603);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n5095);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n5339);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n5340);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n5341);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n4648);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n5096);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n5097);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n5098);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n5099);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n4839);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n4840);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n4841);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n4842);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n4843);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n5100);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n4844);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n5101);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           REGISTERS_23_18_port, QN => n5102);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n5103);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n4845);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n4846);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n4847);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n5604);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n4848);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n4849);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n4850);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n5104);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n5105);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n5106);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n5342);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n5107);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n4851);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n5108);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n5605);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n4852);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n4853);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n5167);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n5606);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n5343);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n5607);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n5608);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n5609);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n5344);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n5345);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n5346);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n5610);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n5611);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n5347);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n5348);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n5349);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n5350);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n5351);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n5352);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n5353);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n5612);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n5613);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n5354);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n5614);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n5355);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n5615);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n5356);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n5616);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n5357);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n5358);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n5617);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n5359);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n5360);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n5361);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n4920);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n5109);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n4854);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n4855);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n5110);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n4856);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n4857);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n4858);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n4859);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n5111);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n5362);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n4860);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n5363);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n5364);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n4861);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n4862);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n4863);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n4864);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n5112);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n5113);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n5114);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n4865);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n4866);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n5365);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n4867);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n5115);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n5116);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n4868);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n4869);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n5117);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n5618);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n4870);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n4921);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n5619);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n4871);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n4872);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n4873);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n5366);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n5118);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n4874);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n5367);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n5368);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n5369);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n4875);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n5119);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n5620);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n5120);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n5121);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n5122);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n4876);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n4877);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n5370);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n5621);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n5123);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n5622);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n5124);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n5623);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n5624);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n4878);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n5625);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n5125);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n5626);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n5126);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n5627);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n4649);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n5127);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n5128);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n5129);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n5130);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n5131);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n4879);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n5132);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n4880);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n4881);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n5133);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n5134);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n4882);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n5135);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n4883);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n4884);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n5136);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n4885);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           REGISTERS_27_13_port, QN => n4886);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n4887);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n4888);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n5137);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n4889);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n5138);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n4890);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n4891);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n5139);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n4892);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n4893);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n5140);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n4894);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n5141);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n4922);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n5371);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n5628);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n5372);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n5373);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n5629);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n5630);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n5374);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n5631);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n5375);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n5632);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n5633);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n5634);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n5635);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n4895);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n5636);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n5376);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n5637);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n5377);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n5638);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n5378);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n5639);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n5142);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n5640);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n5641);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n4896);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n5379);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n5642);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n5643);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n5380);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n5644);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n5645);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n4923);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n5646);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n5143);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n5381);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n5382);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n5144);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n5383);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n5647);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           REGISTERS_29_23_port, QN => n5648);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n5649);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n5650);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n5651);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n5384);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n5385);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n5652);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n5653);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n5386);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n5654);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n5387);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n5655);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n5388);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n5656);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n5389);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n5390);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n5391);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n5145);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n5392);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n5393);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n5657);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n5394);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n5658);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n5395);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n4650);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n4897);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n4898);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n5659);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n4899);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n5146);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n5660);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n5147);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n5396);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n4900);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n4901);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           REGISTERS_30_20_port, QN => n5397);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n5661);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n5148);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n4902);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n5398);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n4903);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n5662);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n5663);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n5399);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n5149);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n5400);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n4904);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n4905);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n4906);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n5401);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n5150);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n5151);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n4907);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n4908);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n5152);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n5153);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n4651);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n4909);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n5664);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n4910);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n5665);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n5154);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n5155);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n5402);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n4911);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n5666);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n5403);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n5667);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n5404);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n4912);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n5668);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n4913);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n5669);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n5156);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n5157);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n5670);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n4914);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n5671);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n5158);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n5405);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n4915);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n5159);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n5160);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n5161);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n5406);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n5162);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n5407);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n5163);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT1(31), QN 
                           => n_1357);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT1(30), QN 
                           => n_1358);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT1(29), QN 
                           => n_1359);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT1(28), QN 
                           => n_1360);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT1(27), QN 
                           => n_1361);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT1(26), QN 
                           => n_1362);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT1(25), QN 
                           => n_1363);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT1(24), QN 
                           => n_1364);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT1(23), QN 
                           => n_1365);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => CLK, Q => OUT1(22), QN 
                           => n_1366);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => CLK, Q => OUT1(21), QN 
                           => n_1367);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => CLK, Q => OUT1(20), QN 
                           => n_1368);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => CLK, Q => OUT1(19), QN 
                           => n_1369);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => CLK, Q => OUT1(18), QN 
                           => n_1370);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => CLK, Q => OUT1(17), QN 
                           => n_1371);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => CLK, Q => OUT1(16), QN 
                           => n_1372);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => CLK, Q => OUT1(15), QN 
                           => n_1373);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => CLK, Q => OUT1(14), QN 
                           => n_1374);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => CLK, Q => OUT1(13), QN 
                           => n_1375);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => CLK, Q => OUT1(12), QN 
                           => n_1376);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => CLK, Q => OUT1(11), QN 
                           => n_1377);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => CLK, Q => OUT1(10), QN 
                           => n_1378);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => CLK, Q => OUT1(9), QN =>
                           n_1379);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => CLK, Q => OUT1(8), QN =>
                           n_1380);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => CLK, Q => OUT1(7), QN =>
                           n_1381);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => CLK, Q => OUT1(6), QN =>
                           n_1382);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => CLK, Q => OUT1(5), QN =>
                           n_1383);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => CLK, Q => OUT1(4), QN =>
                           n_1384);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => CLK, Q => OUT1(3), QN =>
                           n_1385);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => CLK, Q => OUT1(2), QN =>
                           n_1386);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => CLK, Q => OUT1(1), QN =>
                           n_1387);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT2(31), QN 
                           => n_1388);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT2(30), QN 
                           => n_1389);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT2(29), QN 
                           => n_1390);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT2(28), QN 
                           => n_1391);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT2(27), QN 
                           => n_1392);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT2(26), QN 
                           => n_1393);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT2(25), QN 
                           => n_1394);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT2(24), QN 
                           => n_1395);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT2(23), QN 
                           => n_1396);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(22), QN 
                           => n_1397);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(21), QN 
                           => n_1398);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(20), QN 
                           => n_1399);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(19), QN 
                           => n_1400);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(18), QN 
                           => n_1401);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(17), QN 
                           => n_1402);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(16), QN 
                           => n_1403);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(15), QN 
                           => n_1404);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(14), QN 
                           => n_1405);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(13), QN 
                           => n_1406);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(12), QN 
                           => n_1407);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(11), QN 
                           => n_1408);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(10), QN 
                           => n_1409);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(9), QN =>
                           n_1410);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(8), QN =>
                           n_1411);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(7), QN =>
                           n_1412);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(6), QN =>
                           n_1413);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(5), QN =>
                           n_1414);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(4), QN =>
                           n_1415);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(3), QN =>
                           n_1416);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(2), QN =>
                           n_1417);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(1), QN =>
                           n_1418);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(0), QN =>
                           n_1419);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => CLK, Q => OUT1(0), QN =>
                           n_1420);
   U3 : CLKBUF_X1 port map( A => RESET_BAR, Z => n2895);
   U4 : CLKBUF_X1 port map( A => RESET_BAR, Z => n2896);
   U5 : CLKBUF_X1 port map( A => RESET_BAR, Z => n2897);
   U6 : CLKBUF_X1 port map( A => RESET_BAR, Z => n2898);
   U7 : NAND2_X2 port map( A1 => n2895, A2 => n3072, ZN => n3084);
   U8 : NAND2_X2 port map( A1 => n2898, A2 => n3045, ZN => n3047);
   U9 : NAND2_X2 port map( A1 => n2895, A2 => n3041, ZN => n3043);
   U10 : NAND2_X2 port map( A1 => n2896, A2 => n3037, ZN => n3039);
   U11 : NAND2_X2 port map( A1 => n2895, A2 => n3033, ZN => n3035);
   U12 : NAND2_X2 port map( A1 => n2896, A2 => n3029, ZN => n3031);
   U13 : NAND2_X2 port map( A1 => n2898, A2 => n3025, ZN => n3027);
   U14 : NAND2_X2 port map( A1 => n2898, A2 => n3021, ZN => n3023);
   U15 : NAND2_X2 port map( A1 => n2898, A2 => n3015, ZN => n3017);
   U16 : NAND2_X2 port map( A1 => n2898, A2 => n3006, ZN => n3008);
   U17 : NAND2_X2 port map( A1 => n2895, A2 => n3003, ZN => n3005);
   U18 : NAND2_X2 port map( A1 => n2897, A2 => n3000, ZN => n3002);
   U19 : NAND2_X2 port map( A1 => n2895, A2 => n2962, ZN => n2964);
   U20 : NAND2_X2 port map( A1 => n2895, A2 => n2959, ZN => n2961);
   U21 : NAND2_X2 port map( A1 => n2895, A2 => n2956, ZN => n2958);
   U22 : NAND2_X2 port map( A1 => n2895, A2 => n2952, ZN => n2954);
   U23 : NAND2_X2 port map( A1 => n2898, A2 => n2949, ZN => n2951);
   U24 : NAND2_X2 port map( A1 => n2898, A2 => n2946, ZN => n2948);
   U25 : NAND2_X2 port map( A1 => n2895, A2 => n2939, ZN => n2941);
   U26 : NAND2_X2 port map( A1 => n2898, A2 => n2936, ZN => n2938);
   U27 : NAND2_X2 port map( A1 => n2895, A2 => n2933, ZN => n2935);
   U28 : NAND2_X2 port map( A1 => n2895, A2 => n2922, ZN => n2924);
   U29 : NAND2_X2 port map( A1 => n2898, A2 => n2918, ZN => n2920);
   U30 : NAND2_X2 port map( A1 => n2896, A2 => n2914, ZN => n2916);
   U31 : INV_X1 port map( A => ADD_WR(3), ZN => n3019);
   U32 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n2917, A3 => n2926, ZN => 
                           n3040);
   U33 : NOR2_X1 port map( A1 => ADD_WR(3), A2 => n2932, ZN => n2927);
   U34 : CLKBUF_X1 port map( A => n3866, Z => n3814);
   U35 : CLKBUF_X1 port map( A => n4647, Z => n4593);
   U36 : CLKBUF_X1 port map( A => n3029, Z => n3030);
   U37 : NAND2_X1 port map( A1 => n2896, A2 => n3009, ZN => n3012);
   U38 : NAND2_X1 port map( A1 => n2897, A2 => n2986, ZN => n2999);
   U39 : CLKBUF_X1 port map( A => n2995, Z => n3080);
   U40 : CLKBUF_X1 port map( A => n2978, Z => n3064);
   U41 : NAND2_X1 port map( A1 => n2897, A2 => n2942, ZN => n2945);
   U42 : NAND2_X1 port map( A1 => n2897, A2 => n2928, ZN => n2931);
   U43 : CLKBUF_X1 port map( A => n2914, Z => n2915);
   U44 : NAND2_X1 port map( A1 => n2896, A2 => n2904, ZN => n2907);
   U45 : CLKBUF_X1 port map( A => n2901, Z => n2902);
   U46 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1), 
                           ZN => n3020);
   U47 : INV_X1 port map( A => ADD_WR(4), ZN => n2899);
   U48 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n2899, ZN => n2932);
   U49 : NAND2_X1 port map( A1 => n3020, A2 => n2927, ZN => n2901);
   U50 : NAND2_X1 port map( A1 => n2897, A2 => n2902, ZN => n2903);
   U51 : CLKBUF_X1 port map( A => n2903, Z => n2900);
   U52 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(31), ZN => n3050);
   U53 : CLKBUF_X1 port map( A => n3050, Z => n3014);
   U54 : OAI22_X1 port map( A1 => n5168, A2 => n2900, B1 => n3014, B2 => n2902,
                           ZN => n2166);
   U55 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(30), ZN => n2965);
   U56 : OAI22_X1 port map( A1 => n5169, A2 => n2903, B1 => n2902, B2 => n2965,
                           ZN => n2165);
   U57 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(29), ZN => n2966);
   U58 : OAI22_X1 port map( A1 => n5408, A2 => n2900, B1 => n2902, B2 => n2966,
                           ZN => n2164);
   U59 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(28), ZN => n2967);
   U60 : OAI22_X1 port map( A1 => n5170, A2 => n2903, B1 => n2902, B2 => n2967,
                           ZN => n2163);
   U61 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(27), ZN => n2968);
   U62 : OAI22_X1 port map( A1 => n5409, A2 => n2900, B1 => n2902, B2 => n2968,
                           ZN => n2162);
   U63 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(26), ZN => n2969);
   U64 : OAI22_X1 port map( A1 => n5410, A2 => n2903, B1 => n2902, B2 => n2969,
                           ZN => n2161);
   U65 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(25), ZN => n2970);
   U66 : OAI22_X1 port map( A1 => n5171, A2 => n2900, B1 => n2902, B2 => n2970,
                           ZN => n2160);
   U67 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(24), ZN => n2971);
   U68 : OAI22_X1 port map( A1 => n5172, A2 => n2903, B1 => n2902, B2 => n2971,
                           ZN => n2159);
   U69 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(23), ZN => n2972);
   U70 : OAI22_X1 port map( A1 => n5173, A2 => n2900, B1 => n2901, B2 => n2972,
                           ZN => n2158);
   U71 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(22), ZN => n2973);
   U72 : OAI22_X1 port map( A1 => n5174, A2 => n2903, B1 => n2901, B2 => n2973,
                           ZN => n2157);
   U73 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(21), ZN => n2974);
   U74 : OAI22_X1 port map( A1 => n5411, A2 => n2903, B1 => n2901, B2 => n2974,
                           ZN => n2156);
   U75 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(20), ZN => n2975);
   U76 : OAI22_X1 port map( A1 => n5412, A2 => n2903, B1 => n2901, B2 => n2975,
                           ZN => n2155);
   U77 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(19), ZN => n2976);
   U78 : OAI22_X1 port map( A1 => n5413, A2 => n2900, B1 => n2901, B2 => n2976,
                           ZN => n2154);
   U79 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(18), ZN => n2977);
   U80 : OAI22_X1 port map( A1 => n5414, A2 => n2900, B1 => n2901, B2 => n2977,
                           ZN => n2153);
   U81 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(17), ZN => n2978);
   U82 : OAI22_X1 port map( A1 => n5175, A2 => n2900, B1 => n2901, B2 => n2978,
                           ZN => n2152);
   U83 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(16), ZN => n2979);
   U84 : OAI22_X1 port map( A1 => n5415, A2 => n2900, B1 => n2901, B2 => n2979,
                           ZN => n2151);
   U85 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(15), ZN => n2980);
   U86 : OAI22_X1 port map( A1 => n5176, A2 => n2900, B1 => n2902, B2 => n2980,
                           ZN => n2150);
   U87 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(14), ZN => n2981);
   U88 : OAI22_X1 port map( A1 => n5177, A2 => n2900, B1 => n2901, B2 => n2981,
                           ZN => n2149);
   U89 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(13), ZN => n2982);
   U90 : OAI22_X1 port map( A1 => n5416, A2 => n2900, B1 => n2902, B2 => n2982,
                           ZN => n2148);
   U91 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(12), ZN => n2983);
   U92 : OAI22_X1 port map( A1 => n5178, A2 => n2900, B1 => n2901, B2 => n2983,
                           ZN => n2147);
   U93 : NAND2_X1 port map( A1 => n2898, A2 => DATAIN(11), ZN => n2984);
   U94 : OAI22_X1 port map( A1 => n5417, A2 => n2900, B1 => n2901, B2 => n2984,
                           ZN => n2146);
   U95 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(10), ZN => n2985);
   U96 : OAI22_X1 port map( A1 => n5179, A2 => n2900, B1 => n2901, B2 => n2985,
                           ZN => n2145);
   U97 : NAND2_X1 port map( A1 => n2898, A2 => DATAIN(9), ZN => n2987);
   U98 : OAI22_X1 port map( A1 => n5180, A2 => n2900, B1 => n2902, B2 => n2987,
                           ZN => n2144);
   U99 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(8), ZN => n2988);
   U100 : OAI22_X1 port map( A1 => n5418, A2 => n2900, B1 => n2901, B2 => n2988
                           , ZN => n2143);
   U101 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(7), ZN => n2990);
   U102 : OAI22_X1 port map( A1 => n5419, A2 => n2903, B1 => n2902, B2 => n2990
                           , ZN => n2142);
   U103 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(6), ZN => n2991);
   U104 : OAI22_X1 port map( A1 => n5420, A2 => n2903, B1 => n2901, B2 => n2991
                           , ZN => n2141);
   U105 : NAND2_X1 port map( A1 => n2898, A2 => DATAIN(5), ZN => n2992);
   U106 : OAI22_X1 port map( A1 => n5181, A2 => n2903, B1 => n2902, B2 => n2992
                           , ZN => n2140);
   U107 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(4), ZN => n2993);
   U108 : OAI22_X1 port map( A1 => n5182, A2 => n2903, B1 => n2901, B2 => n2993
                           , ZN => n2139);
   U109 : NAND2_X1 port map( A1 => n2897, A2 => DATAIN(3), ZN => n2994);
   U110 : OAI22_X1 port map( A1 => n5421, A2 => n2903, B1 => n2902, B2 => n2994
                           , ZN => n2138);
   U111 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(2), ZN => n2995);
   U112 : OAI22_X1 port map( A1 => n5183, A2 => n2903, B1 => n2901, B2 => n2995
                           , ZN => n2137);
   U113 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(1), ZN => n2996);
   U114 : OAI22_X1 port map( A1 => n5422, A2 => n2903, B1 => n2902, B2 => n2996
                           , ZN => n2136);
   U115 : NAND2_X1 port map( A1 => n2896, A2 => DATAIN(0), ZN => n2998);
   U116 : OAI22_X1 port map( A1 => n5184, A2 => n2903, B1 => n2902, B2 => n2998
                           , ZN => n2135);
   U117 : INV_X1 port map( A => ADD_WR(0), ZN => n2917);
   U118 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n2917, ZN 
                           => n3024);
   U119 : NAND2_X1 port map( A1 => n2927, A2 => n3024, ZN => n2904);
   U120 : CLKBUF_X1 port map( A => n2907, Z => n2905);
   U121 : CLKBUF_X1 port map( A => n2904, Z => n2906);
   U122 : OAI22_X1 port map( A1 => n4924, A2 => n2905, B1 => n3050, B2 => n2906
                           , ZN => n2134);
   U123 : OAI22_X1 port map( A1 => n5423, A2 => n2907, B1 => n2965, B2 => n2904
                           , ZN => n2133);
   U124 : OAI22_X1 port map( A1 => n5185, A2 => n2905, B1 => n2966, B2 => n2906
                           , ZN => n2132);
   U125 : OAI22_X1 port map( A1 => n4652, A2 => n2907, B1 => n2967, B2 => n2904
                           , ZN => n2131);
   U126 : OAI22_X1 port map( A1 => n4925, A2 => n2905, B1 => n2968, B2 => n2906
                           , ZN => n2130);
   U127 : OAI22_X1 port map( A1 => n5424, A2 => n2907, B1 => n2969, B2 => n2904
                           , ZN => n2129);
   U128 : OAI22_X1 port map( A1 => n5425, A2 => n2905, B1 => n2970, B2 => n2906
                           , ZN => n2128);
   U129 : OAI22_X1 port map( A1 => n4926, A2 => n2907, B1 => n2971, B2 => n2904
                           , ZN => n2127);
   U130 : OAI22_X1 port map( A1 => n5426, A2 => n2905, B1 => n2972, B2 => n2906
                           , ZN => n2126);
   U131 : OAI22_X1 port map( A1 => n4927, A2 => n2907, B1 => n2973, B2 => n2904
                           , ZN => n2125);
   U132 : OAI22_X1 port map( A1 => n5186, A2 => n2907, B1 => n2974, B2 => n2904
                           , ZN => n2124);
   U133 : OAI22_X1 port map( A1 => n5427, A2 => n2907, B1 => n2975, B2 => n2906
                           , ZN => n2123);
   U134 : OAI22_X1 port map( A1 => n5187, A2 => n2905, B1 => n2976, B2 => n2904
                           , ZN => n2122);
   U135 : OAI22_X1 port map( A1 => n5428, A2 => n2905, B1 => n2977, B2 => n2906
                           , ZN => n2121);
   U136 : OAI22_X1 port map( A1 => n5188, A2 => n2905, B1 => n2978, B2 => n2904
                           , ZN => n2120);
   U137 : OAI22_X1 port map( A1 => n5429, A2 => n2905, B1 => n2979, B2 => n2906
                           , ZN => n2119);
   U138 : OAI22_X1 port map( A1 => n4928, A2 => n2905, B1 => n2980, B2 => n2904
                           , ZN => n2118);
   U139 : OAI22_X1 port map( A1 => n5430, A2 => n2905, B1 => n2981, B2 => n2904
                           , ZN => n2117);
   U140 : OAI22_X1 port map( A1 => n5189, A2 => n2905, B1 => n2982, B2 => n2904
                           , ZN => n2116);
   U141 : OAI22_X1 port map( A1 => n4929, A2 => n2905, B1 => n2983, B2 => n2904
                           , ZN => n2115);
   U142 : OAI22_X1 port map( A1 => n4930, A2 => n2905, B1 => n2984, B2 => n2904
                           , ZN => n2114);
   U143 : OAI22_X1 port map( A1 => n4653, A2 => n2905, B1 => n2985, B2 => n2904
                           , ZN => n2113);
   U144 : OAI22_X1 port map( A1 => n5431, A2 => n2905, B1 => n2987, B2 => n2904
                           , ZN => n2112);
   U145 : OAI22_X1 port map( A1 => n4654, A2 => n2905, B1 => n2988, B2 => n2906
                           , ZN => n2111);
   U146 : OAI22_X1 port map( A1 => n4655, A2 => n2907, B1 => n2990, B2 => n2906
                           , ZN => n2110);
   U147 : OAI22_X1 port map( A1 => n5190, A2 => n2907, B1 => n2991, B2 => n2906
                           , ZN => n2109);
   U148 : OAI22_X1 port map( A1 => n5432, A2 => n2907, B1 => n2992, B2 => n2906
                           , ZN => n2108);
   U149 : OAI22_X1 port map( A1 => n4656, A2 => n2907, B1 => n2993, B2 => n2906
                           , ZN => n2107);
   U150 : OAI22_X1 port map( A1 => n5191, A2 => n2907, B1 => n2994, B2 => n2906
                           , ZN => n2106);
   U151 : OAI22_X1 port map( A1 => n4657, A2 => n2907, B1 => n2995, B2 => n2906
                           , ZN => n2105);
   U152 : OAI22_X1 port map( A1 => n5192, A2 => n2907, B1 => n2996, B2 => n2906
                           , ZN => n2104);
   U153 : OAI22_X1 port map( A1 => n4658, A2 => n2907, B1 => n2998, B2 => n2906
                           , ZN => n2103);
   U154 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n2917, ZN => n2921);
   U155 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n2921, ZN => n3028);
   U156 : NAND2_X1 port map( A1 => n2927, A2 => n3028, ZN => n2908);
   U157 : NAND2_X2 port map( A1 => n2895, A2 => n2908, ZN => n2910);
   U158 : CLKBUF_X1 port map( A => n2908, Z => n2909);
   U159 : OAI22_X1 port map( A1 => n4659, A2 => n2910, B1 => n3014, B2 => n2909
                           , ZN => n2102);
   U160 : OAI22_X1 port map( A1 => n5433, A2 => n2910, B1 => n2965, B2 => n2908
                           , ZN => n2101);
   U161 : OAI22_X1 port map( A1 => n4931, A2 => n2910, B1 => n2966, B2 => n2909
                           , ZN => n2100);
   U162 : OAI22_X1 port map( A1 => n5193, A2 => n2910, B1 => n2967, B2 => n2908
                           , ZN => n2099);
   U163 : OAI22_X1 port map( A1 => n5434, A2 => n2910, B1 => n2968, B2 => n2909
                           , ZN => n2098);
   U164 : OAI22_X1 port map( A1 => n4660, A2 => n2910, B1 => n2969, B2 => n2908
                           , ZN => n2097);
   U165 : OAI22_X1 port map( A1 => n4932, A2 => n2910, B1 => n2970, B2 => n2909
                           , ZN => n2096);
   U166 : OAI22_X1 port map( A1 => n4661, A2 => n2910, B1 => n2971, B2 => n2908
                           , ZN => n2095);
   U167 : OAI22_X1 port map( A1 => n4933, A2 => n2910, B1 => n2972, B2 => n2909
                           , ZN => n2094);
   U168 : OAI22_X1 port map( A1 => n5194, A2 => n2910, B1 => n2973, B2 => n2908
                           , ZN => n2093);
   U169 : OAI22_X1 port map( A1 => n4934, A2 => n2910, B1 => n2974, B2 => n2908
                           , ZN => n2092);
   U170 : OAI22_X1 port map( A1 => n4662, A2 => n2910, B1 => n2975, B2 => n2909
                           , ZN => n2091);
   U171 : OAI22_X1 port map( A1 => n4663, A2 => n2910, B1 => n2976, B2 => n2908
                           , ZN => n2090);
   U172 : OAI22_X1 port map( A1 => n4664, A2 => n2910, B1 => n2977, B2 => n2909
                           , ZN => n2089);
   U173 : OAI22_X1 port map( A1 => n4935, A2 => n2910, B1 => n2978, B2 => n2908
                           , ZN => n2088);
   U174 : OAI22_X1 port map( A1 => n4665, A2 => n2910, B1 => n2979, B2 => n2909
                           , ZN => n2087);
   U175 : OAI22_X1 port map( A1 => n4936, A2 => n2910, B1 => n2980, B2 => n2908
                           , ZN => n2086);
   U176 : OAI22_X1 port map( A1 => n4937, A2 => n2910, B1 => n2981, B2 => n2908
                           , ZN => n2085);
   U177 : OAI22_X1 port map( A1 => n4666, A2 => n2910, B1 => n2982, B2 => n2908
                           , ZN => n2084);
   U178 : OAI22_X1 port map( A1 => n4938, A2 => n2910, B1 => n2983, B2 => n2908
                           , ZN => n2083);
   U179 : OAI22_X1 port map( A1 => n5195, A2 => n2910, B1 => n2984, B2 => n2908
                           , ZN => n2082);
   U180 : OAI22_X1 port map( A1 => n4939, A2 => n2910, B1 => n2985, B2 => n2908
                           , ZN => n2081);
   U181 : OAI22_X1 port map( A1 => n4940, A2 => n2910, B1 => n2987, B2 => n2908
                           , ZN => n2080);
   U182 : OAI22_X1 port map( A1 => n4667, A2 => n2910, B1 => n2988, B2 => n2909
                           , ZN => n2079);
   U183 : OAI22_X1 port map( A1 => n4941, A2 => n2910, B1 => n2990, B2 => n2909
                           , ZN => n2078);
   U184 : OAI22_X1 port map( A1 => n4942, A2 => n2910, B1 => n2991, B2 => n2909
                           , ZN => n2077);
   U185 : OAI22_X1 port map( A1 => n5435, A2 => n2910, B1 => n2992, B2 => n2909
                           , ZN => n2076);
   U186 : OAI22_X1 port map( A1 => n5436, A2 => n2910, B1 => n2993, B2 => n2909
                           , ZN => n2075);
   U187 : OAI22_X1 port map( A1 => n4943, A2 => n2910, B1 => n2994, B2 => n2909
                           , ZN => n2074);
   U188 : OAI22_X1 port map( A1 => n5437, A2 => n2910, B1 => n2995, B2 => n2909
                           , ZN => n2073);
   U189 : OAI22_X1 port map( A1 => n4668, A2 => n2910, B1 => n2996, B2 => n2909
                           , ZN => n2072);
   U190 : OAI22_X1 port map( A1 => n5438, A2 => n2910, B1 => n2998, B2 => n2909
                           , ZN => n2071);
   U191 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n2925);
   U192 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n2925, ZN => n3032);
   U193 : NAND2_X1 port map( A1 => n2927, A2 => n3032, ZN => n2911);
   U194 : NAND2_X2 port map( A1 => n2895, A2 => n2911, ZN => n2913);
   U195 : CLKBUF_X1 port map( A => n2911, Z => n2912);
   U196 : OAI22_X1 port map( A1 => n5439, A2 => n2913, B1 => n3050, B2 => n2912
                           , ZN => n2070);
   U197 : OAI22_X1 port map( A1 => n4669, A2 => n2913, B1 => n2965, B2 => n2911
                           , ZN => n2069);
   U198 : OAI22_X1 port map( A1 => n4944, A2 => n2913, B1 => n2966, B2 => n2912
                           , ZN => n2068);
   U199 : OAI22_X1 port map( A1 => n4945, A2 => n2913, B1 => n2967, B2 => n2911
                           , ZN => n2067);
   U200 : OAI22_X1 port map( A1 => n4670, A2 => n2913, B1 => n2968, B2 => n2912
                           , ZN => n2066);
   U201 : OAI22_X1 port map( A1 => n4946, A2 => n2913, B1 => n2969, B2 => n2911
                           , ZN => n2065);
   U202 : OAI22_X1 port map( A1 => n4947, A2 => n2913, B1 => n2970, B2 => n2912
                           , ZN => n2064);
   U203 : OAI22_X1 port map( A1 => n5440, A2 => n2913, B1 => n2971, B2 => n2911
                           , ZN => n2063);
   U204 : OAI22_X1 port map( A1 => n4671, A2 => n2913, B1 => n2972, B2 => n2912
                           , ZN => n2062);
   U205 : OAI22_X1 port map( A1 => n4948, A2 => n2913, B1 => n2973, B2 => n2911
                           , ZN => n2061);
   U206 : OAI22_X1 port map( A1 => n4672, A2 => n2913, B1 => n2974, B2 => n2911
                           , ZN => n2060);
   U207 : OAI22_X1 port map( A1 => n4673, A2 => n2913, B1 => n2975, B2 => n2912
                           , ZN => n2059);
   U208 : OAI22_X1 port map( A1 => n4674, A2 => n2913, B1 => n2976, B2 => n2911
                           , ZN => n2058);
   U209 : OAI22_X1 port map( A1 => n4675, A2 => n2913, B1 => n2977, B2 => n2912
                           , ZN => n2057);
   U210 : OAI22_X1 port map( A1 => n4676, A2 => n2913, B1 => n2978, B2 => n2911
                           , ZN => n2056);
   U211 : OAI22_X1 port map( A1 => n4949, A2 => n2913, B1 => n2979, B2 => n2912
                           , ZN => n2055);
   U212 : OAI22_X1 port map( A1 => n5196, A2 => n2913, B1 => n2980, B2 => n2911
                           , ZN => n2054);
   U213 : OAI22_X1 port map( A1 => n5441, A2 => n2913, B1 => n2981, B2 => n2911
                           , ZN => n2053);
   U214 : OAI22_X1 port map( A1 => n4677, A2 => n2913, B1 => n2982, B2 => n2911
                           , ZN => n2052);
   U215 : OAI22_X1 port map( A1 => n4678, A2 => n2913, B1 => n2983, B2 => n2911
                           , ZN => n2051);
   U216 : OAI22_X1 port map( A1 => n4950, A2 => n2913, B1 => n2984, B2 => n2911
                           , ZN => n2050);
   U217 : OAI22_X1 port map( A1 => n5197, A2 => n2913, B1 => n2985, B2 => n2911
                           , ZN => n2049);
   U218 : OAI22_X1 port map( A1 => n4679, A2 => n2913, B1 => n2987, B2 => n2911
                           , ZN => n2048);
   U219 : OAI22_X1 port map( A1 => n4680, A2 => n2913, B1 => n2988, B2 => n2912
                           , ZN => n2047);
   U220 : OAI22_X1 port map( A1 => n5442, A2 => n2913, B1 => n2990, B2 => n2912
                           , ZN => n2046);
   U221 : OAI22_X1 port map( A1 => n4681, A2 => n2913, B1 => n2991, B2 => n2912
                           , ZN => n2045);
   U222 : OAI22_X1 port map( A1 => n4951, A2 => n2913, B1 => n2992, B2 => n2912
                           , ZN => n2044);
   U223 : OAI22_X1 port map( A1 => n4682, A2 => n2913, B1 => n2993, B2 => n2912
                           , ZN => n2043);
   U224 : OAI22_X1 port map( A1 => n4952, A2 => n2913, B1 => n2994, B2 => n2912
                           , ZN => n2042);
   U225 : OAI22_X1 port map( A1 => n4953, A2 => n2913, B1 => n2995, B2 => n2912
                           , ZN => n2041);
   U226 : OAI22_X1 port map( A1 => n4683, A2 => n2913, B1 => n2996, B2 => n2912
                           , ZN => n2040);
   U227 : OAI22_X1 port map( A1 => n4684, A2 => n2913, B1 => n2998, B2 => n2912
                           , ZN => n2039);
   U228 : INV_X1 port map( A => ADD_WR(2), ZN => n2926);
   U229 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n2926, ZN 
                           => n3036);
   U230 : NAND2_X1 port map( A1 => n2927, A2 => n3036, ZN => n2914);
   U231 : OAI22_X1 port map( A1 => n5443, A2 => n2916, B1 => n3014, B2 => n2915
                           , ZN => n2038);
   U232 : OAI22_X1 port map( A1 => n4685, A2 => n2916, B1 => n2965, B2 => n2914
                           , ZN => n2037);
   U233 : OAI22_X1 port map( A1 => n5198, A2 => n2916, B1 => n2966, B2 => n2915
                           , ZN => n2036);
   U234 : OAI22_X1 port map( A1 => n5444, A2 => n2916, B1 => n2967, B2 => n2914
                           , ZN => n2035);
   U235 : OAI22_X1 port map( A1 => n5199, A2 => n2916, B1 => n2968, B2 => n2915
                           , ZN => n2034);
   U236 : OAI22_X1 port map( A1 => n5200, A2 => n2916, B1 => n2969, B2 => n2914
                           , ZN => n2033);
   U237 : OAI22_X1 port map( A1 => n5201, A2 => n2916, B1 => n2970, B2 => n2915
                           , ZN => n2032);
   U238 : OAI22_X1 port map( A1 => n5445, A2 => n2916, B1 => n2971, B2 => n2914
                           , ZN => n2031);
   U239 : OAI22_X1 port map( A1 => n5202, A2 => n2916, B1 => n2972, B2 => n2915
                           , ZN => n2030);
   U240 : OAI22_X1 port map( A1 => n5446, A2 => n2916, B1 => n2973, B2 => n2914
                           , ZN => n2029);
   U241 : OAI22_X1 port map( A1 => n4686, A2 => n2916, B1 => n2974, B2 => n2914
                           , ZN => n2028);
   U242 : OAI22_X1 port map( A1 => n5203, A2 => n2916, B1 => n2975, B2 => n2915
                           , ZN => n2027);
   U243 : OAI22_X1 port map( A1 => n5447, A2 => n2916, B1 => n2976, B2 => n2914
                           , ZN => n2026);
   U244 : OAI22_X1 port map( A1 => n5204, A2 => n2916, B1 => n2977, B2 => n2915
                           , ZN => n2025);
   U245 : OAI22_X1 port map( A1 => n5448, A2 => n2916, B1 => n2978, B2 => n2914
                           , ZN => n2024);
   U246 : OAI22_X1 port map( A1 => n5205, A2 => n2916, B1 => n2979, B2 => n2915
                           , ZN => n2023);
   U247 : OAI22_X1 port map( A1 => n5449, A2 => n2916, B1 => n2980, B2 => n2914
                           , ZN => n2022);
   U248 : OAI22_X1 port map( A1 => n5206, A2 => n2916, B1 => n2981, B2 => n2914
                           , ZN => n2021);
   U249 : OAI22_X1 port map( A1 => n5207, A2 => n2916, B1 => n2982, B2 => n2914
                           , ZN => n2020);
   U250 : OAI22_X1 port map( A1 => n5450, A2 => n2916, B1 => n2983, B2 => n2914
                           , ZN => n2019);
   U251 : OAI22_X1 port map( A1 => n4687, A2 => n2916, B1 => n2984, B2 => n2914
                           , ZN => n2018);
   U252 : OAI22_X1 port map( A1 => n5451, A2 => n2916, B1 => n2985, B2 => n2914
                           , ZN => n2017);
   U253 : OAI22_X1 port map( A1 => n5208, A2 => n2916, B1 => n2987, B2 => n2914
                           , ZN => n2016);
   U254 : OAI22_X1 port map( A1 => n5209, A2 => n2916, B1 => n2988, B2 => n2915
                           , ZN => n2015);
   U255 : OAI22_X1 port map( A1 => n5210, A2 => n2916, B1 => n2990, B2 => n2915
                           , ZN => n2014);
   U256 : OAI22_X1 port map( A1 => n5211, A2 => n2916, B1 => n2991, B2 => n2915
                           , ZN => n2013);
   U257 : OAI22_X1 port map( A1 => n4688, A2 => n2916, B1 => n2992, B2 => n2915
                           , ZN => n2012);
   U258 : OAI22_X1 port map( A1 => n5452, A2 => n2916, B1 => n2993, B2 => n2915
                           , ZN => n2011);
   U259 : OAI22_X1 port map( A1 => n5453, A2 => n2916, B1 => n2994, B2 => n2915
                           , ZN => n2010);
   U260 : OAI22_X1 port map( A1 => n4954, A2 => n2916, B1 => n2995, B2 => n2915
                           , ZN => n2009);
   U261 : OAI22_X1 port map( A1 => n4689, A2 => n2916, B1 => n2996, B2 => n2915
                           , ZN => n2008);
   U262 : OAI22_X1 port map( A1 => n5212, A2 => n2916, B1 => n2998, B2 => n2915
                           , ZN => n2007);
   U263 : NAND2_X1 port map( A1 => n2927, A2 => n3040, ZN => n2918);
   U264 : CLKBUF_X1 port map( A => n2918, Z => n2919);
   U265 : OAI22_X1 port map( A1 => n4690, A2 => n2920, B1 => n3050, B2 => n2919
                           , ZN => n2006);
   U266 : OAI22_X1 port map( A1 => n5454, A2 => n2920, B1 => n2965, B2 => n2918
                           , ZN => n2005);
   U267 : OAI22_X1 port map( A1 => n4691, A2 => n2920, B1 => n2966, B2 => n2919
                           , ZN => n2004);
   U268 : OAI22_X1 port map( A1 => n4955, A2 => n2920, B1 => n2967, B2 => n2918
                           , ZN => n2003);
   U269 : OAI22_X1 port map( A1 => n5213, A2 => n2920, B1 => n2968, B2 => n2919
                           , ZN => n2002);
   U270 : OAI22_X1 port map( A1 => n5214, A2 => n2920, B1 => n2969, B2 => n2918
                           , ZN => n2001);
   U271 : OAI22_X1 port map( A1 => n4692, A2 => n2920, B1 => n2970, B2 => n2919
                           , ZN => n2000);
   U272 : OAI22_X1 port map( A1 => n5215, A2 => n2920, B1 => n2971, B2 => n2918
                           , ZN => n1999);
   U273 : OAI22_X1 port map( A1 => n5455, A2 => n2920, B1 => n2972, B2 => n2919
                           , ZN => n1998);
   U274 : OAI22_X1 port map( A1 => n5216, A2 => n2920, B1 => n2973, B2 => n2918
                           , ZN => n1997);
   U275 : OAI22_X1 port map( A1 => n5217, A2 => n2920, B1 => n2974, B2 => n2918
                           , ZN => n1996);
   U276 : OAI22_X1 port map( A1 => n5218, A2 => n2920, B1 => n2975, B2 => n2919
                           , ZN => n1995);
   U277 : OAI22_X1 port map( A1 => n5456, A2 => n2920, B1 => n2976, B2 => n2918
                           , ZN => n1994);
   U278 : OAI22_X1 port map( A1 => n4956, A2 => n2920, B1 => n2977, B2 => n2919
                           , ZN => n1993);
   U279 : OAI22_X1 port map( A1 => n5219, A2 => n2920, B1 => n2978, B2 => n2918
                           , ZN => n1992);
   U280 : OAI22_X1 port map( A1 => n5220, A2 => n2920, B1 => n2979, B2 => n2919
                           , ZN => n1991);
   U281 : OAI22_X1 port map( A1 => n4957, A2 => n2920, B1 => n2980, B2 => n2918
                           , ZN => n1990);
   U282 : OAI22_X1 port map( A1 => n4693, A2 => n2920, B1 => n2981, B2 => n2918
                           , ZN => n1989);
   U283 : OAI22_X1 port map( A1 => n5457, A2 => n2920, B1 => n2982, B2 => n2918
                           , ZN => n1988);
   U284 : OAI22_X1 port map( A1 => n5458, A2 => n2920, B1 => n2983, B2 => n2918
                           , ZN => n1987);
   U285 : OAI22_X1 port map( A1 => n5221, A2 => n2920, B1 => n2984, B2 => n2918
                           , ZN => n1986);
   U286 : OAI22_X1 port map( A1 => n5459, A2 => n2920, B1 => n2985, B2 => n2918
                           , ZN => n1985);
   U287 : OAI22_X1 port map( A1 => n5222, A2 => n2920, B1 => n2987, B2 => n2918
                           , ZN => n1984);
   U288 : OAI22_X1 port map( A1 => n5460, A2 => n2920, B1 => n2988, B2 => n2919
                           , ZN => n1983);
   U289 : OAI22_X1 port map( A1 => n5461, A2 => n2920, B1 => n2990, B2 => n2919
                           , ZN => n1982);
   U290 : OAI22_X1 port map( A1 => n4958, A2 => n2920, B1 => n2991, B2 => n2919
                           , ZN => n1981);
   U291 : OAI22_X1 port map( A1 => n5223, A2 => n2920, B1 => n2992, B2 => n2919
                           , ZN => n1980);
   U292 : OAI22_X1 port map( A1 => n5224, A2 => n2920, B1 => n2993, B2 => n2919
                           , ZN => n1979);
   U293 : OAI22_X1 port map( A1 => n5225, A2 => n2920, B1 => n2994, B2 => n2919
                           , ZN => n1978);
   U294 : OAI22_X1 port map( A1 => n5226, A2 => n2920, B1 => n2995, B2 => n2919
                           , ZN => n1977);
   U295 : OAI22_X1 port map( A1 => n5462, A2 => n2920, B1 => n2996, B2 => n2919
                           , ZN => n1976);
   U296 : OAI22_X1 port map( A1 => n5463, A2 => n2920, B1 => n2998, B2 => n2919
                           , ZN => n1975);
   U297 : NOR2_X1 port map( A1 => n2926, A2 => n2921, ZN => n3044);
   U298 : NAND2_X1 port map( A1 => n2927, A2 => n3044, ZN => n2922);
   U299 : CLKBUF_X1 port map( A => n2922, Z => n2923);
   U300 : OAI22_X1 port map( A1 => n5227, A2 => n2924, B1 => n3014, B2 => n2923
                           , ZN => n1974);
   U301 : OAI22_X1 port map( A1 => n4959, A2 => n2924, B1 => n2965, B2 => n2922
                           , ZN => n1973);
   U302 : OAI22_X1 port map( A1 => n5464, A2 => n2924, B1 => n2966, B2 => n2923
                           , ZN => n1972);
   U303 : OAI22_X1 port map( A1 => n5465, A2 => n2924, B1 => n2967, B2 => n2922
                           , ZN => n1971);
   U304 : OAI22_X1 port map( A1 => n4694, A2 => n2924, B1 => n2968, B2 => n2923
                           , ZN => n1970);
   U305 : OAI22_X1 port map( A1 => n4695, A2 => n2924, B1 => n2969, B2 => n2922
                           , ZN => n1969);
   U306 : OAI22_X1 port map( A1 => n5466, A2 => n2924, B1 => n2970, B2 => n2923
                           , ZN => n1968);
   U307 : OAI22_X1 port map( A1 => n4696, A2 => n2924, B1 => n2971, B2 => n2922
                           , ZN => n1967);
   U308 : OAI22_X1 port map( A1 => n4697, A2 => n2924, B1 => n2972, B2 => n2923
                           , ZN => n1966);
   U309 : OAI22_X1 port map( A1 => n4960, A2 => n2924, B1 => n2973, B2 => n2922
                           , ZN => n1965);
   U310 : OAI22_X1 port map( A1 => n5467, A2 => n2924, B1 => n2974, B2 => n2922
                           , ZN => n1964);
   U311 : OAI22_X1 port map( A1 => n4961, A2 => n2924, B1 => n2975, B2 => n2923
                           , ZN => n1963);
   U312 : OAI22_X1 port map( A1 => n4698, A2 => n2924, B1 => n2976, B2 => n2922
                           , ZN => n1962);
   U313 : OAI22_X1 port map( A1 => n5468, A2 => n2924, B1 => n2977, B2 => n2923
                           , ZN => n1961);
   U314 : OAI22_X1 port map( A1 => n4962, A2 => n2924, B1 => n2978, B2 => n2922
                           , ZN => n1960);
   U315 : OAI22_X1 port map( A1 => n4699, A2 => n2924, B1 => n2979, B2 => n2923
                           , ZN => n1959);
   U316 : OAI22_X1 port map( A1 => n5228, A2 => n2924, B1 => n2980, B2 => n2922
                           , ZN => n1958);
   U317 : OAI22_X1 port map( A1 => n4963, A2 => n2924, B1 => n2981, B2 => n2922
                           , ZN => n1957);
   U318 : OAI22_X1 port map( A1 => n4964, A2 => n2924, B1 => n2982, B2 => n2922
                           , ZN => n1956);
   U319 : OAI22_X1 port map( A1 => n5229, A2 => n2924, B1 => n2983, B2 => n2922
                           , ZN => n1955);
   U320 : OAI22_X1 port map( A1 => n5469, A2 => n2924, B1 => n2984, B2 => n2922
                           , ZN => n1954);
   U321 : OAI22_X1 port map( A1 => n4965, A2 => n2924, B1 => n2985, B2 => n2922
                           , ZN => n1953);
   U322 : OAI22_X1 port map( A1 => n4966, A2 => n2924, B1 => n2987, B2 => n2922
                           , ZN => n1952);
   U323 : OAI22_X1 port map( A1 => n5470, A2 => n2924, B1 => n2988, B2 => n2923
                           , ZN => n1951);
   U324 : OAI22_X1 port map( A1 => n4700, A2 => n2924, B1 => n2990, B2 => n2923
                           , ZN => n1950);
   U325 : OAI22_X1 port map( A1 => n5471, A2 => n2924, B1 => n2991, B2 => n2923
                           , ZN => n1949);
   U326 : OAI22_X1 port map( A1 => n4701, A2 => n2924, B1 => n2992, B2 => n2923
                           , ZN => n1948);
   U327 : OAI22_X1 port map( A1 => n4967, A2 => n2924, B1 => n2993, B2 => n2923
                           , ZN => n1947);
   U328 : OAI22_X1 port map( A1 => n4702, A2 => n2924, B1 => n2994, B2 => n2923
                           , ZN => n1946);
   U329 : OAI22_X1 port map( A1 => n5230, A2 => n2924, B1 => n2995, B2 => n2923
                           , ZN => n1945);
   U330 : OAI22_X1 port map( A1 => n5472, A2 => n2924, B1 => n2996, B2 => n2923
                           , ZN => n1944);
   U331 : OAI22_X1 port map( A1 => n4968, A2 => n2924, B1 => n2998, B2 => n2923
                           , ZN => n1943);
   U332 : NOR2_X1 port map( A1 => n2926, A2 => n2925, ZN => n3049);
   U333 : NAND2_X1 port map( A1 => n2927, A2 => n3049, ZN => n2928);
   U334 : CLKBUF_X1 port map( A => n2931, Z => n2929);
   U335 : CLKBUF_X1 port map( A => n2928, Z => n2930);
   U336 : OAI22_X1 port map( A1 => n4969, A2 => n2929, B1 => n3050, B2 => n2930
                           , ZN => n1942);
   U337 : OAI22_X1 port map( A1 => n4703, A2 => n2931, B1 => n2965, B2 => n2928
                           , ZN => n1941);
   U338 : OAI22_X1 port map( A1 => n4704, A2 => n2929, B1 => n2966, B2 => n2930
                           , ZN => n1940);
   U339 : OAI22_X1 port map( A1 => n4705, A2 => n2931, B1 => n2967, B2 => n2928
                           , ZN => n1939);
   U340 : OAI22_X1 port map( A1 => n4970, A2 => n2929, B1 => n2968, B2 => n2930
                           , ZN => n1938);
   U341 : OAI22_X1 port map( A1 => n4971, A2 => n2931, B1 => n2969, B2 => n2928
                           , ZN => n1937);
   U342 : OAI22_X1 port map( A1 => n4706, A2 => n2929, B1 => n2970, B2 => n2930
                           , ZN => n1936);
   U343 : OAI22_X1 port map( A1 => n4972, A2 => n2931, B1 => n2971, B2 => n2928
                           , ZN => n1935);
   U344 : OAI22_X1 port map( A1 => n4973, A2 => n2929, B1 => n2972, B2 => n2930
                           , ZN => n1934);
   U345 : OAI22_X1 port map( A1 => n4707, A2 => n2931, B1 => n2973, B2 => n2928
                           , ZN => n1933);
   U346 : OAI22_X1 port map( A1 => n4974, A2 => n2931, B1 => n2974, B2 => n2928
                           , ZN => n1932);
   U347 : OAI22_X1 port map( A1 => n4975, A2 => n2931, B1 => n2975, B2 => n2930
                           , ZN => n1931);
   U348 : OAI22_X1 port map( A1 => n4976, A2 => n2929, B1 => n2976, B2 => n2928
                           , ZN => n1930);
   U349 : OAI22_X1 port map( A1 => n4708, A2 => n2929, B1 => n2977, B2 => n2930
                           , ZN => n1929);
   U350 : OAI22_X1 port map( A1 => n4977, A2 => n2929, B1 => n2978, B2 => n2928
                           , ZN => n1928);
   U351 : OAI22_X1 port map( A1 => n4978, A2 => n2929, B1 => n2979, B2 => n2930
                           , ZN => n1927);
   U352 : OAI22_X1 port map( A1 => n4709, A2 => n2929, B1 => n2980, B2 => n2928
                           , ZN => n1926);
   U353 : OAI22_X1 port map( A1 => n4710, A2 => n2929, B1 => n2981, B2 => n2928
                           , ZN => n1925);
   U354 : OAI22_X1 port map( A1 => n4979, A2 => n2929, B1 => n2982, B2 => n2928
                           , ZN => n1924);
   U355 : OAI22_X1 port map( A1 => n4711, A2 => n2929, B1 => n2983, B2 => n2928
                           , ZN => n1923);
   U356 : OAI22_X1 port map( A1 => n4712, A2 => n2929, B1 => n2984, B2 => n2928
                           , ZN => n1922);
   U357 : OAI22_X1 port map( A1 => n4713, A2 => n2929, B1 => n2985, B2 => n2928
                           , ZN => n1921);
   U358 : OAI22_X1 port map( A1 => n4980, A2 => n2929, B1 => n2987, B2 => n2928
                           , ZN => n1920);
   U359 : OAI22_X1 port map( A1 => n4981, A2 => n2929, B1 => n2988, B2 => n2930
                           , ZN => n1919);
   U360 : OAI22_X1 port map( A1 => n4714, A2 => n2931, B1 => n2990, B2 => n2930
                           , ZN => n1918);
   U361 : OAI22_X1 port map( A1 => n4715, A2 => n2931, B1 => n2991, B2 => n2930
                           , ZN => n1917);
   U362 : OAI22_X1 port map( A1 => n4982, A2 => n2931, B1 => n2992, B2 => n2930
                           , ZN => n1916);
   U363 : OAI22_X1 port map( A1 => n4983, A2 => n2931, B1 => n2993, B2 => n2930
                           , ZN => n1915);
   U364 : OAI22_X1 port map( A1 => n4716, A2 => n2931, B1 => n2994, B2 => n2930
                           , ZN => n1914);
   U365 : OAI22_X1 port map( A1 => n4984, A2 => n2931, B1 => n2995, B2 => n2930
                           , ZN => n1913);
   U366 : OAI22_X1 port map( A1 => n4985, A2 => n2931, B1 => n2996, B2 => n2930
                           , ZN => n1912);
   U367 : OAI22_X1 port map( A1 => n4986, A2 => n2931, B1 => n2998, B2 => n2930
                           , ZN => n1911);
   U368 : NOR2_X1 port map( A1 => n3019, A2 => n2932, ZN => n2955);
   U369 : NAND2_X1 port map( A1 => n3020, A2 => n2955, ZN => n2933);
   U370 : CLKBUF_X1 port map( A => n2933, Z => n2934);
   U371 : OAI22_X1 port map( A1 => n5473, A2 => n2935, B1 => n3014, B2 => n2934
                           , ZN => n1910);
   U372 : OAI22_X1 port map( A1 => n5474, A2 => n2935, B1 => n2965, B2 => n2933
                           , ZN => n1909);
   U373 : OAI22_X1 port map( A1 => n5231, A2 => n2935, B1 => n2966, B2 => n2934
                           , ZN => n1908);
   U374 : OAI22_X1 port map( A1 => n5232, A2 => n2935, B1 => n2967, B2 => n2933
                           , ZN => n1907);
   U375 : OAI22_X1 port map( A1 => n5475, A2 => n2935, B1 => n2968, B2 => n2934
                           , ZN => n1906);
   U376 : OAI22_X1 port map( A1 => n5233, A2 => n2935, B1 => n2969, B2 => n2933
                           , ZN => n1905);
   U377 : OAI22_X1 port map( A1 => n5476, A2 => n2935, B1 => n2970, B2 => n2934
                           , ZN => n1904);
   U378 : OAI22_X1 port map( A1 => n5234, A2 => n2935, B1 => n2971, B2 => n2933
                           , ZN => n1903);
   U379 : OAI22_X1 port map( A1 => n5235, A2 => n2935, B1 => n2972, B2 => n2934
                           , ZN => n1902);
   U380 : OAI22_X1 port map( A1 => n5236, A2 => n2935, B1 => n2973, B2 => n2933
                           , ZN => n1901);
   U381 : OAI22_X1 port map( A1 => n5477, A2 => n2935, B1 => n2974, B2 => n2933
                           , ZN => n1900);
   U382 : OAI22_X1 port map( A1 => n5478, A2 => n2935, B1 => n2975, B2 => n2934
                           , ZN => n1899);
   U383 : OAI22_X1 port map( A1 => n5237, A2 => n2935, B1 => n2976, B2 => n2933
                           , ZN => n1898);
   U384 : OAI22_X1 port map( A1 => n5238, A2 => n2935, B1 => n2977, B2 => n2934
                           , ZN => n1897);
   U385 : OAI22_X1 port map( A1 => n5239, A2 => n2935, B1 => n2978, B2 => n2933
                           , ZN => n1896);
   U386 : OAI22_X1 port map( A1 => n5240, A2 => n2935, B1 => n2979, B2 => n2934
                           , ZN => n1895);
   U387 : OAI22_X1 port map( A1 => n5479, A2 => n2935, B1 => n2980, B2 => n2933
                           , ZN => n1894);
   U388 : OAI22_X1 port map( A1 => n5480, A2 => n2935, B1 => n2981, B2 => n2933
                           , ZN => n1893);
   U389 : OAI22_X1 port map( A1 => n5481, A2 => n2935, B1 => n2982, B2 => n2933
                           , ZN => n1892);
   U390 : OAI22_X1 port map( A1 => n5482, A2 => n2935, B1 => n2983, B2 => n2933
                           , ZN => n1891);
   U391 : OAI22_X1 port map( A1 => n5241, A2 => n2935, B1 => n2984, B2 => n2933
                           , ZN => n1890);
   U392 : OAI22_X1 port map( A1 => n5242, A2 => n2935, B1 => n2985, B2 => n2933
                           , ZN => n1889);
   U393 : OAI22_X1 port map( A1 => n5243, A2 => n2935, B1 => n2987, B2 => n2933
                           , ZN => n1888);
   U394 : OAI22_X1 port map( A1 => n5244, A2 => n2935, B1 => n2988, B2 => n2934
                           , ZN => n1887);
   U395 : OAI22_X1 port map( A1 => n5483, A2 => n2935, B1 => n2990, B2 => n2934
                           , ZN => n1886);
   U396 : OAI22_X1 port map( A1 => n5245, A2 => n2935, B1 => n2991, B2 => n2934
                           , ZN => n1885);
   U397 : OAI22_X1 port map( A1 => n5484, A2 => n2935, B1 => n2992, B2 => n2934
                           , ZN => n1884);
   U398 : OAI22_X1 port map( A1 => n5246, A2 => n2935, B1 => n2993, B2 => n2934
                           , ZN => n1883);
   U399 : OAI22_X1 port map( A1 => n5485, A2 => n2935, B1 => n2994, B2 => n2934
                           , ZN => n1882);
   U400 : OAI22_X1 port map( A1 => n5247, A2 => n2935, B1 => n2995, B2 => n2934
                           , ZN => n1881);
   U401 : OAI22_X1 port map( A1 => n5248, A2 => n2935, B1 => n2996, B2 => n2934
                           , ZN => n1880);
   U402 : OAI22_X1 port map( A1 => n5486, A2 => n2935, B1 => n2998, B2 => n2934
                           , ZN => n1879);
   U403 : NAND2_X1 port map( A1 => n3024, A2 => n2955, ZN => n2936);
   U404 : CLKBUF_X1 port map( A => n2936, Z => n2937);
   U405 : OAI22_X1 port map( A1 => n4717, A2 => n2938, B1 => n3050, B2 => n2937
                           , ZN => n1878);
   U406 : OAI22_X1 port map( A1 => n5487, A2 => n2938, B1 => n2965, B2 => n2936
                           , ZN => n1877);
   U407 : OAI22_X1 port map( A1 => n4718, A2 => n2938, B1 => n2966, B2 => n2937
                           , ZN => n1876);
   U408 : OAI22_X1 port map( A1 => n4987, A2 => n2938, B1 => n2967, B2 => n2936
                           , ZN => n1875);
   U409 : OAI22_X1 port map( A1 => n4988, A2 => n2938, B1 => n2968, B2 => n2937
                           , ZN => n1874);
   U410 : OAI22_X1 port map( A1 => n4719, A2 => n2938, B1 => n2969, B2 => n2936
                           , ZN => n1873);
   U411 : OAI22_X1 port map( A1 => n4720, A2 => n2938, B1 => n2970, B2 => n2937
                           , ZN => n1872);
   U412 : OAI22_X1 port map( A1 => n4989, A2 => n2938, B1 => n2971, B2 => n2936
                           , ZN => n1871);
   U413 : OAI22_X1 port map( A1 => n4990, A2 => n2938, B1 => n2972, B2 => n2937
                           , ZN => n1870);
   U414 : OAI22_X1 port map( A1 => n5249, A2 => n2938, B1 => n2973, B2 => n2936
                           , ZN => n1869);
   U415 : OAI22_X1 port map( A1 => n5488, A2 => n2938, B1 => n2974, B2 => n2936
                           , ZN => n1868);
   U416 : OAI22_X1 port map( A1 => n5489, A2 => n2938, B1 => n2975, B2 => n2937
                           , ZN => n1867);
   U417 : OAI22_X1 port map( A1 => n4721, A2 => n2938, B1 => n2976, B2 => n2936
                           , ZN => n1866);
   U418 : OAI22_X1 port map( A1 => n5490, A2 => n2938, B1 => n2977, B2 => n2937
                           , ZN => n1865);
   U419 : OAI22_X1 port map( A1 => n5250, A2 => n2938, B1 => n2978, B2 => n2936
                           , ZN => n1864);
   U420 : OAI22_X1 port map( A1 => n4722, A2 => n2938, B1 => n2979, B2 => n2937
                           , ZN => n1863);
   U421 : OAI22_X1 port map( A1 => n4991, A2 => n2938, B1 => n2980, B2 => n2936
                           , ZN => n1862);
   U422 : OAI22_X1 port map( A1 => n4723, A2 => n2938, B1 => n2981, B2 => n2936
                           , ZN => n1861);
   U423 : OAI22_X1 port map( A1 => n5251, A2 => n2938, B1 => n2982, B2 => n2936
                           , ZN => n1860);
   U424 : OAI22_X1 port map( A1 => n4992, A2 => n2938, B1 => n2983, B2 => n2936
                           , ZN => n1859);
   U425 : OAI22_X1 port map( A1 => n4724, A2 => n2938, B1 => n2984, B2 => n2936
                           , ZN => n1858);
   U426 : OAI22_X1 port map( A1 => n5491, A2 => n2938, B1 => n2985, B2 => n2936
                           , ZN => n1857);
   U427 : OAI22_X1 port map( A1 => n5492, A2 => n2938, B1 => n2987, B2 => n2936
                           , ZN => n1856);
   U428 : OAI22_X1 port map( A1 => n5493, A2 => n2938, B1 => n2988, B2 => n2937
                           , ZN => n1855);
   U429 : OAI22_X1 port map( A1 => n5494, A2 => n2938, B1 => n2990, B2 => n2937
                           , ZN => n1854);
   U430 : OAI22_X1 port map( A1 => n5495, A2 => n2938, B1 => n2991, B2 => n2937
                           , ZN => n1853);
   U431 : OAI22_X1 port map( A1 => n5252, A2 => n2938, B1 => n2992, B2 => n2937
                           , ZN => n1852);
   U432 : OAI22_X1 port map( A1 => n5496, A2 => n2938, B1 => n2993, B2 => n2937
                           , ZN => n1851);
   U433 : OAI22_X1 port map( A1 => n5253, A2 => n2938, B1 => n2994, B2 => n2937
                           , ZN => n1850);
   U434 : OAI22_X1 port map( A1 => n5497, A2 => n2938, B1 => n2995, B2 => n2937
                           , ZN => n1849);
   U435 : OAI22_X1 port map( A1 => n4725, A2 => n2938, B1 => n2996, B2 => n2937
                           , ZN => n1848);
   U436 : OAI22_X1 port map( A1 => n4726, A2 => n2938, B1 => n2998, B2 => n2937
                           , ZN => n1847);
   U437 : NAND2_X1 port map( A1 => n3028, A2 => n2955, ZN => n2939);
   U438 : CLKBUF_X1 port map( A => n2939, Z => n2940);
   U439 : OAI22_X1 port map( A1 => n4727, A2 => n2941, B1 => n3050, B2 => n2940
                           , ZN => n1846);
   U440 : OAI22_X1 port map( A1 => n4993, A2 => n2941, B1 => n2965, B2 => n2939
                           , ZN => n1845);
   U441 : OAI22_X1 port map( A1 => n4728, A2 => n2941, B1 => n2966, B2 => n2940
                           , ZN => n1844);
   U442 : OAI22_X1 port map( A1 => n4729, A2 => n2941, B1 => n2967, B2 => n2939
                           , ZN => n1843);
   U443 : OAI22_X1 port map( A1 => n5254, A2 => n2941, B1 => n2968, B2 => n2940
                           , ZN => n1842);
   U444 : OAI22_X1 port map( A1 => n4730, A2 => n2941, B1 => n2969, B2 => n2939
                           , ZN => n1841);
   U445 : OAI22_X1 port map( A1 => n4731, A2 => n2941, B1 => n2970, B2 => n2940
                           , ZN => n1840);
   U446 : OAI22_X1 port map( A1 => n4994, A2 => n2941, B1 => n2971, B2 => n2939
                           , ZN => n1839);
   U447 : OAI22_X1 port map( A1 => n5255, A2 => n2941, B1 => n2972, B2 => n2940
                           , ZN => n1838);
   U448 : OAI22_X1 port map( A1 => n4732, A2 => n2941, B1 => n2973, B2 => n2939
                           , ZN => n1837);
   U449 : OAI22_X1 port map( A1 => n4995, A2 => n2941, B1 => n2974, B2 => n2939
                           , ZN => n1836);
   U450 : OAI22_X1 port map( A1 => n4733, A2 => n2941, B1 => n2975, B2 => n2940
                           , ZN => n1835);
   U451 : OAI22_X1 port map( A1 => n4734, A2 => n2941, B1 => n2976, B2 => n2939
                           , ZN => n1834);
   U452 : OAI22_X1 port map( A1 => n4735, A2 => n2941, B1 => n2977, B2 => n2940
                           , ZN => n1833);
   U453 : OAI22_X1 port map( A1 => n4996, A2 => n2941, B1 => n2978, B2 => n2939
                           , ZN => n1832);
   U454 : OAI22_X1 port map( A1 => n4997, A2 => n2941, B1 => n2979, B2 => n2940
                           , ZN => n1831);
   U455 : OAI22_X1 port map( A1 => n4736, A2 => n2941, B1 => n2980, B2 => n2939
                           , ZN => n1830);
   U456 : OAI22_X1 port map( A1 => n4998, A2 => n2941, B1 => n2981, B2 => n2939
                           , ZN => n1829);
   U457 : OAI22_X1 port map( A1 => n4737, A2 => n2941, B1 => n2982, B2 => n2939
                           , ZN => n1828);
   U458 : OAI22_X1 port map( A1 => n4738, A2 => n2941, B1 => n2983, B2 => n2939
                           , ZN => n1827);
   U459 : OAI22_X1 port map( A1 => n4999, A2 => n2941, B1 => n2984, B2 => n2939
                           , ZN => n1826);
   U460 : OAI22_X1 port map( A1 => n5000, A2 => n2941, B1 => n2985, B2 => n2939
                           , ZN => n1825);
   U461 : OAI22_X1 port map( A1 => n5001, A2 => n2941, B1 => n2987, B2 => n2939
                           , ZN => n1824);
   U462 : OAI22_X1 port map( A1 => n4739, A2 => n2941, B1 => n2988, B2 => n2940
                           , ZN => n1823);
   U463 : OAI22_X1 port map( A1 => n4740, A2 => n2941, B1 => n2990, B2 => n2940
                           , ZN => n1822);
   U464 : OAI22_X1 port map( A1 => n4741, A2 => n2941, B1 => n2991, B2 => n2940
                           , ZN => n1821);
   U465 : OAI22_X1 port map( A1 => n4742, A2 => n2941, B1 => n2992, B2 => n2940
                           , ZN => n1820);
   U466 : OAI22_X1 port map( A1 => n4743, A2 => n2941, B1 => n2993, B2 => n2940
                           , ZN => n1819);
   U467 : OAI22_X1 port map( A1 => n4744, A2 => n2941, B1 => n2994, B2 => n2940
                           , ZN => n1818);
   U468 : OAI22_X1 port map( A1 => n5002, A2 => n2941, B1 => n2995, B2 => n2940
                           , ZN => n1817);
   U469 : OAI22_X1 port map( A1 => n5498, A2 => n2941, B1 => n2996, B2 => n2940
                           , ZN => n1816);
   U470 : OAI22_X1 port map( A1 => n4745, A2 => n2941, B1 => n2998, B2 => n2940
                           , ZN => n1815);
   U471 : NAND2_X1 port map( A1 => n3032, A2 => n2955, ZN => n2942);
   U472 : CLKBUF_X1 port map( A => n2945, Z => n2943);
   U473 : CLKBUF_X1 port map( A => n2942, Z => n2944);
   U474 : OAI22_X1 port map( A1 => n5256, A2 => n2943, B1 => n3050, B2 => n2944
                           , ZN => n1814);
   U475 : CLKBUF_X1 port map( A => n2965, Z => n3051);
   U476 : OAI22_X1 port map( A1 => n4746, A2 => n2945, B1 => n3051, B2 => n2942
                           , ZN => n1813);
   U477 : CLKBUF_X1 port map( A => n2966, Z => n3052);
   U478 : OAI22_X1 port map( A1 => n5003, A2 => n2943, B1 => n3052, B2 => n2944
                           , ZN => n1812);
   U479 : CLKBUF_X1 port map( A => n2967, Z => n3053);
   U480 : OAI22_X1 port map( A1 => n5004, A2 => n2945, B1 => n3053, B2 => n2942
                           , ZN => n1811);
   U481 : CLKBUF_X1 port map( A => n2968, Z => n3054);
   U482 : OAI22_X1 port map( A1 => n5005, A2 => n2943, B1 => n3054, B2 => n2944
                           , ZN => n1810);
   U483 : CLKBUF_X1 port map( A => n2969, Z => n3055);
   U484 : OAI22_X1 port map( A1 => n5499, A2 => n2945, B1 => n3055, B2 => n2942
                           , ZN => n1809);
   U485 : CLKBUF_X1 port map( A => n2970, Z => n3056);
   U486 : OAI22_X1 port map( A1 => n5006, A2 => n2943, B1 => n3056, B2 => n2944
                           , ZN => n1808);
   U487 : CLKBUF_X1 port map( A => n2971, Z => n3057);
   U488 : OAI22_X1 port map( A1 => n5007, A2 => n2945, B1 => n3057, B2 => n2942
                           , ZN => n1807);
   U489 : CLKBUF_X1 port map( A => n2972, Z => n3058);
   U490 : OAI22_X1 port map( A1 => n5008, A2 => n2943, B1 => n3058, B2 => n2944
                           , ZN => n1806);
   U491 : CLKBUF_X1 port map( A => n2973, Z => n3059);
   U492 : OAI22_X1 port map( A1 => n5500, A2 => n2945, B1 => n3059, B2 => n2942
                           , ZN => n1805);
   U493 : CLKBUF_X1 port map( A => n2974, Z => n3060);
   U494 : OAI22_X1 port map( A1 => n4747, A2 => n2945, B1 => n3060, B2 => n2942
                           , ZN => n1804);
   U495 : CLKBUF_X1 port map( A => n2975, Z => n3061);
   U496 : OAI22_X1 port map( A1 => n5009, A2 => n2945, B1 => n3061, B2 => n2944
                           , ZN => n1803);
   U497 : CLKBUF_X1 port map( A => n2976, Z => n3062);
   U498 : OAI22_X1 port map( A1 => n5501, A2 => n2943, B1 => n3062, B2 => n2942
                           , ZN => n1802);
   U499 : CLKBUF_X1 port map( A => n2977, Z => n3063);
   U500 : OAI22_X1 port map( A1 => n4748, A2 => n2943, B1 => n3063, B2 => n2944
                           , ZN => n1801);
   U501 : OAI22_X1 port map( A1 => n5010, A2 => n2943, B1 => n3064, B2 => n2942
                           , ZN => n1800);
   U502 : CLKBUF_X1 port map( A => n2979, Z => n3065);
   U503 : OAI22_X1 port map( A1 => n5502, A2 => n2943, B1 => n3065, B2 => n2944
                           , ZN => n1799);
   U504 : CLKBUF_X1 port map( A => n2980, Z => n3066);
   U505 : OAI22_X1 port map( A1 => n4749, A2 => n2943, B1 => n3066, B2 => n2942
                           , ZN => n1798);
   U506 : CLKBUF_X1 port map( A => n2981, Z => n3067);
   U507 : OAI22_X1 port map( A1 => n5257, A2 => n2943, B1 => n3067, B2 => n2942
                           , ZN => n1797);
   U508 : CLKBUF_X1 port map( A => n2982, Z => n3068);
   U509 : OAI22_X1 port map( A1 => n4750, A2 => n2943, B1 => n3068, B2 => n2942
                           , ZN => n1796);
   U510 : CLKBUF_X1 port map( A => n2983, Z => n3069);
   U511 : OAI22_X1 port map( A1 => n5011, A2 => n2943, B1 => n3069, B2 => n2942
                           , ZN => n1795);
   U512 : CLKBUF_X1 port map( A => n2984, Z => n3070);
   U513 : OAI22_X1 port map( A1 => n5258, A2 => n2943, B1 => n3070, B2 => n2942
                           , ZN => n1794);
   U514 : CLKBUF_X1 port map( A => n2985, Z => n3071);
   U515 : OAI22_X1 port map( A1 => n4751, A2 => n2943, B1 => n3071, B2 => n2942
                           , ZN => n1793);
   U516 : CLKBUF_X1 port map( A => n2987, Z => n3073);
   U517 : OAI22_X1 port map( A1 => n4752, A2 => n2943, B1 => n3073, B2 => n2942
                           , ZN => n1792);
   U518 : CLKBUF_X1 port map( A => n2988, Z => n3074);
   U519 : OAI22_X1 port map( A1 => n4753, A2 => n2943, B1 => n3074, B2 => n2944
                           , ZN => n1791);
   U520 : CLKBUF_X1 port map( A => n2990, Z => n3075);
   U521 : OAI22_X1 port map( A1 => n5012, A2 => n2945, B1 => n3075, B2 => n2944
                           , ZN => n1790);
   U522 : CLKBUF_X1 port map( A => n2991, Z => n3076);
   U523 : OAI22_X1 port map( A1 => n5013, A2 => n2945, B1 => n3076, B2 => n2944
                           , ZN => n1789);
   U524 : CLKBUF_X1 port map( A => n2992, Z => n3077);
   U525 : OAI22_X1 port map( A1 => n4754, A2 => n2945, B1 => n3077, B2 => n2944
                           , ZN => n1788);
   U526 : CLKBUF_X1 port map( A => n2993, Z => n3078);
   U527 : OAI22_X1 port map( A1 => n5014, A2 => n2945, B1 => n3078, B2 => n2944
                           , ZN => n1787);
   U528 : CLKBUF_X1 port map( A => n2994, Z => n3079);
   U529 : OAI22_X1 port map( A1 => n5015, A2 => n2945, B1 => n3079, B2 => n2944
                           , ZN => n1786);
   U530 : OAI22_X1 port map( A1 => n4755, A2 => n2945, B1 => n3080, B2 => n2944
                           , ZN => n1785);
   U531 : CLKBUF_X1 port map( A => n2996, Z => n3081);
   U532 : OAI22_X1 port map( A1 => n4756, A2 => n2945, B1 => n3081, B2 => n2944
                           , ZN => n1784);
   U533 : CLKBUF_X1 port map( A => n2998, Z => n3083);
   U534 : OAI22_X1 port map( A1 => n5503, A2 => n2945, B1 => n3083, B2 => n2944
                           , ZN => n1783);
   U535 : NAND2_X1 port map( A1 => n3036, A2 => n2955, ZN => n2946);
   U536 : CLKBUF_X1 port map( A => n2946, Z => n2947);
   U537 : OAI22_X1 port map( A1 => n5504, A2 => n2948, B1 => n3014, B2 => n2947
                           , ZN => n1782);
   U538 : OAI22_X1 port map( A1 => n4757, A2 => n2948, B1 => n2965, B2 => n2946
                           , ZN => n1781);
   U539 : OAI22_X1 port map( A1 => n5505, A2 => n2948, B1 => n2966, B2 => n2947
                           , ZN => n1780);
   U540 : OAI22_X1 port map( A1 => n5259, A2 => n2948, B1 => n2967, B2 => n2946
                           , ZN => n1779);
   U541 : OAI22_X1 port map( A1 => n5260, A2 => n2948, B1 => n2968, B2 => n2947
                           , ZN => n1778);
   U542 : OAI22_X1 port map( A1 => n5506, A2 => n2948, B1 => n2969, B2 => n2946
                           , ZN => n1777);
   U543 : OAI22_X1 port map( A1 => n5261, A2 => n2948, B1 => n2970, B2 => n2947
                           , ZN => n1776);
   U544 : OAI22_X1 port map( A1 => n5507, A2 => n2948, B1 => n2971, B2 => n2946
                           , ZN => n1775);
   U545 : OAI22_X1 port map( A1 => n5262, A2 => n2948, B1 => n2972, B2 => n2947
                           , ZN => n1774);
   U546 : OAI22_X1 port map( A1 => n5016, A2 => n2948, B1 => n2973, B2 => n2946
                           , ZN => n1773);
   U547 : OAI22_X1 port map( A1 => n5263, A2 => n2948, B1 => n2974, B2 => n2946
                           , ZN => n1772);
   U548 : OAI22_X1 port map( A1 => n4758, A2 => n2948, B1 => n2975, B2 => n2947
                           , ZN => n1771);
   U549 : OAI22_X1 port map( A1 => n5017, A2 => n2948, B1 => n2976, B2 => n2946
                           , ZN => n1770);
   U550 : OAI22_X1 port map( A1 => n4759, A2 => n2948, B1 => n2977, B2 => n2947
                           , ZN => n1769);
   U551 : OAI22_X1 port map( A1 => n5018, A2 => n2948, B1 => n2978, B2 => n2946
                           , ZN => n1768);
   U552 : OAI22_X1 port map( A1 => n5508, A2 => n2948, B1 => n2979, B2 => n2947
                           , ZN => n1767);
   U553 : OAI22_X1 port map( A1 => n5264, A2 => n2948, B1 => n2980, B2 => n2946
                           , ZN => n1766);
   U554 : OAI22_X1 port map( A1 => n4760, A2 => n2948, B1 => n2981, B2 => n2946
                           , ZN => n1765);
   U555 : OAI22_X1 port map( A1 => n5265, A2 => n2948, B1 => n2982, B2 => n2946
                           , ZN => n1764);
   U556 : OAI22_X1 port map( A1 => n5266, A2 => n2948, B1 => n2983, B2 => n2946
                           , ZN => n1763);
   U557 : OAI22_X1 port map( A1 => n5267, A2 => n2948, B1 => n2984, B2 => n2946
                           , ZN => n1762);
   U558 : OAI22_X1 port map( A1 => n5019, A2 => n2948, B1 => n2985, B2 => n2946
                           , ZN => n1761);
   U559 : OAI22_X1 port map( A1 => n4761, A2 => n2948, B1 => n2987, B2 => n2946
                           , ZN => n1760);
   U560 : OAI22_X1 port map( A1 => n4762, A2 => n2948, B1 => n2988, B2 => n2947
                           , ZN => n1759);
   U561 : OAI22_X1 port map( A1 => n5509, A2 => n2948, B1 => n2990, B2 => n2947
                           , ZN => n1758);
   U562 : OAI22_X1 port map( A1 => n5268, A2 => n2948, B1 => n2991, B2 => n2947
                           , ZN => n1757);
   U563 : OAI22_X1 port map( A1 => n5020, A2 => n2948, B1 => n2992, B2 => n2947
                           , ZN => n1756);
   U564 : OAI22_X1 port map( A1 => n5510, A2 => n2948, B1 => n2993, B2 => n2947
                           , ZN => n1755);
   U565 : OAI22_X1 port map( A1 => n5511, A2 => n2948, B1 => n2994, B2 => n2947
                           , ZN => n1754);
   U566 : OAI22_X1 port map( A1 => n4763, A2 => n2948, B1 => n2995, B2 => n2947
                           , ZN => n1753);
   U567 : OAI22_X1 port map( A1 => n5512, A2 => n2948, B1 => n2996, B2 => n2947
                           , ZN => n1752);
   U568 : OAI22_X1 port map( A1 => n5513, A2 => n2948, B1 => n2998, B2 => n2947
                           , ZN => n1751);
   U569 : NAND2_X1 port map( A1 => n3040, A2 => n2955, ZN => n2949);
   U570 : CLKBUF_X1 port map( A => n2949, Z => n2950);
   U571 : OAI22_X1 port map( A1 => n5514, A2 => n2951, B1 => n3014, B2 => n2950
                           , ZN => n1750);
   U572 : OAI22_X1 port map( A1 => n5269, A2 => n2951, B1 => n3051, B2 => n2949
                           , ZN => n1749);
   U573 : OAI22_X1 port map( A1 => n5270, A2 => n2951, B1 => n3052, B2 => n2950
                           , ZN => n1748);
   U574 : OAI22_X1 port map( A1 => n5515, A2 => n2951, B1 => n3053, B2 => n2949
                           , ZN => n1747);
   U575 : OAI22_X1 port map( A1 => n5271, A2 => n2951, B1 => n3054, B2 => n2950
                           , ZN => n1746);
   U576 : OAI22_X1 port map( A1 => n5516, A2 => n2951, B1 => n3055, B2 => n2949
                           , ZN => n1745);
   U577 : OAI22_X1 port map( A1 => n5272, A2 => n2951, B1 => n3056, B2 => n2950
                           , ZN => n1744);
   U578 : OAI22_X1 port map( A1 => n5273, A2 => n2951, B1 => n3057, B2 => n2949
                           , ZN => n1743);
   U579 : OAI22_X1 port map( A1 => n5517, A2 => n2951, B1 => n3058, B2 => n2950
                           , ZN => n1742);
   U580 : OAI22_X1 port map( A1 => n5518, A2 => n2951, B1 => n3059, B2 => n2949
                           , ZN => n1741);
   U581 : OAI22_X1 port map( A1 => n5274, A2 => n2951, B1 => n3060, B2 => n2949
                           , ZN => n1740);
   U582 : OAI22_X1 port map( A1 => n5275, A2 => n2951, B1 => n3061, B2 => n2950
                           , ZN => n1739);
   U583 : OAI22_X1 port map( A1 => n5276, A2 => n2951, B1 => n3062, B2 => n2949
                           , ZN => n1738);
   U584 : OAI22_X1 port map( A1 => n5519, A2 => n2951, B1 => n3063, B2 => n2950
                           , ZN => n1737);
   U585 : OAI22_X1 port map( A1 => n5520, A2 => n2951, B1 => n3064, B2 => n2949
                           , ZN => n1736);
   U586 : OAI22_X1 port map( A1 => n5277, A2 => n2951, B1 => n3065, B2 => n2950
                           , ZN => n1735);
   U587 : OAI22_X1 port map( A1 => n5521, A2 => n2951, B1 => n3066, B2 => n2949
                           , ZN => n1734);
   U588 : OAI22_X1 port map( A1 => n5522, A2 => n2951, B1 => n3067, B2 => n2949
                           , ZN => n1733);
   U589 : OAI22_X1 port map( A1 => n5523, A2 => n2951, B1 => n3068, B2 => n2949
                           , ZN => n1732);
   U590 : OAI22_X1 port map( A1 => n5278, A2 => n2951, B1 => n3069, B2 => n2949
                           , ZN => n1731);
   U591 : OAI22_X1 port map( A1 => n5524, A2 => n2951, B1 => n3070, B2 => n2949
                           , ZN => n1730);
   U592 : OAI22_X1 port map( A1 => n5279, A2 => n2951, B1 => n3071, B2 => n2949
                           , ZN => n1729);
   U593 : OAI22_X1 port map( A1 => n5525, A2 => n2951, B1 => n3073, B2 => n2949
                           , ZN => n1728);
   U594 : OAI22_X1 port map( A1 => n5526, A2 => n2951, B1 => n3074, B2 => n2950
                           , ZN => n1727);
   U595 : OAI22_X1 port map( A1 => n5280, A2 => n2951, B1 => n3075, B2 => n2950
                           , ZN => n1726);
   U596 : OAI22_X1 port map( A1 => n5527, A2 => n2951, B1 => n3076, B2 => n2950
                           , ZN => n1725);
   U597 : OAI22_X1 port map( A1 => n5528, A2 => n2951, B1 => n3077, B2 => n2950
                           , ZN => n1724);
   U598 : OAI22_X1 port map( A1 => n5281, A2 => n2951, B1 => n3078, B2 => n2950
                           , ZN => n1723);
   U599 : OAI22_X1 port map( A1 => n5021, A2 => n2951, B1 => n3079, B2 => n2950
                           , ZN => n1722);
   U600 : OAI22_X1 port map( A1 => n5282, A2 => n2951, B1 => n3080, B2 => n2950
                           , ZN => n1721);
   U601 : OAI22_X1 port map( A1 => n5529, A2 => n2951, B1 => n3081, B2 => n2950
                           , ZN => n1720);
   U602 : OAI22_X1 port map( A1 => n5022, A2 => n2951, B1 => n3083, B2 => n2950
                           , ZN => n1719);
   U603 : NAND2_X1 port map( A1 => n3044, A2 => n2955, ZN => n2952);
   U604 : CLKBUF_X1 port map( A => n2952, Z => n2953);
   U605 : OAI22_X1 port map( A1 => n4764, A2 => n2954, B1 => n3014, B2 => n2953
                           , ZN => n1718);
   U606 : OAI22_X1 port map( A1 => n5530, A2 => n2954, B1 => n2965, B2 => n2952
                           , ZN => n1717);
   U607 : OAI22_X1 port map( A1 => n5531, A2 => n2954, B1 => n2966, B2 => n2953
                           , ZN => n1716);
   U608 : OAI22_X1 port map( A1 => n5283, A2 => n2954, B1 => n2967, B2 => n2952
                           , ZN => n1715);
   U609 : OAI22_X1 port map( A1 => n5023, A2 => n2954, B1 => n2968, B2 => n2953
                           , ZN => n1714);
   U610 : OAI22_X1 port map( A1 => n4765, A2 => n2954, B1 => n2969, B2 => n2952
                           , ZN => n1713);
   U611 : OAI22_X1 port map( A1 => n5532, A2 => n2954, B1 => n2970, B2 => n2953
                           , ZN => n1712);
   U612 : OAI22_X1 port map( A1 => n5284, A2 => n2954, B1 => n2971, B2 => n2952
                           , ZN => n1711);
   U613 : OAI22_X1 port map( A1 => n5024, A2 => n2954, B1 => n2972, B2 => n2953
                           , ZN => n1710);
   U614 : OAI22_X1 port map( A1 => n4766, A2 => n2954, B1 => n2973, B2 => n2952
                           , ZN => n1709);
   U615 : OAI22_X1 port map( A1 => n5025, A2 => n2954, B1 => n2974, B2 => n2952
                           , ZN => n1708);
   U616 : OAI22_X1 port map( A1 => n5285, A2 => n2954, B1 => n2975, B2 => n2953
                           , ZN => n1707);
   U617 : OAI22_X1 port map( A1 => n5533, A2 => n2954, B1 => n2976, B2 => n2952
                           , ZN => n1706);
   U618 : OAI22_X1 port map( A1 => n5534, A2 => n2954, B1 => n2977, B2 => n2953
                           , ZN => n1705);
   U619 : OAI22_X1 port map( A1 => n5286, A2 => n2954, B1 => n2978, B2 => n2952
                           , ZN => n1704);
   U620 : OAI22_X1 port map( A1 => n5026, A2 => n2954, B1 => n2979, B2 => n2953
                           , ZN => n1703);
   U621 : OAI22_X1 port map( A1 => n5287, A2 => n2954, B1 => n2980, B2 => n2952
                           , ZN => n1702);
   U622 : OAI22_X1 port map( A1 => n5535, A2 => n2954, B1 => n2981, B2 => n2952
                           , ZN => n1701);
   U623 : OAI22_X1 port map( A1 => n5027, A2 => n2954, B1 => n2982, B2 => n2952
                           , ZN => n1700);
   U624 : OAI22_X1 port map( A1 => n5536, A2 => n2954, B1 => n2983, B2 => n2952
                           , ZN => n1699);
   U625 : OAI22_X1 port map( A1 => n5028, A2 => n2954, B1 => n2984, B2 => n2952
                           , ZN => n1698);
   U626 : OAI22_X1 port map( A1 => n5537, A2 => n2954, B1 => n2985, B2 => n2952
                           , ZN => n1697);
   U627 : OAI22_X1 port map( A1 => n5288, A2 => n2954, B1 => n2987, B2 => n2952
                           , ZN => n1696);
   U628 : OAI22_X1 port map( A1 => n5538, A2 => n2954, B1 => n2988, B2 => n2953
                           , ZN => n1695);
   U629 : OAI22_X1 port map( A1 => n4767, A2 => n2954, B1 => n2990, B2 => n2953
                           , ZN => n1694);
   U630 : OAI22_X1 port map( A1 => n4768, A2 => n2954, B1 => n2991, B2 => n2953
                           , ZN => n1693);
   U631 : OAI22_X1 port map( A1 => n5289, A2 => n2954, B1 => n2992, B2 => n2953
                           , ZN => n1692);
   U632 : OAI22_X1 port map( A1 => n4769, A2 => n2954, B1 => n2993, B2 => n2953
                           , ZN => n1691);
   U633 : OAI22_X1 port map( A1 => n5290, A2 => n2954, B1 => n2994, B2 => n2953
                           , ZN => n1690);
   U634 : OAI22_X1 port map( A1 => n5539, A2 => n2954, B1 => n2995, B2 => n2953
                           , ZN => n1689);
   U635 : OAI22_X1 port map( A1 => n4770, A2 => n2954, B1 => n2996, B2 => n2953
                           , ZN => n1688);
   U636 : OAI22_X1 port map( A1 => n5291, A2 => n2954, B1 => n2998, B2 => n2953
                           , ZN => n1687);
   U637 : NAND2_X1 port map( A1 => n3049, A2 => n2955, ZN => n2956);
   U638 : CLKBUF_X1 port map( A => n2956, Z => n2957);
   U639 : OAI22_X1 port map( A1 => n5029, A2 => n2958, B1 => n3014, B2 => n2957
                           , ZN => n1686);
   U640 : OAI22_X1 port map( A1 => n4771, A2 => n2958, B1 => n3051, B2 => n2956
                           , ZN => n1685);
   U641 : OAI22_X1 port map( A1 => n5030, A2 => n2958, B1 => n3052, B2 => n2957
                           , ZN => n1684);
   U642 : OAI22_X1 port map( A1 => n5031, A2 => n2958, B1 => n3053, B2 => n2956
                           , ZN => n1683);
   U643 : OAI22_X1 port map( A1 => n4772, A2 => n2958, B1 => n3054, B2 => n2957
                           , ZN => n1682);
   U644 : OAI22_X1 port map( A1 => n5032, A2 => n2958, B1 => n3055, B2 => n2956
                           , ZN => n1681);
   U645 : OAI22_X1 port map( A1 => n5033, A2 => n2958, B1 => n3056, B2 => n2957
                           , ZN => n1680);
   U646 : OAI22_X1 port map( A1 => n4773, A2 => n2958, B1 => n3057, B2 => n2956
                           , ZN => n1679);
   U647 : OAI22_X1 port map( A1 => n4774, A2 => n2958, B1 => n3058, B2 => n2957
                           , ZN => n1678);
   U648 : OAI22_X1 port map( A1 => n5034, A2 => n2958, B1 => n3059, B2 => n2956
                           , ZN => n1677);
   U649 : OAI22_X1 port map( A1 => n4775, A2 => n2958, B1 => n3060, B2 => n2956
                           , ZN => n1676);
   U650 : OAI22_X1 port map( A1 => n5035, A2 => n2958, B1 => n3061, B2 => n2957
                           , ZN => n1675);
   U651 : OAI22_X1 port map( A1 => n5036, A2 => n2958, B1 => n3062, B2 => n2956
                           , ZN => n1674);
   U652 : OAI22_X1 port map( A1 => n5037, A2 => n2958, B1 => n3063, B2 => n2957
                           , ZN => n1673);
   U653 : OAI22_X1 port map( A1 => n4776, A2 => n2958, B1 => n3064, B2 => n2956
                           , ZN => n1672);
   U654 : OAI22_X1 port map( A1 => n4777, A2 => n2958, B1 => n3065, B2 => n2957
                           , ZN => n1671);
   U655 : OAI22_X1 port map( A1 => n5038, A2 => n2958, B1 => n3066, B2 => n2956
                           , ZN => n1670);
   U656 : OAI22_X1 port map( A1 => n4778, A2 => n2958, B1 => n3067, B2 => n2956
                           , ZN => n1669);
   U657 : OAI22_X1 port map( A1 => n5039, A2 => n2958, B1 => n3068, B2 => n2956
                           , ZN => n1668);
   U658 : OAI22_X1 port map( A1 => n4779, A2 => n2958, B1 => n3069, B2 => n2956
                           , ZN => n1667);
   U659 : OAI22_X1 port map( A1 => n5040, A2 => n2958, B1 => n3070, B2 => n2956
                           , ZN => n1666);
   U660 : OAI22_X1 port map( A1 => n4780, A2 => n2958, B1 => n3071, B2 => n2956
                           , ZN => n1665);
   U661 : OAI22_X1 port map( A1 => n5041, A2 => n2958, B1 => n3073, B2 => n2956
                           , ZN => n1664);
   U662 : OAI22_X1 port map( A1 => n5042, A2 => n2958, B1 => n3074, B2 => n2957
                           , ZN => n1663);
   U663 : OAI22_X1 port map( A1 => n4781, A2 => n2958, B1 => n3075, B2 => n2957
                           , ZN => n1662);
   U664 : OAI22_X1 port map( A1 => n5043, A2 => n2958, B1 => n3076, B2 => n2957
                           , ZN => n1661);
   U665 : OAI22_X1 port map( A1 => n5044, A2 => n2958, B1 => n3077, B2 => n2957
                           , ZN => n1660);
   U666 : OAI22_X1 port map( A1 => n5045, A2 => n2958, B1 => n3078, B2 => n2957
                           , ZN => n1659);
   U667 : OAI22_X1 port map( A1 => n4782, A2 => n2958, B1 => n3079, B2 => n2957
                           , ZN => n1658);
   U668 : OAI22_X1 port map( A1 => n5046, A2 => n2958, B1 => n3080, B2 => n2957
                           , ZN => n1657);
   U669 : OAI22_X1 port map( A1 => n5047, A2 => n2958, B1 => n3081, B2 => n2957
                           , ZN => n1656);
   U670 : OAI22_X1 port map( A1 => n4783, A2 => n2958, B1 => n3083, B2 => n2957
                           , ZN => n1655);
   U671 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => ADD_WR(4), ZN => 
                           n3018);
   U672 : NOR2_X1 port map( A1 => ADD_WR(3), A2 => n3018, ZN => n3013);
   U673 : NAND2_X1 port map( A1 => n3020, A2 => n3013, ZN => n2959);
   U674 : CLKBUF_X1 port map( A => n2959, Z => n2960);
   U675 : OAI22_X1 port map( A1 => n5164, A2 => n2961, B1 => n3014, B2 => n2960
                           , ZN => n1654);
   U676 : OAI22_X1 port map( A1 => n5292, A2 => n2961, B1 => n2965, B2 => n2959
                           , ZN => n1653);
   U677 : OAI22_X1 port map( A1 => n5293, A2 => n2961, B1 => n2966, B2 => n2960
                           , ZN => n1652);
   U678 : OAI22_X1 port map( A1 => n5540, A2 => n2961, B1 => n2967, B2 => n2959
                           , ZN => n1651);
   U679 : OAI22_X1 port map( A1 => n5294, A2 => n2961, B1 => n2968, B2 => n2960
                           , ZN => n1650);
   U680 : OAI22_X1 port map( A1 => n5295, A2 => n2961, B1 => n2969, B2 => n2959
                           , ZN => n1649);
   U681 : OAI22_X1 port map( A1 => n5296, A2 => n2961, B1 => n2970, B2 => n2960
                           , ZN => n1648);
   U682 : OAI22_X1 port map( A1 => n5541, A2 => n2961, B1 => n2971, B2 => n2959
                           , ZN => n1647);
   U683 : OAI22_X1 port map( A1 => n4784, A2 => n2961, B1 => n2972, B2 => n2960
                           , ZN => n1646);
   U684 : OAI22_X1 port map( A1 => n5542, A2 => n2961, B1 => n2973, B2 => n2959
                           , ZN => n1645);
   U685 : OAI22_X1 port map( A1 => n5297, A2 => n2961, B1 => n2974, B2 => n2959
                           , ZN => n1644);
   U686 : OAI22_X1 port map( A1 => n5298, A2 => n2961, B1 => n2975, B2 => n2960
                           , ZN => n1643);
   U687 : OAI22_X1 port map( A1 => n4785, A2 => n2961, B1 => n2976, B2 => n2959
                           , ZN => n1642);
   U688 : OAI22_X1 port map( A1 => n5543, A2 => n2961, B1 => n2977, B2 => n2960
                           , ZN => n1641);
   U689 : OAI22_X1 port map( A1 => n5299, A2 => n2961, B1 => n2978, B2 => n2959
                           , ZN => n1640);
   U690 : OAI22_X1 port map( A1 => n5544, A2 => n2961, B1 => n2979, B2 => n2960
                           , ZN => n1639);
   U691 : OAI22_X1 port map( A1 => n5545, A2 => n2961, B1 => n2980, B2 => n2959
                           , ZN => n1638);
   U692 : OAI22_X1 port map( A1 => n5300, A2 => n2961, B1 => n2981, B2 => n2959
                           , ZN => n1637);
   U693 : OAI22_X1 port map( A1 => n5546, A2 => n2961, B1 => n2982, B2 => n2959
                           , ZN => n1636);
   U694 : OAI22_X1 port map( A1 => n5301, A2 => n2961, B1 => n2983, B2 => n2959
                           , ZN => n1635);
   U695 : OAI22_X1 port map( A1 => n5547, A2 => n2961, B1 => n2984, B2 => n2959
                           , ZN => n1634);
   U696 : OAI22_X1 port map( A1 => n4786, A2 => n2961, B1 => n2985, B2 => n2959
                           , ZN => n1633);
   U697 : OAI22_X1 port map( A1 => n5548, A2 => n2961, B1 => n2987, B2 => n2959
                           , ZN => n1632);
   U698 : OAI22_X1 port map( A1 => n5549, A2 => n2961, B1 => n2988, B2 => n2960
                           , ZN => n1631);
   U699 : OAI22_X1 port map( A1 => n5550, A2 => n2961, B1 => n2990, B2 => n2960
                           , ZN => n1630);
   U700 : OAI22_X1 port map( A1 => n5302, A2 => n2961, B1 => n2991, B2 => n2960
                           , ZN => n1629);
   U701 : OAI22_X1 port map( A1 => n5303, A2 => n2961, B1 => n2992, B2 => n2960
                           , ZN => n1628);
   U702 : OAI22_X1 port map( A1 => n5551, A2 => n2961, B1 => n2993, B2 => n2960
                           , ZN => n1627);
   U703 : OAI22_X1 port map( A1 => n5304, A2 => n2961, B1 => n2994, B2 => n2960
                           , ZN => n1626);
   U704 : OAI22_X1 port map( A1 => n5552, A2 => n2961, B1 => n2995, B2 => n2960
                           , ZN => n1625);
   U705 : OAI22_X1 port map( A1 => n4787, A2 => n2961, B1 => n2996, B2 => n2960
                           , ZN => n1624);
   U706 : OAI22_X1 port map( A1 => n5048, A2 => n2961, B1 => n2998, B2 => n2960
                           , ZN => n1623);
   U707 : NAND2_X1 port map( A1 => n3024, A2 => n3013, ZN => n2962);
   U708 : CLKBUF_X1 port map( A => n2962, Z => n2963);
   U709 : OAI22_X1 port map( A1 => n4916, A2 => n2964, B1 => n3014, B2 => n2963
                           , ZN => n1622);
   U710 : OAI22_X1 port map( A1 => n5553, A2 => n2964, B1 => n3051, B2 => n2962
                           , ZN => n1621);
   U711 : OAI22_X1 port map( A1 => n5305, A2 => n2964, B1 => n3052, B2 => n2963
                           , ZN => n1620);
   U712 : OAI22_X1 port map( A1 => n5049, A2 => n2964, B1 => n3053, B2 => n2962
                           , ZN => n1619);
   U713 : OAI22_X1 port map( A1 => n4788, A2 => n2964, B1 => n3054, B2 => n2963
                           , ZN => n1618);
   U714 : OAI22_X1 port map( A1 => n5554, A2 => n2964, B1 => n3055, B2 => n2962
                           , ZN => n1617);
   U715 : OAI22_X1 port map( A1 => n5555, A2 => n2964, B1 => n3056, B2 => n2963
                           , ZN => n1616);
   U716 : OAI22_X1 port map( A1 => n5306, A2 => n2964, B1 => n3057, B2 => n2962
                           , ZN => n1615);
   U717 : OAI22_X1 port map( A1 => n5556, A2 => n2964, B1 => n3058, B2 => n2963
                           , ZN => n1614);
   U718 : OAI22_X1 port map( A1 => n4789, A2 => n2964, B1 => n3059, B2 => n2962
                           , ZN => n1613);
   U719 : OAI22_X1 port map( A1 => n4790, A2 => n2964, B1 => n3060, B2 => n2962
                           , ZN => n1612);
   U720 : OAI22_X1 port map( A1 => n4791, A2 => n2964, B1 => n3061, B2 => n2963
                           , ZN => n1611);
   U721 : OAI22_X1 port map( A1 => n5050, A2 => n2964, B1 => n3062, B2 => n2962
                           , ZN => n1610);
   U722 : OAI22_X1 port map( A1 => n5051, A2 => n2964, B1 => n3063, B2 => n2963
                           , ZN => n1609);
   U723 : OAI22_X1 port map( A1 => n5307, A2 => n2964, B1 => n3064, B2 => n2962
                           , ZN => n1608);
   U724 : OAI22_X1 port map( A1 => n5557, A2 => n2964, B1 => n3065, B2 => n2963
                           , ZN => n1607);
   U725 : OAI22_X1 port map( A1 => n5308, A2 => n2964, B1 => n3066, B2 => n2962
                           , ZN => n1606);
   U726 : OAI22_X1 port map( A1 => n5558, A2 => n2964, B1 => n3067, B2 => n2962
                           , ZN => n1605);
   U727 : OAI22_X1 port map( A1 => n4792, A2 => n2964, B1 => n3068, B2 => n2962
                           , ZN => n1604);
   U728 : OAI22_X1 port map( A1 => n5309, A2 => n2964, B1 => n3069, B2 => n2962
                           , ZN => n1603);
   U729 : OAI22_X1 port map( A1 => n5310, A2 => n2964, B1 => n3070, B2 => n2962
                           , ZN => n1602);
   U730 : OAI22_X1 port map( A1 => n5052, A2 => n2964, B1 => n3071, B2 => n2962
                           , ZN => n1601);
   U731 : OAI22_X1 port map( A1 => n5311, A2 => n2964, B1 => n3073, B2 => n2962
                           , ZN => n1600);
   U732 : OAI22_X1 port map( A1 => n4793, A2 => n2964, B1 => n3074, B2 => n2963
                           , ZN => n1599);
   U733 : OAI22_X1 port map( A1 => n5559, A2 => n2964, B1 => n3075, B2 => n2963
                           , ZN => n1598);
   U734 : OAI22_X1 port map( A1 => n5560, A2 => n2964, B1 => n3076, B2 => n2963
                           , ZN => n1597);
   U735 : OAI22_X1 port map( A1 => n5312, A2 => n2964, B1 => n3077, B2 => n2963
                           , ZN => n1596);
   U736 : OAI22_X1 port map( A1 => n5561, A2 => n2964, B1 => n3078, B2 => n2963
                           , ZN => n1595);
   U737 : OAI22_X1 port map( A1 => n4794, A2 => n2964, B1 => n3079, B2 => n2963
                           , ZN => n1594);
   U738 : OAI22_X1 port map( A1 => n5562, A2 => n2964, B1 => n3080, B2 => n2963
                           , ZN => n1593);
   U739 : OAI22_X1 port map( A1 => n4795, A2 => n2964, B1 => n3081, B2 => n2963
                           , ZN => n1592);
   U740 : OAI22_X1 port map( A1 => n4796, A2 => n2964, B1 => n3083, B2 => n2963
                           , ZN => n1591);
   U741 : NAND2_X1 port map( A1 => n3028, A2 => n3013, ZN => n2986);
   U742 : CLKBUF_X1 port map( A => n2999, Z => n2989);
   U743 : CLKBUF_X1 port map( A => n2986, Z => n2997);
   U744 : OAI22_X1 port map( A1 => n4917, A2 => n2989, B1 => n3014, B2 => n2997
                           , ZN => n1590);
   U745 : OAI22_X1 port map( A1 => n5053, A2 => n2999, B1 => n2965, B2 => n2986
                           , ZN => n1589);
   U746 : OAI22_X1 port map( A1 => n5054, A2 => n2989, B1 => n2966, B2 => n2997
                           , ZN => n1588);
   U747 : OAI22_X1 port map( A1 => n5055, A2 => n2999, B1 => n2967, B2 => n2986
                           , ZN => n1587);
   U748 : OAI22_X1 port map( A1 => n5056, A2 => n2989, B1 => n2968, B2 => n2997
                           , ZN => n1586);
   U749 : OAI22_X1 port map( A1 => n4797, A2 => n2999, B1 => n2969, B2 => n2986
                           , ZN => n1585);
   U750 : OAI22_X1 port map( A1 => n5057, A2 => n2989, B1 => n2970, B2 => n2997
                           , ZN => n1584);
   U751 : OAI22_X1 port map( A1 => n5058, A2 => n2999, B1 => n2971, B2 => n2986
                           , ZN => n1583);
   U752 : OAI22_X1 port map( A1 => n5059, A2 => n2989, B1 => n2972, B2 => n2997
                           , ZN => n1582);
   U753 : OAI22_X1 port map( A1 => n4798, A2 => n2999, B1 => n2973, B2 => n2986
                           , ZN => n1581);
   U754 : OAI22_X1 port map( A1 => n4799, A2 => n2999, B1 => n2974, B2 => n2986
                           , ZN => n1580);
   U755 : OAI22_X1 port map( A1 => n5060, A2 => n2999, B1 => n2975, B2 => n2997
                           , ZN => n1579);
   U756 : OAI22_X1 port map( A1 => n4800, A2 => n2989, B1 => n2976, B2 => n2986
                           , ZN => n1578);
   U757 : OAI22_X1 port map( A1 => n4801, A2 => n2989, B1 => n2977, B2 => n2997
                           , ZN => n1577);
   U758 : OAI22_X1 port map( A1 => n5061, A2 => n2989, B1 => n2978, B2 => n2986
                           , ZN => n1576);
   U759 : OAI22_X1 port map( A1 => n5062, A2 => n2989, B1 => n2979, B2 => n2997
                           , ZN => n1575);
   U760 : OAI22_X1 port map( A1 => n5063, A2 => n2989, B1 => n2980, B2 => n2986
                           , ZN => n1574);
   U761 : OAI22_X1 port map( A1 => n5313, A2 => n2989, B1 => n2981, B2 => n2986
                           , ZN => n1573);
   U762 : OAI22_X1 port map( A1 => n5064, A2 => n2989, B1 => n2982, B2 => n2986
                           , ZN => n1572);
   U763 : OAI22_X1 port map( A1 => n4802, A2 => n2989, B1 => n2983, B2 => n2986
                           , ZN => n1571);
   U764 : OAI22_X1 port map( A1 => n5065, A2 => n2989, B1 => n2984, B2 => n2986
                           , ZN => n1570);
   U765 : OAI22_X1 port map( A1 => n4803, A2 => n2989, B1 => n2985, B2 => n2986
                           , ZN => n1569);
   U766 : OAI22_X1 port map( A1 => n5066, A2 => n2989, B1 => n2987, B2 => n2986
                           , ZN => n1568);
   U767 : OAI22_X1 port map( A1 => n4804, A2 => n2989, B1 => n2988, B2 => n2997
                           , ZN => n1567);
   U768 : OAI22_X1 port map( A1 => n4805, A2 => n2999, B1 => n2990, B2 => n2997
                           , ZN => n1566);
   U769 : OAI22_X1 port map( A1 => n5067, A2 => n2999, B1 => n2991, B2 => n2997
                           , ZN => n1565);
   U770 : OAI22_X1 port map( A1 => n5068, A2 => n2999, B1 => n2992, B2 => n2997
                           , ZN => n1564);
   U771 : OAI22_X1 port map( A1 => n4806, A2 => n2999, B1 => n2993, B2 => n2997
                           , ZN => n1563);
   U772 : OAI22_X1 port map( A1 => n5069, A2 => n2999, B1 => n2994, B2 => n2997
                           , ZN => n1562);
   U773 : OAI22_X1 port map( A1 => n4807, A2 => n2999, B1 => n2995, B2 => n2997
                           , ZN => n1561);
   U774 : OAI22_X1 port map( A1 => n5070, A2 => n2999, B1 => n2996, B2 => n2997
                           , ZN => n1560);
   U775 : OAI22_X1 port map( A1 => n5071, A2 => n2999, B1 => n2998, B2 => n2997
                           , ZN => n1559);
   U776 : NAND2_X1 port map( A1 => n3032, A2 => n3013, ZN => n3000);
   U777 : CLKBUF_X1 port map( A => n3000, Z => n3001);
   U778 : OAI22_X1 port map( A1 => n4918, A2 => n3002, B1 => n3014, B2 => n3001
                           , ZN => n1558);
   U779 : OAI22_X1 port map( A1 => n4808, A2 => n3002, B1 => n3051, B2 => n3000
                           , ZN => n1557);
   U780 : OAI22_X1 port map( A1 => n5563, A2 => n3002, B1 => n3052, B2 => n3001
                           , ZN => n1556);
   U781 : OAI22_X1 port map( A1 => n4809, A2 => n3002, B1 => n3053, B2 => n3000
                           , ZN => n1555);
   U782 : OAI22_X1 port map( A1 => n4810, A2 => n3002, B1 => n3054, B2 => n3001
                           , ZN => n1554);
   U783 : OAI22_X1 port map( A1 => n5564, A2 => n3002, B1 => n3055, B2 => n3000
                           , ZN => n1553);
   U784 : OAI22_X1 port map( A1 => n5072, A2 => n3002, B1 => n3056, B2 => n3001
                           , ZN => n1552);
   U785 : OAI22_X1 port map( A1 => n4811, A2 => n3002, B1 => n3057, B2 => n3000
                           , ZN => n1551);
   U786 : OAI22_X1 port map( A1 => n5073, A2 => n3002, B1 => n3058, B2 => n3001
                           , ZN => n1550);
   U787 : OAI22_X1 port map( A1 => n5074, A2 => n3002, B1 => n3059, B2 => n3000
                           , ZN => n1549);
   U788 : OAI22_X1 port map( A1 => n5075, A2 => n3002, B1 => n3060, B2 => n3000
                           , ZN => n1548);
   U789 : OAI22_X1 port map( A1 => n5565, A2 => n3002, B1 => n3061, B2 => n3001
                           , ZN => n1547);
   U790 : OAI22_X1 port map( A1 => n5076, A2 => n3002, B1 => n3062, B2 => n3000
                           , ZN => n1546);
   U791 : OAI22_X1 port map( A1 => n5566, A2 => n3002, B1 => n3063, B2 => n3001
                           , ZN => n1545);
   U792 : OAI22_X1 port map( A1 => n5314, A2 => n3002, B1 => n3064, B2 => n3000
                           , ZN => n1544);
   U793 : OAI22_X1 port map( A1 => n5567, A2 => n3002, B1 => n3065, B2 => n3001
                           , ZN => n1543);
   U794 : OAI22_X1 port map( A1 => n5077, A2 => n3002, B1 => n3066, B2 => n3000
                           , ZN => n1542);
   U795 : OAI22_X1 port map( A1 => n5078, A2 => n3002, B1 => n3067, B2 => n3000
                           , ZN => n1541);
   U796 : OAI22_X1 port map( A1 => n4812, A2 => n3002, B1 => n3068, B2 => n3000
                           , ZN => n1540);
   U797 : OAI22_X1 port map( A1 => n5079, A2 => n3002, B1 => n3069, B2 => n3000
                           , ZN => n1539);
   U798 : OAI22_X1 port map( A1 => n5080, A2 => n3002, B1 => n3070, B2 => n3000
                           , ZN => n1538);
   U799 : OAI22_X1 port map( A1 => n5568, A2 => n3002, B1 => n3071, B2 => n3000
                           , ZN => n1537);
   U800 : OAI22_X1 port map( A1 => n4813, A2 => n3002, B1 => n3073, B2 => n3000
                           , ZN => n1536);
   U801 : OAI22_X1 port map( A1 => n4814, A2 => n3002, B1 => n3074, B2 => n3001
                           , ZN => n1535);
   U802 : OAI22_X1 port map( A1 => n4815, A2 => n3002, B1 => n3075, B2 => n3001
                           , ZN => n1534);
   U803 : OAI22_X1 port map( A1 => n4816, A2 => n3002, B1 => n3076, B2 => n3001
                           , ZN => n1533);
   U804 : OAI22_X1 port map( A1 => n5315, A2 => n3002, B1 => n3077, B2 => n3001
                           , ZN => n1532);
   U805 : OAI22_X1 port map( A1 => n4817, A2 => n3002, B1 => n3078, B2 => n3001
                           , ZN => n1531);
   U806 : OAI22_X1 port map( A1 => n5316, A2 => n3002, B1 => n3079, B2 => n3001
                           , ZN => n1530);
   U807 : OAI22_X1 port map( A1 => n4818, A2 => n3002, B1 => n3080, B2 => n3001
                           , ZN => n1529);
   U808 : OAI22_X1 port map( A1 => n5569, A2 => n3002, B1 => n3081, B2 => n3001
                           , ZN => n1528);
   U809 : OAI22_X1 port map( A1 => n5570, A2 => n3002, B1 => n3083, B2 => n3001
                           , ZN => n1527);
   U810 : NAND2_X1 port map( A1 => n3036, A2 => n3013, ZN => n3003);
   U811 : CLKBUF_X1 port map( A => n3003, Z => n3004);
   U812 : OAI22_X1 port map( A1 => n4919, A2 => n3005, B1 => n3014, B2 => n3004
                           , ZN => n1526);
   U813 : OAI22_X1 port map( A1 => n4819, A2 => n3005, B1 => n3051, B2 => n3003
                           , ZN => n1525);
   U814 : OAI22_X1 port map( A1 => n4820, A2 => n3005, B1 => n3052, B2 => n3004
                           , ZN => n1524);
   U815 : OAI22_X1 port map( A1 => n5571, A2 => n3005, B1 => n3053, B2 => n3003
                           , ZN => n1523);
   U816 : OAI22_X1 port map( A1 => n5317, A2 => n3005, B1 => n3054, B2 => n3004
                           , ZN => n1522);
   U817 : OAI22_X1 port map( A1 => n4821, A2 => n3005, B1 => n3055, B2 => n3003
                           , ZN => n1521);
   U818 : OAI22_X1 port map( A1 => n4822, A2 => n3005, B1 => n3056, B2 => n3004
                           , ZN => n1520);
   U819 : OAI22_X1 port map( A1 => n5081, A2 => n3005, B1 => n3057, B2 => n3003
                           , ZN => n1519);
   U820 : OAI22_X1 port map( A1 => n5572, A2 => n3005, B1 => n3058, B2 => n3004
                           , ZN => n1518);
   U821 : OAI22_X1 port map( A1 => n5573, A2 => n3005, B1 => n3059, B2 => n3003
                           , ZN => n1517);
   U822 : OAI22_X1 port map( A1 => n4823, A2 => n3005, B1 => n3060, B2 => n3003
                           , ZN => n1516);
   U823 : OAI22_X1 port map( A1 => n5082, A2 => n3005, B1 => n3061, B2 => n3004
                           , ZN => n1515);
   U824 : OAI22_X1 port map( A1 => n4824, A2 => n3005, B1 => n3062, B2 => n3003
                           , ZN => n1514);
   U825 : OAI22_X1 port map( A1 => n5318, A2 => n3005, B1 => n3063, B2 => n3004
                           , ZN => n1513);
   U826 : OAI22_X1 port map( A1 => n5083, A2 => n3005, B1 => n3064, B2 => n3003
                           , ZN => n1512);
   U827 : OAI22_X1 port map( A1 => n4825, A2 => n3005, B1 => n3065, B2 => n3004
                           , ZN => n1511);
   U828 : OAI22_X1 port map( A1 => n5574, A2 => n3005, B1 => n3066, B2 => n3003
                           , ZN => n1510);
   U829 : OAI22_X1 port map( A1 => n5084, A2 => n3005, B1 => n3067, B2 => n3003
                           , ZN => n1509);
   U830 : OAI22_X1 port map( A1 => n4826, A2 => n3005, B1 => n3068, B2 => n3003
                           , ZN => n1508);
   U831 : OAI22_X1 port map( A1 => n4827, A2 => n3005, B1 => n3069, B2 => n3003
                           , ZN => n1507);
   U832 : OAI22_X1 port map( A1 => n4828, A2 => n3005, B1 => n3070, B2 => n3003
                           , ZN => n1506);
   U833 : OAI22_X1 port map( A1 => n5319, A2 => n3005, B1 => n3071, B2 => n3003
                           , ZN => n1505);
   U834 : OAI22_X1 port map( A1 => n5320, A2 => n3005, B1 => n3073, B2 => n3003
                           , ZN => n1504);
   U835 : OAI22_X1 port map( A1 => n5085, A2 => n3005, B1 => n3074, B2 => n3004
                           , ZN => n1503);
   U836 : OAI22_X1 port map( A1 => n5575, A2 => n3005, B1 => n3075, B2 => n3004
                           , ZN => n1502);
   U837 : OAI22_X1 port map( A1 => n4829, A2 => n3005, B1 => n3076, B2 => n3004
                           , ZN => n1501);
   U838 : OAI22_X1 port map( A1 => n5576, A2 => n3005, B1 => n3077, B2 => n3004
                           , ZN => n1500);
   U839 : OAI22_X1 port map( A1 => n4830, A2 => n3005, B1 => n3078, B2 => n3004
                           , ZN => n1499);
   U840 : OAI22_X1 port map( A1 => n5577, A2 => n3005, B1 => n3079, B2 => n3004
                           , ZN => n1498);
   U841 : OAI22_X1 port map( A1 => n4831, A2 => n3005, B1 => n3080, B2 => n3004
                           , ZN => n1497);
   U842 : OAI22_X1 port map( A1 => n4832, A2 => n3005, B1 => n3081, B2 => n3004
                           , ZN => n1496);
   U843 : OAI22_X1 port map( A1 => n5321, A2 => n3005, B1 => n3083, B2 => n3004
                           , ZN => n1495);
   U844 : NAND2_X1 port map( A1 => n3040, A2 => n3013, ZN => n3006);
   U845 : CLKBUF_X1 port map( A => n3006, Z => n3007);
   U846 : OAI22_X1 port map( A1 => n5165, A2 => n3008, B1 => n3014, B2 => n3007
                           , ZN => n1494);
   U847 : OAI22_X1 port map( A1 => n5322, A2 => n3008, B1 => n3051, B2 => n3006
                           , ZN => n1493);
   U848 : OAI22_X1 port map( A1 => n5323, A2 => n3008, B1 => n3052, B2 => n3007
                           , ZN => n1492);
   U849 : OAI22_X1 port map( A1 => n5324, A2 => n3008, B1 => n3053, B2 => n3006
                           , ZN => n1491);
   U850 : OAI22_X1 port map( A1 => n5578, A2 => n3008, B1 => n3054, B2 => n3007
                           , ZN => n1490);
   U851 : OAI22_X1 port map( A1 => n5325, A2 => n3008, B1 => n3055, B2 => n3006
                           , ZN => n1489);
   U852 : OAI22_X1 port map( A1 => n5579, A2 => n3008, B1 => n3056, B2 => n3007
                           , ZN => n1488);
   U853 : OAI22_X1 port map( A1 => n5580, A2 => n3008, B1 => n3057, B2 => n3006
                           , ZN => n1487);
   U854 : OAI22_X1 port map( A1 => n5581, A2 => n3008, B1 => n3058, B2 => n3007
                           , ZN => n1486);
   U855 : OAI22_X1 port map( A1 => n5086, A2 => n3008, B1 => n3059, B2 => n3006
                           , ZN => n1485);
   U856 : OAI22_X1 port map( A1 => n5582, A2 => n3008, B1 => n3060, B2 => n3006
                           , ZN => n1484);
   U857 : OAI22_X1 port map( A1 => n4833, A2 => n3008, B1 => n3061, B2 => n3007
                           , ZN => n1483);
   U858 : OAI22_X1 port map( A1 => n5583, A2 => n3008, B1 => n3062, B2 => n3006
                           , ZN => n1482);
   U859 : OAI22_X1 port map( A1 => n4834, A2 => n3008, B1 => n3063, B2 => n3007
                           , ZN => n1481);
   U860 : OAI22_X1 port map( A1 => n5584, A2 => n3008, B1 => n3064, B2 => n3006
                           , ZN => n1480);
   U861 : OAI22_X1 port map( A1 => n5326, A2 => n3008, B1 => n3065, B2 => n3007
                           , ZN => n1479);
   U862 : OAI22_X1 port map( A1 => n5087, A2 => n3008, B1 => n3066, B2 => n3006
                           , ZN => n1478);
   U863 : OAI22_X1 port map( A1 => n4835, A2 => n3008, B1 => n3067, B2 => n3006
                           , ZN => n1477);
   U864 : OAI22_X1 port map( A1 => n5585, A2 => n3008, B1 => n3068, B2 => n3006
                           , ZN => n1476);
   U865 : OAI22_X1 port map( A1 => n5088, A2 => n3008, B1 => n3069, B2 => n3006
                           , ZN => n1475);
   U866 : OAI22_X1 port map( A1 => n5586, A2 => n3008, B1 => n3070, B2 => n3006
                           , ZN => n1474);
   U867 : OAI22_X1 port map( A1 => n4836, A2 => n3008, B1 => n3071, B2 => n3006
                           , ZN => n1473);
   U868 : OAI22_X1 port map( A1 => n5587, A2 => n3008, B1 => n3073, B2 => n3006
                           , ZN => n1472);
   U869 : OAI22_X1 port map( A1 => n5588, A2 => n3008, B1 => n3074, B2 => n3007
                           , ZN => n1471);
   U870 : OAI22_X1 port map( A1 => n5089, A2 => n3008, B1 => n3075, B2 => n3007
                           , ZN => n1470);
   U871 : OAI22_X1 port map( A1 => n5327, A2 => n3008, B1 => n3076, B2 => n3007
                           , ZN => n1469);
   U872 : OAI22_X1 port map( A1 => n5589, A2 => n3008, B1 => n3077, B2 => n3007
                           , ZN => n1468);
   U873 : OAI22_X1 port map( A1 => n5590, A2 => n3008, B1 => n3078, B2 => n3007
                           , ZN => n1467);
   U874 : OAI22_X1 port map( A1 => n5328, A2 => n3008, B1 => n3079, B2 => n3007
                           , ZN => n1466);
   U875 : OAI22_X1 port map( A1 => n5090, A2 => n3008, B1 => n3080, B2 => n3007
                           , ZN => n1465);
   U876 : OAI22_X1 port map( A1 => n5591, A2 => n3008, B1 => n3081, B2 => n3007
                           , ZN => n1464);
   U877 : OAI22_X1 port map( A1 => n5329, A2 => n3008, B1 => n3083, B2 => n3007
                           , ZN => n1463);
   U878 : NAND2_X1 port map( A1 => n3044, A2 => n3013, ZN => n3009);
   U879 : CLKBUF_X1 port map( A => n3012, Z => n3010);
   U880 : CLKBUF_X1 port map( A => n3009, Z => n3011);
   U881 : OAI22_X1 port map( A1 => n5166, A2 => n3010, B1 => n3014, B2 => n3011
                           , ZN => n1462);
   U882 : OAI22_X1 port map( A1 => n5330, A2 => n3012, B1 => n3051, B2 => n3009
                           , ZN => n1461);
   U883 : OAI22_X1 port map( A1 => n5592, A2 => n3010, B1 => n3052, B2 => n3011
                           , ZN => n1460);
   U884 : OAI22_X1 port map( A1 => n5331, A2 => n3012, B1 => n3053, B2 => n3009
                           , ZN => n1459);
   U885 : OAI22_X1 port map( A1 => n5593, A2 => n3010, B1 => n3054, B2 => n3011
                           , ZN => n1458);
   U886 : OAI22_X1 port map( A1 => n5332, A2 => n3012, B1 => n3055, B2 => n3009
                           , ZN => n1457);
   U887 : OAI22_X1 port map( A1 => n5333, A2 => n3010, B1 => n3056, B2 => n3011
                           , ZN => n1456);
   U888 : OAI22_X1 port map( A1 => n5594, A2 => n3012, B1 => n3057, B2 => n3009
                           , ZN => n1455);
   U889 : OAI22_X1 port map( A1 => n5091, A2 => n3010, B1 => n3058, B2 => n3011
                           , ZN => n1454);
   U890 : OAI22_X1 port map( A1 => n5334, A2 => n3012, B1 => n3059, B2 => n3009
                           , ZN => n1453);
   U891 : OAI22_X1 port map( A1 => n5092, A2 => n3012, B1 => n3060, B2 => n3009
                           , ZN => n1452);
   U892 : OAI22_X1 port map( A1 => n5595, A2 => n3012, B1 => n3061, B2 => n3011
                           , ZN => n1451);
   U893 : OAI22_X1 port map( A1 => n5596, A2 => n3010, B1 => n3062, B2 => n3009
                           , ZN => n1450);
   U894 : OAI22_X1 port map( A1 => n4837, A2 => n3010, B1 => n3063, B2 => n3011
                           , ZN => n1449);
   U895 : OAI22_X1 port map( A1 => n5597, A2 => n3010, B1 => n3064, B2 => n3009
                           , ZN => n1448);
   U896 : OAI22_X1 port map( A1 => n5093, A2 => n3010, B1 => n3065, B2 => n3011
                           , ZN => n1447);
   U897 : OAI22_X1 port map( A1 => n5335, A2 => n3010, B1 => n3066, B2 => n3009
                           , ZN => n1446);
   U898 : OAI22_X1 port map( A1 => n5598, A2 => n3010, B1 => n3067, B2 => n3009
                           , ZN => n1445);
   U899 : OAI22_X1 port map( A1 => n5336, A2 => n3010, B1 => n3068, B2 => n3009
                           , ZN => n1444);
   U900 : OAI22_X1 port map( A1 => n5094, A2 => n3010, B1 => n3069, B2 => n3009
                           , ZN => n1443);
   U901 : OAI22_X1 port map( A1 => n5599, A2 => n3010, B1 => n3070, B2 => n3009
                           , ZN => n1442);
   U902 : OAI22_X1 port map( A1 => n5337, A2 => n3010, B1 => n3071, B2 => n3009
                           , ZN => n1441);
   U903 : OAI22_X1 port map( A1 => n5600, A2 => n3010, B1 => n3073, B2 => n3009
                           , ZN => n1440);
   U904 : OAI22_X1 port map( A1 => n5338, A2 => n3010, B1 => n3074, B2 => n3011
                           , ZN => n1439);
   U905 : OAI22_X1 port map( A1 => n5601, A2 => n3012, B1 => n3075, B2 => n3011
                           , ZN => n1438);
   U906 : OAI22_X1 port map( A1 => n5602, A2 => n3012, B1 => n3076, B2 => n3011
                           , ZN => n1437);
   U907 : OAI22_X1 port map( A1 => n4838, A2 => n3012, B1 => n3077, B2 => n3011
                           , ZN => n1436);
   U908 : OAI22_X1 port map( A1 => n5603, A2 => n3012, B1 => n3078, B2 => n3011
                           , ZN => n1435);
   U909 : OAI22_X1 port map( A1 => n5095, A2 => n3012, B1 => n3079, B2 => n3011
                           , ZN => n1434);
   U910 : OAI22_X1 port map( A1 => n5339, A2 => n3012, B1 => n3080, B2 => n3011
                           , ZN => n1433);
   U911 : OAI22_X1 port map( A1 => n5340, A2 => n3012, B1 => n3081, B2 => n3011
                           , ZN => n1432);
   U912 : OAI22_X1 port map( A1 => n5341, A2 => n3012, B1 => n3083, B2 => n3011
                           , ZN => n1431);
   U913 : NAND2_X1 port map( A1 => n3049, A2 => n3013, ZN => n3015);
   U914 : CLKBUF_X1 port map( A => n3015, Z => n3016);
   U915 : OAI22_X1 port map( A1 => n4648, A2 => n3017, B1 => n3014, B2 => n3016
                           , ZN => n1430);
   U916 : OAI22_X1 port map( A1 => n5096, A2 => n3017, B1 => n3051, B2 => n3015
                           , ZN => n1429);
   U917 : OAI22_X1 port map( A1 => n5097, A2 => n3017, B1 => n3052, B2 => n3016
                           , ZN => n1428);
   U918 : OAI22_X1 port map( A1 => n5098, A2 => n3017, B1 => n3053, B2 => n3015
                           , ZN => n1427);
   U919 : OAI22_X1 port map( A1 => n5099, A2 => n3017, B1 => n3054, B2 => n3016
                           , ZN => n1426);
   U920 : OAI22_X1 port map( A1 => n4839, A2 => n3017, B1 => n3055, B2 => n3015
                           , ZN => n1425);
   U921 : OAI22_X1 port map( A1 => n4840, A2 => n3017, B1 => n3056, B2 => n3016
                           , ZN => n1424);
   U922 : OAI22_X1 port map( A1 => n4841, A2 => n3017, B1 => n3057, B2 => n3015
                           , ZN => n1423);
   U923 : OAI22_X1 port map( A1 => n4842, A2 => n3017, B1 => n3058, B2 => n3016
                           , ZN => n1422);
   U924 : OAI22_X1 port map( A1 => n4843, A2 => n3017, B1 => n3059, B2 => n3015
                           , ZN => n1421);
   U925 : OAI22_X1 port map( A1 => n5100, A2 => n3017, B1 => n3060, B2 => n3015
                           , ZN => n1420);
   U926 : OAI22_X1 port map( A1 => n4844, A2 => n3017, B1 => n3061, B2 => n3016
                           , ZN => n1419);
   U927 : OAI22_X1 port map( A1 => n5101, A2 => n3017, B1 => n3062, B2 => n3015
                           , ZN => n1418);
   U928 : OAI22_X1 port map( A1 => n5102, A2 => n3017, B1 => n3063, B2 => n3016
                           , ZN => n1417);
   U929 : OAI22_X1 port map( A1 => n5103, A2 => n3017, B1 => n3064, B2 => n3015
                           , ZN => n1416);
   U930 : OAI22_X1 port map( A1 => n4845, A2 => n3017, B1 => n3065, B2 => n3016
                           , ZN => n1415);
   U931 : OAI22_X1 port map( A1 => n4846, A2 => n3017, B1 => n3066, B2 => n3015
                           , ZN => n1414);
   U932 : OAI22_X1 port map( A1 => n4847, A2 => n3017, B1 => n3067, B2 => n3015
                           , ZN => n1413);
   U933 : OAI22_X1 port map( A1 => n5604, A2 => n3017, B1 => n3068, B2 => n3015
                           , ZN => n1412);
   U934 : OAI22_X1 port map( A1 => n4848, A2 => n3017, B1 => n3069, B2 => n3015
                           , ZN => n1411);
   U935 : OAI22_X1 port map( A1 => n4849, A2 => n3017, B1 => n3070, B2 => n3015
                           , ZN => n1410);
   U936 : OAI22_X1 port map( A1 => n4850, A2 => n3017, B1 => n3071, B2 => n3015
                           , ZN => n1409);
   U937 : OAI22_X1 port map( A1 => n5104, A2 => n3017, B1 => n3073, B2 => n3015
                           , ZN => n1408);
   U938 : OAI22_X1 port map( A1 => n5105, A2 => n3017, B1 => n3074, B2 => n3016
                           , ZN => n1407);
   U939 : OAI22_X1 port map( A1 => n5106, A2 => n3017, B1 => n3075, B2 => n3016
                           , ZN => n1406);
   U940 : OAI22_X1 port map( A1 => n5342, A2 => n3017, B1 => n3076, B2 => n3016
                           , ZN => n1405);
   U941 : OAI22_X1 port map( A1 => n5107, A2 => n3017, B1 => n3077, B2 => n3016
                           , ZN => n1404);
   U942 : OAI22_X1 port map( A1 => n4851, A2 => n3017, B1 => n3078, B2 => n3016
                           , ZN => n1403);
   U943 : OAI22_X1 port map( A1 => n5108, A2 => n3017, B1 => n3079, B2 => n3016
                           , ZN => n1402);
   U944 : OAI22_X1 port map( A1 => n5605, A2 => n3017, B1 => n3080, B2 => n3016
                           , ZN => n1401);
   U945 : OAI22_X1 port map( A1 => n4852, A2 => n3017, B1 => n3081, B2 => n3016
                           , ZN => n1400);
   U946 : OAI22_X1 port map( A1 => n4853, A2 => n3017, B1 => n3083, B2 => n3016
                           , ZN => n1399);
   U947 : NOR2_X1 port map( A1 => n3019, A2 => n3018, ZN => n3048);
   U948 : NAND2_X1 port map( A1 => n3020, A2 => n3048, ZN => n3021);
   U949 : CLKBUF_X1 port map( A => n3021, Z => n3022);
   U950 : OAI22_X1 port map( A1 => n5167, A2 => n3023, B1 => n3050, B2 => n3022
                           , ZN => n1398);
   U951 : OAI22_X1 port map( A1 => n5606, A2 => n3023, B1 => n3051, B2 => n3021
                           , ZN => n1397);
   U952 : OAI22_X1 port map( A1 => n5343, A2 => n3023, B1 => n3052, B2 => n3022
                           , ZN => n1396);
   U953 : OAI22_X1 port map( A1 => n5607, A2 => n3023, B1 => n3053, B2 => n3021
                           , ZN => n1395);
   U954 : OAI22_X1 port map( A1 => n5608, A2 => n3023, B1 => n3054, B2 => n3022
                           , ZN => n1394);
   U955 : OAI22_X1 port map( A1 => n5609, A2 => n3023, B1 => n3055, B2 => n3021
                           , ZN => n1393);
   U956 : OAI22_X1 port map( A1 => n5344, A2 => n3023, B1 => n3056, B2 => n3022
                           , ZN => n1392);
   U957 : OAI22_X1 port map( A1 => n5345, A2 => n3023, B1 => n3057, B2 => n3021
                           , ZN => n1391);
   U958 : OAI22_X1 port map( A1 => n5346, A2 => n3023, B1 => n3058, B2 => n3022
                           , ZN => n1390);
   U959 : OAI22_X1 port map( A1 => n5610, A2 => n3023, B1 => n3059, B2 => n3021
                           , ZN => n1389);
   U960 : OAI22_X1 port map( A1 => n5611, A2 => n3023, B1 => n3060, B2 => n3021
                           , ZN => n1388);
   U961 : OAI22_X1 port map( A1 => n5347, A2 => n3023, B1 => n3061, B2 => n3022
                           , ZN => n1387);
   U962 : OAI22_X1 port map( A1 => n5348, A2 => n3023, B1 => n3062, B2 => n3021
                           , ZN => n1386);
   U963 : OAI22_X1 port map( A1 => n5349, A2 => n3023, B1 => n3063, B2 => n3022
                           , ZN => n1385);
   U964 : OAI22_X1 port map( A1 => n5350, A2 => n3023, B1 => n3064, B2 => n3021
                           , ZN => n1384);
   U965 : OAI22_X1 port map( A1 => n5351, A2 => n3023, B1 => n3065, B2 => n3022
                           , ZN => n1383);
   U966 : OAI22_X1 port map( A1 => n5352, A2 => n3023, B1 => n3066, B2 => n3021
                           , ZN => n1382);
   U967 : OAI22_X1 port map( A1 => n5353, A2 => n3023, B1 => n3067, B2 => n3021
                           , ZN => n1381);
   U968 : OAI22_X1 port map( A1 => n5612, A2 => n3023, B1 => n3068, B2 => n3021
                           , ZN => n1380);
   U969 : OAI22_X1 port map( A1 => n5613, A2 => n3023, B1 => n3069, B2 => n3021
                           , ZN => n1379);
   U970 : OAI22_X1 port map( A1 => n5354, A2 => n3023, B1 => n3070, B2 => n3021
                           , ZN => n1378);
   U971 : OAI22_X1 port map( A1 => n5614, A2 => n3023, B1 => n3071, B2 => n3021
                           , ZN => n1377);
   U972 : OAI22_X1 port map( A1 => n5355, A2 => n3023, B1 => n3073, B2 => n3021
                           , ZN => n1376);
   U973 : OAI22_X1 port map( A1 => n5615, A2 => n3023, B1 => n3074, B2 => n3022
                           , ZN => n1375);
   U974 : OAI22_X1 port map( A1 => n5356, A2 => n3023, B1 => n3075, B2 => n3022
                           , ZN => n1374);
   U975 : OAI22_X1 port map( A1 => n5616, A2 => n3023, B1 => n3076, B2 => n3022
                           , ZN => n1373);
   U976 : OAI22_X1 port map( A1 => n5357, A2 => n3023, B1 => n3077, B2 => n3022
                           , ZN => n1372);
   U977 : OAI22_X1 port map( A1 => n5358, A2 => n3023, B1 => n3078, B2 => n3022
                           , ZN => n1371);
   U978 : OAI22_X1 port map( A1 => n5617, A2 => n3023, B1 => n3079, B2 => n3022
                           , ZN => n1370);
   U979 : OAI22_X1 port map( A1 => n5359, A2 => n3023, B1 => n3080, B2 => n3022
                           , ZN => n1369);
   U980 : OAI22_X1 port map( A1 => n5360, A2 => n3023, B1 => n3081, B2 => n3022
                           , ZN => n1368);
   U981 : OAI22_X1 port map( A1 => n5361, A2 => n3023, B1 => n3083, B2 => n3022
                           , ZN => n1367);
   U982 : NAND2_X1 port map( A1 => n3024, A2 => n3048, ZN => n3025);
   U983 : CLKBUF_X1 port map( A => n3025, Z => n3026);
   U984 : OAI22_X1 port map( A1 => n4920, A2 => n3027, B1 => n3050, B2 => n3026
                           , ZN => n1366);
   U985 : OAI22_X1 port map( A1 => n5109, A2 => n3027, B1 => n3051, B2 => n3025
                           , ZN => n1365);
   U986 : OAI22_X1 port map( A1 => n4854, A2 => n3027, B1 => n3052, B2 => n3026
                           , ZN => n1364);
   U987 : OAI22_X1 port map( A1 => n4855, A2 => n3027, B1 => n3053, B2 => n3025
                           , ZN => n1363);
   U988 : OAI22_X1 port map( A1 => n5110, A2 => n3027, B1 => n3054, B2 => n3026
                           , ZN => n1362);
   U989 : OAI22_X1 port map( A1 => n4856, A2 => n3027, B1 => n3055, B2 => n3025
                           , ZN => n1361);
   U990 : OAI22_X1 port map( A1 => n4857, A2 => n3027, B1 => n3056, B2 => n3026
                           , ZN => n1360);
   U991 : OAI22_X1 port map( A1 => n4858, A2 => n3027, B1 => n3057, B2 => n3025
                           , ZN => n1359);
   U992 : OAI22_X1 port map( A1 => n4859, A2 => n3027, B1 => n3058, B2 => n3026
                           , ZN => n1358);
   U993 : OAI22_X1 port map( A1 => n5111, A2 => n3027, B1 => n3059, B2 => n3025
                           , ZN => n1357);
   U994 : OAI22_X1 port map( A1 => n5362, A2 => n3027, B1 => n3060, B2 => n3025
                           , ZN => n1356);
   U995 : OAI22_X1 port map( A1 => n4860, A2 => n3027, B1 => n3061, B2 => n3026
                           , ZN => n1355);
   U996 : OAI22_X1 port map( A1 => n5363, A2 => n3027, B1 => n3062, B2 => n3025
                           , ZN => n1354);
   U997 : OAI22_X1 port map( A1 => n5364, A2 => n3027, B1 => n3063, B2 => n3026
                           , ZN => n1353);
   U998 : OAI22_X1 port map( A1 => n4861, A2 => n3027, B1 => n3064, B2 => n3025
                           , ZN => n1352);
   U999 : OAI22_X1 port map( A1 => n4862, A2 => n3027, B1 => n3065, B2 => n3026
                           , ZN => n1351);
   U1000 : OAI22_X1 port map( A1 => n4863, A2 => n3027, B1 => n3066, B2 => 
                           n3025, ZN => n1350);
   U1001 : OAI22_X1 port map( A1 => n4864, A2 => n3027, B1 => n3067, B2 => 
                           n3025, ZN => n1349);
   U1002 : OAI22_X1 port map( A1 => n5112, A2 => n3027, B1 => n3068, B2 => 
                           n3025, ZN => n1348);
   U1003 : OAI22_X1 port map( A1 => n5113, A2 => n3027, B1 => n3069, B2 => 
                           n3025, ZN => n1347);
   U1004 : OAI22_X1 port map( A1 => n5114, A2 => n3027, B1 => n3070, B2 => 
                           n3025, ZN => n1346);
   U1005 : OAI22_X1 port map( A1 => n4865, A2 => n3027, B1 => n3071, B2 => 
                           n3025, ZN => n1345);
   U1006 : OAI22_X1 port map( A1 => n4866, A2 => n3027, B1 => n3073, B2 => 
                           n3025, ZN => n1344);
   U1007 : OAI22_X1 port map( A1 => n5365, A2 => n3027, B1 => n3074, B2 => 
                           n3026, ZN => n1343);
   U1008 : OAI22_X1 port map( A1 => n4867, A2 => n3027, B1 => n3075, B2 => 
                           n3026, ZN => n1342);
   U1009 : OAI22_X1 port map( A1 => n5115, A2 => n3027, B1 => n3076, B2 => 
                           n3026, ZN => n1341);
   U1010 : OAI22_X1 port map( A1 => n5116, A2 => n3027, B1 => n3077, B2 => 
                           n3026, ZN => n1340);
   U1011 : OAI22_X1 port map( A1 => n4868, A2 => n3027, B1 => n3078, B2 => 
                           n3026, ZN => n1339);
   U1012 : OAI22_X1 port map( A1 => n4869, A2 => n3027, B1 => n3079, B2 => 
                           n3026, ZN => n1338);
   U1013 : OAI22_X1 port map( A1 => n5117, A2 => n3027, B1 => n3080, B2 => 
                           n3026, ZN => n1337);
   U1014 : OAI22_X1 port map( A1 => n5618, A2 => n3027, B1 => n3081, B2 => 
                           n3026, ZN => n1336);
   U1015 : OAI22_X1 port map( A1 => n4870, A2 => n3027, B1 => n3083, B2 => 
                           n3026, ZN => n1335);
   U1016 : NAND2_X1 port map( A1 => n3028, A2 => n3048, ZN => n3029);
   U1017 : OAI22_X1 port map( A1 => n4921, A2 => n3031, B1 => n3050, B2 => 
                           n3030, ZN => n1334);
   U1018 : OAI22_X1 port map( A1 => n5619, A2 => n3031, B1 => n3051, B2 => 
                           n3029, ZN => n1333);
   U1019 : OAI22_X1 port map( A1 => n4871, A2 => n3031, B1 => n3052, B2 => 
                           n3030, ZN => n1332);
   U1020 : OAI22_X1 port map( A1 => n4872, A2 => n3031, B1 => n3053, B2 => 
                           n3029, ZN => n1331);
   U1021 : OAI22_X1 port map( A1 => n4873, A2 => n3031, B1 => n3054, B2 => 
                           n3030, ZN => n1330);
   U1022 : OAI22_X1 port map( A1 => n5366, A2 => n3031, B1 => n3055, B2 => 
                           n3029, ZN => n1329);
   U1023 : OAI22_X1 port map( A1 => n5118, A2 => n3031, B1 => n3056, B2 => 
                           n3030, ZN => n1328);
   U1024 : OAI22_X1 port map( A1 => n4874, A2 => n3031, B1 => n3057, B2 => 
                           n3029, ZN => n1327);
   U1025 : OAI22_X1 port map( A1 => n5367, A2 => n3031, B1 => n3058, B2 => 
                           n3030, ZN => n1326);
   U1026 : OAI22_X1 port map( A1 => n5368, A2 => n3031, B1 => n3059, B2 => 
                           n3029, ZN => n1325);
   U1027 : OAI22_X1 port map( A1 => n5369, A2 => n3031, B1 => n3060, B2 => 
                           n3029, ZN => n1324);
   U1028 : OAI22_X1 port map( A1 => n4875, A2 => n3031, B1 => n3061, B2 => 
                           n3030, ZN => n1323);
   U1029 : OAI22_X1 port map( A1 => n5119, A2 => n3031, B1 => n3062, B2 => 
                           n3029, ZN => n1322);
   U1030 : OAI22_X1 port map( A1 => n5620, A2 => n3031, B1 => n3063, B2 => 
                           n3030, ZN => n1321);
   U1031 : OAI22_X1 port map( A1 => n5120, A2 => n3031, B1 => n3064, B2 => 
                           n3029, ZN => n1320);
   U1032 : OAI22_X1 port map( A1 => n5121, A2 => n3031, B1 => n3065, B2 => 
                           n3030, ZN => n1319);
   U1033 : OAI22_X1 port map( A1 => n5122, A2 => n3031, B1 => n3066, B2 => 
                           n3029, ZN => n1318);
   U1034 : OAI22_X1 port map( A1 => n4876, A2 => n3031, B1 => n3067, B2 => 
                           n3029, ZN => n1317);
   U1035 : OAI22_X1 port map( A1 => n4877, A2 => n3031, B1 => n3068, B2 => 
                           n3029, ZN => n1316);
   U1036 : OAI22_X1 port map( A1 => n5370, A2 => n3031, B1 => n3069, B2 => 
                           n3029, ZN => n1315);
   U1037 : OAI22_X1 port map( A1 => n5621, A2 => n3031, B1 => n3070, B2 => 
                           n3029, ZN => n1314);
   U1038 : OAI22_X1 port map( A1 => n5123, A2 => n3031, B1 => n3071, B2 => 
                           n3029, ZN => n1313);
   U1039 : OAI22_X1 port map( A1 => n5622, A2 => n3031, B1 => n3073, B2 => 
                           n3029, ZN => n1312);
   U1040 : OAI22_X1 port map( A1 => n5124, A2 => n3031, B1 => n3074, B2 => 
                           n3030, ZN => n1311);
   U1041 : OAI22_X1 port map( A1 => n5623, A2 => n3031, B1 => n3075, B2 => 
                           n3030, ZN => n1310);
   U1042 : OAI22_X1 port map( A1 => n5624, A2 => n3031, B1 => n3076, B2 => 
                           n3030, ZN => n1309);
   U1043 : OAI22_X1 port map( A1 => n4878, A2 => n3031, B1 => n3077, B2 => 
                           n3030, ZN => n1308);
   U1044 : OAI22_X1 port map( A1 => n5625, A2 => n3031, B1 => n3078, B2 => 
                           n3030, ZN => n1307);
   U1045 : OAI22_X1 port map( A1 => n5125, A2 => n3031, B1 => n3079, B2 => 
                           n3030, ZN => n1306);
   U1046 : OAI22_X1 port map( A1 => n5626, A2 => n3031, B1 => n3080, B2 => 
                           n3030, ZN => n1305);
   U1047 : OAI22_X1 port map( A1 => n5126, A2 => n3031, B1 => n3081, B2 => 
                           n3030, ZN => n1304);
   U1048 : OAI22_X1 port map( A1 => n5627, A2 => n3031, B1 => n3083, B2 => 
                           n3030, ZN => n1303);
   U1049 : NAND2_X1 port map( A1 => n3032, A2 => n3048, ZN => n3033);
   U1050 : CLKBUF_X1 port map( A => n3033, Z => n3034);
   U1051 : OAI22_X1 port map( A1 => n4649, A2 => n3035, B1 => n3050, B2 => 
                           n3034, ZN => n1302);
   U1052 : OAI22_X1 port map( A1 => n5127, A2 => n3035, B1 => n3051, B2 => 
                           n3033, ZN => n1301);
   U1053 : OAI22_X1 port map( A1 => n5128, A2 => n3035, B1 => n3052, B2 => 
                           n3034, ZN => n1300);
   U1054 : OAI22_X1 port map( A1 => n5129, A2 => n3035, B1 => n3053, B2 => 
                           n3033, ZN => n1299);
   U1055 : OAI22_X1 port map( A1 => n5130, A2 => n3035, B1 => n3054, B2 => 
                           n3034, ZN => n1298);
   U1056 : OAI22_X1 port map( A1 => n5131, A2 => n3035, B1 => n3055, B2 => 
                           n3033, ZN => n1297);
   U1057 : OAI22_X1 port map( A1 => n4879, A2 => n3035, B1 => n3056, B2 => 
                           n3034, ZN => n1296);
   U1058 : OAI22_X1 port map( A1 => n5132, A2 => n3035, B1 => n3057, B2 => 
                           n3033, ZN => n1295);
   U1059 : OAI22_X1 port map( A1 => n4880, A2 => n3035, B1 => n3058, B2 => 
                           n3034, ZN => n1294);
   U1060 : OAI22_X1 port map( A1 => n4881, A2 => n3035, B1 => n3059, B2 => 
                           n3033, ZN => n1293);
   U1061 : OAI22_X1 port map( A1 => n5133, A2 => n3035, B1 => n3060, B2 => 
                           n3033, ZN => n1292);
   U1062 : OAI22_X1 port map( A1 => n5134, A2 => n3035, B1 => n3061, B2 => 
                           n3034, ZN => n1291);
   U1063 : OAI22_X1 port map( A1 => n4882, A2 => n3035, B1 => n3062, B2 => 
                           n3033, ZN => n1290);
   U1064 : OAI22_X1 port map( A1 => n5135, A2 => n3035, B1 => n3063, B2 => 
                           n3034, ZN => n1289);
   U1065 : OAI22_X1 port map( A1 => n4883, A2 => n3035, B1 => n3064, B2 => 
                           n3033, ZN => n1288);
   U1066 : OAI22_X1 port map( A1 => n4884, A2 => n3035, B1 => n3065, B2 => 
                           n3034, ZN => n1287);
   U1067 : OAI22_X1 port map( A1 => n5136, A2 => n3035, B1 => n3066, B2 => 
                           n3033, ZN => n1286);
   U1068 : OAI22_X1 port map( A1 => n4885, A2 => n3035, B1 => n3067, B2 => 
                           n3033, ZN => n1285);
   U1069 : OAI22_X1 port map( A1 => n4886, A2 => n3035, B1 => n3068, B2 => 
                           n3033, ZN => n1284);
   U1070 : OAI22_X1 port map( A1 => n4887, A2 => n3035, B1 => n3069, B2 => 
                           n3033, ZN => n1283);
   U1071 : OAI22_X1 port map( A1 => n4888, A2 => n3035, B1 => n3070, B2 => 
                           n3033, ZN => n1282);
   U1072 : OAI22_X1 port map( A1 => n5137, A2 => n3035, B1 => n3071, B2 => 
                           n3033, ZN => n1281);
   U1073 : OAI22_X1 port map( A1 => n4889, A2 => n3035, B1 => n3073, B2 => 
                           n3033, ZN => n1280);
   U1074 : OAI22_X1 port map( A1 => n5138, A2 => n3035, B1 => n3074, B2 => 
                           n3034, ZN => n1279);
   U1075 : OAI22_X1 port map( A1 => n4890, A2 => n3035, B1 => n3075, B2 => 
                           n3034, ZN => n1278);
   U1076 : OAI22_X1 port map( A1 => n4891, A2 => n3035, B1 => n3076, B2 => 
                           n3034, ZN => n1277);
   U1077 : OAI22_X1 port map( A1 => n5139, A2 => n3035, B1 => n3077, B2 => 
                           n3034, ZN => n1276);
   U1078 : OAI22_X1 port map( A1 => n4892, A2 => n3035, B1 => n3078, B2 => 
                           n3034, ZN => n1275);
   U1079 : OAI22_X1 port map( A1 => n4893, A2 => n3035, B1 => n3079, B2 => 
                           n3034, ZN => n1274);
   U1080 : OAI22_X1 port map( A1 => n5140, A2 => n3035, B1 => n3080, B2 => 
                           n3034, ZN => n1273);
   U1081 : OAI22_X1 port map( A1 => n4894, A2 => n3035, B1 => n3081, B2 => 
                           n3034, ZN => n1272);
   U1082 : OAI22_X1 port map( A1 => n5141, A2 => n3035, B1 => n3083, B2 => 
                           n3034, ZN => n1271);
   U1083 : NAND2_X1 port map( A1 => n3036, A2 => n3048, ZN => n3037);
   U1084 : CLKBUF_X1 port map( A => n3037, Z => n3038);
   U1085 : OAI22_X1 port map( A1 => n4922, A2 => n3039, B1 => n3050, B2 => 
                           n3038, ZN => n1270);
   U1086 : OAI22_X1 port map( A1 => n5371, A2 => n3039, B1 => n3051, B2 => 
                           n3037, ZN => n1269);
   U1087 : OAI22_X1 port map( A1 => n5628, A2 => n3039, B1 => n3052, B2 => 
                           n3038, ZN => n1268);
   U1088 : OAI22_X1 port map( A1 => n5372, A2 => n3039, B1 => n3053, B2 => 
                           n3037, ZN => n1267);
   U1089 : OAI22_X1 port map( A1 => n5373, A2 => n3039, B1 => n3054, B2 => 
                           n3038, ZN => n1266);
   U1090 : OAI22_X1 port map( A1 => n5629, A2 => n3039, B1 => n3055, B2 => 
                           n3037, ZN => n1265);
   U1091 : OAI22_X1 port map( A1 => n5630, A2 => n3039, B1 => n3056, B2 => 
                           n3038, ZN => n1264);
   U1092 : OAI22_X1 port map( A1 => n5374, A2 => n3039, B1 => n3057, B2 => 
                           n3037, ZN => n1263);
   U1093 : OAI22_X1 port map( A1 => n5631, A2 => n3039, B1 => n3058, B2 => 
                           n3038, ZN => n1262);
   U1094 : OAI22_X1 port map( A1 => n5375, A2 => n3039, B1 => n3059, B2 => 
                           n3037, ZN => n1261);
   U1095 : OAI22_X1 port map( A1 => n5632, A2 => n3039, B1 => n3060, B2 => 
                           n3037, ZN => n1260);
   U1096 : OAI22_X1 port map( A1 => n5633, A2 => n3039, B1 => n3061, B2 => 
                           n3038, ZN => n1259);
   U1097 : OAI22_X1 port map( A1 => n5634, A2 => n3039, B1 => n3062, B2 => 
                           n3037, ZN => n1258);
   U1098 : OAI22_X1 port map( A1 => n5635, A2 => n3039, B1 => n3063, B2 => 
                           n3038, ZN => n1257);
   U1099 : OAI22_X1 port map( A1 => n4895, A2 => n3039, B1 => n3064, B2 => 
                           n3037, ZN => n1256);
   U1100 : OAI22_X1 port map( A1 => n5636, A2 => n3039, B1 => n3065, B2 => 
                           n3038, ZN => n1255);
   U1101 : OAI22_X1 port map( A1 => n5376, A2 => n3039, B1 => n3066, B2 => 
                           n3037, ZN => n1254);
   U1102 : OAI22_X1 port map( A1 => n5637, A2 => n3039, B1 => n3067, B2 => 
                           n3037, ZN => n1253);
   U1103 : OAI22_X1 port map( A1 => n5377, A2 => n3039, B1 => n3068, B2 => 
                           n3037, ZN => n1252);
   U1104 : OAI22_X1 port map( A1 => n5638, A2 => n3039, B1 => n3069, B2 => 
                           n3037, ZN => n1251);
   U1105 : OAI22_X1 port map( A1 => n5378, A2 => n3039, B1 => n3070, B2 => 
                           n3037, ZN => n1250);
   U1106 : OAI22_X1 port map( A1 => n5639, A2 => n3039, B1 => n3071, B2 => 
                           n3037, ZN => n1249);
   U1107 : OAI22_X1 port map( A1 => n5142, A2 => n3039, B1 => n3073, B2 => 
                           n3037, ZN => n1248);
   U1108 : OAI22_X1 port map( A1 => n5640, A2 => n3039, B1 => n3074, B2 => 
                           n3038, ZN => n1247);
   U1109 : OAI22_X1 port map( A1 => n5641, A2 => n3039, B1 => n3075, B2 => 
                           n3038, ZN => n1246);
   U1110 : OAI22_X1 port map( A1 => n4896, A2 => n3039, B1 => n3076, B2 => 
                           n3038, ZN => n1245);
   U1111 : OAI22_X1 port map( A1 => n5379, A2 => n3039, B1 => n3077, B2 => 
                           n3038, ZN => n1244);
   U1112 : OAI22_X1 port map( A1 => n5642, A2 => n3039, B1 => n3078, B2 => 
                           n3038, ZN => n1243);
   U1113 : OAI22_X1 port map( A1 => n5643, A2 => n3039, B1 => n3079, B2 => 
                           n3038, ZN => n1242);
   U1114 : OAI22_X1 port map( A1 => n5380, A2 => n3039, B1 => n3080, B2 => 
                           n3038, ZN => n1241);
   U1115 : OAI22_X1 port map( A1 => n5644, A2 => n3039, B1 => n3081, B2 => 
                           n3038, ZN => n1240);
   U1116 : OAI22_X1 port map( A1 => n5645, A2 => n3039, B1 => n3083, B2 => 
                           n3038, ZN => n1239);
   U1117 : NAND2_X1 port map( A1 => n3040, A2 => n3048, ZN => n3041);
   U1118 : CLKBUF_X1 port map( A => n3041, Z => n3042);
   U1119 : OAI22_X1 port map( A1 => n4923, A2 => n3043, B1 => n3050, B2 => 
                           n3042, ZN => n1238);
   U1120 : OAI22_X1 port map( A1 => n5646, A2 => n3043, B1 => n3051, B2 => 
                           n3041, ZN => n1237);
   U1121 : OAI22_X1 port map( A1 => n5143, A2 => n3043, B1 => n3052, B2 => 
                           n3042, ZN => n1236);
   U1122 : OAI22_X1 port map( A1 => n5381, A2 => n3043, B1 => n3053, B2 => 
                           n3041, ZN => n1235);
   U1123 : OAI22_X1 port map( A1 => n5382, A2 => n3043, B1 => n3054, B2 => 
                           n3042, ZN => n1234);
   U1124 : OAI22_X1 port map( A1 => n5144, A2 => n3043, B1 => n3055, B2 => 
                           n3041, ZN => n1233);
   U1125 : OAI22_X1 port map( A1 => n5383, A2 => n3043, B1 => n3056, B2 => 
                           n3042, ZN => n1232);
   U1126 : OAI22_X1 port map( A1 => n5647, A2 => n3043, B1 => n3057, B2 => 
                           n3041, ZN => n1231);
   U1127 : OAI22_X1 port map( A1 => n5648, A2 => n3043, B1 => n3058, B2 => 
                           n3042, ZN => n1230);
   U1128 : OAI22_X1 port map( A1 => n5649, A2 => n3043, B1 => n3059, B2 => 
                           n3041, ZN => n1229);
   U1129 : OAI22_X1 port map( A1 => n5650, A2 => n3043, B1 => n3060, B2 => 
                           n3041, ZN => n1228);
   U1130 : OAI22_X1 port map( A1 => n5651, A2 => n3043, B1 => n3061, B2 => 
                           n3042, ZN => n1227);
   U1131 : OAI22_X1 port map( A1 => n5384, A2 => n3043, B1 => n3062, B2 => 
                           n3041, ZN => n1226);
   U1132 : OAI22_X1 port map( A1 => n5385, A2 => n3043, B1 => n3063, B2 => 
                           n3042, ZN => n1225);
   U1133 : OAI22_X1 port map( A1 => n5652, A2 => n3043, B1 => n3064, B2 => 
                           n3041, ZN => n1224);
   U1134 : OAI22_X1 port map( A1 => n5653, A2 => n3043, B1 => n3065, B2 => 
                           n3042, ZN => n1223);
   U1135 : OAI22_X1 port map( A1 => n5386, A2 => n3043, B1 => n3066, B2 => 
                           n3041, ZN => n1222);
   U1136 : OAI22_X1 port map( A1 => n5654, A2 => n3043, B1 => n3067, B2 => 
                           n3041, ZN => n1221);
   U1137 : OAI22_X1 port map( A1 => n5387, A2 => n3043, B1 => n3068, B2 => 
                           n3041, ZN => n1220);
   U1138 : OAI22_X1 port map( A1 => n5655, A2 => n3043, B1 => n3069, B2 => 
                           n3041, ZN => n1219);
   U1139 : OAI22_X1 port map( A1 => n5388, A2 => n3043, B1 => n3070, B2 => 
                           n3041, ZN => n1218);
   U1140 : OAI22_X1 port map( A1 => n5656, A2 => n3043, B1 => n3071, B2 => 
                           n3041, ZN => n1217);
   U1141 : OAI22_X1 port map( A1 => n5389, A2 => n3043, B1 => n3073, B2 => 
                           n3041, ZN => n1216);
   U1142 : OAI22_X1 port map( A1 => n5390, A2 => n3043, B1 => n3074, B2 => 
                           n3042, ZN => n1215);
   U1143 : OAI22_X1 port map( A1 => n5391, A2 => n3043, B1 => n3075, B2 => 
                           n3042, ZN => n1214);
   U1144 : OAI22_X1 port map( A1 => n5145, A2 => n3043, B1 => n3076, B2 => 
                           n3042, ZN => n1213);
   U1145 : OAI22_X1 port map( A1 => n5392, A2 => n3043, B1 => n3077, B2 => 
                           n3042, ZN => n1212);
   U1146 : OAI22_X1 port map( A1 => n5393, A2 => n3043, B1 => n3078, B2 => 
                           n3042, ZN => n1211);
   U1147 : OAI22_X1 port map( A1 => n5657, A2 => n3043, B1 => n3079, B2 => 
                           n3042, ZN => n1210);
   U1148 : OAI22_X1 port map( A1 => n5394, A2 => n3043, B1 => n3080, B2 => 
                           n3042, ZN => n1209);
   U1149 : OAI22_X1 port map( A1 => n5658, A2 => n3043, B1 => n3081, B2 => 
                           n3042, ZN => n1208);
   U1150 : OAI22_X1 port map( A1 => n5395, A2 => n3043, B1 => n3083, B2 => 
                           n3042, ZN => n1207);
   U1151 : NAND2_X1 port map( A1 => n3044, A2 => n3048, ZN => n3045);
   U1152 : CLKBUF_X1 port map( A => n3045, Z => n3046);
   U1153 : OAI22_X1 port map( A1 => n4650, A2 => n3047, B1 => n3050, B2 => 
                           n3046, ZN => n1206);
   U1154 : OAI22_X1 port map( A1 => n4897, A2 => n3047, B1 => n3051, B2 => 
                           n3045, ZN => n1205);
   U1155 : OAI22_X1 port map( A1 => n4898, A2 => n3047, B1 => n3052, B2 => 
                           n3046, ZN => n1204);
   U1156 : OAI22_X1 port map( A1 => n5659, A2 => n3047, B1 => n3053, B2 => 
                           n3045, ZN => n1203);
   U1157 : OAI22_X1 port map( A1 => n4899, A2 => n3047, B1 => n3054, B2 => 
                           n3046, ZN => n1202);
   U1158 : OAI22_X1 port map( A1 => n5146, A2 => n3047, B1 => n3055, B2 => 
                           n3045, ZN => n1201);
   U1159 : OAI22_X1 port map( A1 => n5660, A2 => n3047, B1 => n3056, B2 => 
                           n3046, ZN => n1200);
   U1160 : OAI22_X1 port map( A1 => n5147, A2 => n3047, B1 => n3057, B2 => 
                           n3045, ZN => n1199);
   U1161 : OAI22_X1 port map( A1 => n5396, A2 => n3047, B1 => n3058, B2 => 
                           n3046, ZN => n1198);
   U1162 : OAI22_X1 port map( A1 => n4900, A2 => n3047, B1 => n3059, B2 => 
                           n3045, ZN => n1197);
   U1163 : OAI22_X1 port map( A1 => n4901, A2 => n3047, B1 => n3060, B2 => 
                           n3045, ZN => n1196);
   U1164 : OAI22_X1 port map( A1 => n5397, A2 => n3047, B1 => n3061, B2 => 
                           n3046, ZN => n1195);
   U1165 : OAI22_X1 port map( A1 => n5661, A2 => n3047, B1 => n3062, B2 => 
                           n3045, ZN => n1194);
   U1166 : OAI22_X1 port map( A1 => n5148, A2 => n3047, B1 => n3063, B2 => 
                           n3046, ZN => n1193);
   U1167 : OAI22_X1 port map( A1 => n4902, A2 => n3047, B1 => n3064, B2 => 
                           n3045, ZN => n1192);
   U1168 : OAI22_X1 port map( A1 => n5398, A2 => n3047, B1 => n3065, B2 => 
                           n3046, ZN => n1191);
   U1169 : OAI22_X1 port map( A1 => n4903, A2 => n3047, B1 => n3066, B2 => 
                           n3045, ZN => n1190);
   U1170 : OAI22_X1 port map( A1 => n5662, A2 => n3047, B1 => n3067, B2 => 
                           n3045, ZN => n1189);
   U1171 : OAI22_X1 port map( A1 => n5663, A2 => n3047, B1 => n3068, B2 => 
                           n3045, ZN => n1188);
   U1172 : OAI22_X1 port map( A1 => n5399, A2 => n3047, B1 => n3069, B2 => 
                           n3045, ZN => n1187);
   U1173 : OAI22_X1 port map( A1 => n5149, A2 => n3047, B1 => n3070, B2 => 
                           n3045, ZN => n1186);
   U1174 : OAI22_X1 port map( A1 => n5400, A2 => n3047, B1 => n3071, B2 => 
                           n3045, ZN => n1185);
   U1175 : OAI22_X1 port map( A1 => n4904, A2 => n3047, B1 => n3073, B2 => 
                           n3045, ZN => n1184);
   U1176 : OAI22_X1 port map( A1 => n4905, A2 => n3047, B1 => n3074, B2 => 
                           n3046, ZN => n1183);
   U1177 : OAI22_X1 port map( A1 => n4906, A2 => n3047, B1 => n3075, B2 => 
                           n3046, ZN => n1182);
   U1178 : OAI22_X1 port map( A1 => n5401, A2 => n3047, B1 => n3076, B2 => 
                           n3046, ZN => n1181);
   U1179 : OAI22_X1 port map( A1 => n5150, A2 => n3047, B1 => n3077, B2 => 
                           n3046, ZN => n1180);
   U1180 : OAI22_X1 port map( A1 => n5151, A2 => n3047, B1 => n3078, B2 => 
                           n3046, ZN => n1179);
   U1181 : OAI22_X1 port map( A1 => n4907, A2 => n3047, B1 => n3079, B2 => 
                           n3046, ZN => n1178);
   U1182 : OAI22_X1 port map( A1 => n4908, A2 => n3047, B1 => n3080, B2 => 
                           n3046, ZN => n1177);
   U1183 : OAI22_X1 port map( A1 => n5152, A2 => n3047, B1 => n3081, B2 => 
                           n3046, ZN => n1176);
   U1184 : OAI22_X1 port map( A1 => n5153, A2 => n3047, B1 => n3083, B2 => 
                           n3046, ZN => n1175);
   U1185 : NAND2_X1 port map( A1 => n3049, A2 => n3048, ZN => n3072);
   U1186 : CLKBUF_X1 port map( A => n3072, Z => n3082);
   U1187 : OAI22_X1 port map( A1 => n4651, A2 => n3084, B1 => n3050, B2 => 
                           n3082, ZN => n1174);
   U1188 : OAI22_X1 port map( A1 => n4909, A2 => n3084, B1 => n3051, B2 => 
                           n3072, ZN => n1173);
   U1189 : OAI22_X1 port map( A1 => n5664, A2 => n3084, B1 => n3052, B2 => 
                           n3082, ZN => n1172);
   U1190 : OAI22_X1 port map( A1 => n4910, A2 => n3084, B1 => n3053, B2 => 
                           n3072, ZN => n1171);
   U1191 : OAI22_X1 port map( A1 => n5665, A2 => n3084, B1 => n3054, B2 => 
                           n3082, ZN => n1170);
   U1192 : OAI22_X1 port map( A1 => n5154, A2 => n3084, B1 => n3055, B2 => 
                           n3072, ZN => n1169);
   U1193 : OAI22_X1 port map( A1 => n5155, A2 => n3084, B1 => n3056, B2 => 
                           n3082, ZN => n1168);
   U1194 : OAI22_X1 port map( A1 => n5402, A2 => n3084, B1 => n3057, B2 => 
                           n3072, ZN => n1167);
   U1195 : OAI22_X1 port map( A1 => n4911, A2 => n3084, B1 => n3058, B2 => 
                           n3082, ZN => n1166);
   U1196 : OAI22_X1 port map( A1 => n5666, A2 => n3084, B1 => n3059, B2 => 
                           n3072, ZN => n1165);
   U1197 : OAI22_X1 port map( A1 => n5403, A2 => n3084, B1 => n3060, B2 => 
                           n3072, ZN => n1164);
   U1198 : OAI22_X1 port map( A1 => n5667, A2 => n3084, B1 => n3061, B2 => 
                           n3082, ZN => n1163);
   U1199 : OAI22_X1 port map( A1 => n5404, A2 => n3084, B1 => n3062, B2 => 
                           n3072, ZN => n1162);
   U1200 : OAI22_X1 port map( A1 => n4912, A2 => n3084, B1 => n3063, B2 => 
                           n3082, ZN => n1161);
   U1201 : OAI22_X1 port map( A1 => n5668, A2 => n3084, B1 => n3064, B2 => 
                           n3072, ZN => n1160);
   U1202 : OAI22_X1 port map( A1 => n4913, A2 => n3084, B1 => n3065, B2 => 
                           n3082, ZN => n1159);
   U1203 : OAI22_X1 port map( A1 => n5669, A2 => n3084, B1 => n3066, B2 => 
                           n3072, ZN => n1158);
   U1204 : OAI22_X1 port map( A1 => n5156, A2 => n3084, B1 => n3067, B2 => 
                           n3072, ZN => n1157);
   U1205 : OAI22_X1 port map( A1 => n5157, A2 => n3084, B1 => n3068, B2 => 
                           n3072, ZN => n1156);
   U1206 : OAI22_X1 port map( A1 => n5670, A2 => n3084, B1 => n3069, B2 => 
                           n3072, ZN => n1155);
   U1207 : OAI22_X1 port map( A1 => n4914, A2 => n3084, B1 => n3070, B2 => 
                           n3072, ZN => n1154);
   U1208 : OAI22_X1 port map( A1 => n5671, A2 => n3084, B1 => n3071, B2 => 
                           n3072, ZN => n1153);
   U1209 : OAI22_X1 port map( A1 => n5158, A2 => n3084, B1 => n3073, B2 => 
                           n3072, ZN => n1152);
   U1210 : OAI22_X1 port map( A1 => n5405, A2 => n3084, B1 => n3074, B2 => 
                           n3082, ZN => n1151);
   U1211 : OAI22_X1 port map( A1 => n4915, A2 => n3084, B1 => n3075, B2 => 
                           n3082, ZN => n1150);
   U1212 : OAI22_X1 port map( A1 => n5159, A2 => n3084, B1 => n3076, B2 => 
                           n3082, ZN => n1149);
   U1213 : OAI22_X1 port map( A1 => n5160, A2 => n3084, B1 => n3077, B2 => 
                           n3082, ZN => n1148);
   U1214 : OAI22_X1 port map( A1 => n5161, A2 => n3084, B1 => n3078, B2 => 
                           n3082, ZN => n1147);
   U1215 : OAI22_X1 port map( A1 => n5406, A2 => n3084, B1 => n3079, B2 => 
                           n3082, ZN => n1146);
   U1216 : OAI22_X1 port map( A1 => n5162, A2 => n3084, B1 => n3080, B2 => 
                           n3082, ZN => n1145);
   U1217 : OAI22_X1 port map( A1 => n5407, A2 => n3084, B1 => n3081, B2 => 
                           n3082, ZN => n1144);
   U1218 : OAI22_X1 port map( A1 => n5163, A2 => n3084, B1 => n3083, B2 => 
                           n3082, ZN => n1143);
   U1219 : NAND3_X1 port map( A1 => n2898, A2 => ENABLE, A3 => RD2, ZN => n3866
                           );
   U1220 : INV_X1 port map( A => ADD_RD2(3), ZN => n3107);
   U1221 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n3107, ZN => n3094);
   U1222 : INV_X1 port map( A => ADD_RD2(2), ZN => n3091);
   U1223 : OR3_X1 port map( A1 => n3091, A2 => ADD_RD2(0), A3 => ADD_RD2(1), ZN
                           => n3151);
   U1224 : NOR2_X1 port map( A1 => n3094, A2 => n3151, ZN => n3588);
   U1225 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n3093);
   U1226 : INV_X1 port map( A => ADD_RD2(1), ZN => n3089);
   U1227 : OR3_X1 port map( A1 => n3091, A2 => n3089, A3 => ADD_RD2(0), ZN => 
                           n3222);
   U1228 : NOR2_X1 port map( A1 => n3093, A2 => n3222, ZN => n3831);
   U1229 : CLKBUF_X1 port map( A => n3831, Z => n3658);
   U1230 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n3588, B1 => 
                           REGISTERS_30_31_port, B2 => n3658, ZN => n3088);
   U1231 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), ZN => n3090);
   U1232 : NAND2_X1 port map( A1 => n3090, A2 => ADD_RD2(1), ZN => n3101);
   U1233 : NOR2_X1 port map( A1 => n3093, A2 => n3101, ZN => n3786);
   U1234 : INV_X1 port map( A => ADD_RD2(0), ZN => n3092);
   U1235 : OR3_X1 port map( A1 => n3091, A2 => n3092, A3 => n3089, ZN => n3126)
                           ;
   U1236 : NOR2_X1 port map( A1 => n3093, A2 => n3126, ZN => n3833);
   U1237 : CLKBUF_X1 port map( A => n3833, Z => n3787);
   U1238 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n3786, B1 => 
                           REGISTERS_31_31_port, B2 => n3787, ZN => n3087);
   U1239 : NOR2_X1 port map( A1 => n3094, A2 => n3101, ZN => n3568);
   U1240 : OR3_X1 port map( A1 => n3092, A2 => n3089, A3 => ADD_RD2(2), ZN => 
                           n3128);
   U1241 : NOR2_X1 port map( A1 => n3093, A2 => n3128, ZN => n3827);
   U1242 : AOI22_X1 port map( A1 => REGISTERS_18_31_port, A2 => n3568, B1 => 
                           REGISTERS_27_31_port, B2 => n3827, ZN => n3086);
   U1243 : OR3_X1 port map( A1 => n3092, A2 => ADD_RD2(2), A3 => ADD_RD2(1), ZN
                           => n3127);
   U1244 : NOR2_X1 port map( A1 => n3093, A2 => n3127, ZN => n3390);
   U1245 : NOR2_X1 port map( A1 => n3094, A2 => n3126, ZN => n3756);
   U1246 : CLKBUF_X1 port map( A => n3756, Z => n3817);
   U1247 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n3390, B1 => 
                           REGISTERS_23_31_port, B2 => n3817, ZN => n3085);
   U1248 : NAND4_X1 port map( A1 => n3088, A2 => n3087, A3 => n3086, A4 => 
                           n3085, ZN => n3100);
   U1249 : NAND2_X1 port map( A1 => n3090, A2 => n3089, ZN => n3102);
   U1250 : NOR2_X1 port map( A1 => n3102, A2 => n3094, ZN => n3815);
   U1251 : NOR2_X1 port map( A1 => n3093, A2 => n3151, ZN => n3659);
   U1252 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n3815, B1 => 
                           REGISTERS_28_31_port, B2 => n3659, ZN => n3098);
   U1253 : NOR2_X1 port map( A1 => n3093, A2 => n3102, ZN => n3816);
   U1254 : OR3_X1 port map( A1 => n3092, A2 => n3091, A3 => ADD_RD2(1), ZN => 
                           n3333);
   U1255 : NOR2_X1 port map( A1 => n3093, A2 => n3333, ZN => n3664);
   U1256 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n3816, B1 => 
                           REGISTERS_29_31_port, B2 => n3664, ZN => n3097);
   U1257 : NOR2_X1 port map( A1 => n3333, A2 => n3094, ZN => n3761);
   U1258 : NOR2_X1 port map( A1 => n3094, A2 => n3128, ZN => n3569);
   U1259 : CLKBUF_X1 port map( A => n3569, Z => n3832);
   U1260 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n3761, B1 => 
                           REGISTERS_19_31_port, B2 => n3832, ZN => n3096);
   U1261 : NOR2_X1 port map( A1 => n3094, A2 => n3222, ZN => n3734);
   U1262 : NOR2_X1 port map( A1 => n3094, A2 => n3127, ZN => n3821);
   U1263 : CLKBUF_X1 port map( A => n3821, Z => n3755);
   U1264 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n3734, B1 => 
                           REGISTERS_17_31_port, B2 => n3755, ZN => n3095);
   U1265 : NAND4_X1 port map( A1 => n3098, A2 => n3097, A3 => n3096, A4 => 
                           n3095, ZN => n3099);
   U1266 : NOR2_X1 port map( A1 => n3100, A2 => n3099, ZN => n3115);
   U1267 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n3814, 
                           ZN => n3863);
   U1268 : CLKBUF_X1 port map( A => n3863, Z => n3681);
   U1269 : INV_X1 port map( A => n3128, ZN => n3805);
   U1270 : INV_X1 port map( A => n3101, ZN => n3854);
   U1271 : CLKBUF_X1 port map( A => n3854, Z => n3746);
   U1272 : AOI22_X1 port map( A1 => n3805, A2 => REGISTERS_3_31_port, B1 => 
                           n3746, B2 => REGISTERS_2_31_port, ZN => n3106);
   U1273 : INV_X1 port map( A => n3222, ZN => n3855);
   U1274 : INV_X1 port map( A => n3126, ZN => n3852);
   U1275 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_31_port, B1 => 
                           n3852, B2 => REGISTERS_7_31_port, ZN => n3105);
   U1276 : INV_X1 port map( A => n3151, ZN => n3777);
   U1277 : INV_X1 port map( A => n3127, ZN => n3850);
   U1278 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_4_31_port, B1 => 
                           n3850, B2 => REGISTERS_1_31_port, ZN => n3104);
   U1279 : INV_X1 port map( A => n3102, ZN => n3769);
   U1280 : CLKBUF_X1 port map( A => n3769, Z => n3555);
   U1281 : INV_X1 port map( A => n3333, ZN => n3798);
   U1282 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_31_port, B1 => 
                           n3798, B2 => REGISTERS_5_31_port, ZN => n3103);
   U1283 : NAND4_X1 port map( A1 => n3106, A2 => n3105, A3 => n3104, A4 => 
                           n3103, ZN => n3113);
   U1284 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n3107, A3 => n3814, ZN => 
                           n3861);
   U1285 : CLKBUF_X1 port map( A => n3861, Z => n3703);
   U1286 : INV_X1 port map( A => n3126, ZN => n3775);
   U1287 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_31_port, B1 => 
                           n3775, B2 => REGISTERS_15_31_port, ZN => n3111);
   U1288 : INV_X1 port map( A => n3151, ZN => n3851);
   U1289 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_31_port, B1 => 
                           n3855, B2 => REGISTERS_14_31_port, ZN => n3110);
   U1290 : INV_X1 port map( A => n3333, ZN => n3848);
   U1291 : INV_X1 port map( A => n3127, ZN => n3774);
   U1292 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_31_port, B1 => 
                           n3774, B2 => REGISTERS_9_31_port, ZN => n3109);
   U1293 : INV_X1 port map( A => n3128, ZN => n3843);
   U1294 : AOI22_X1 port map( A1 => n3843, A2 => REGISTERS_11_31_port, B1 => 
                           n3746, B2 => REGISTERS_10_31_port, ZN => n3108);
   U1295 : NAND4_X1 port map( A1 => n3111, A2 => n3110, A3 => n3109, A4 => 
                           n3108, ZN => n3112);
   U1296 : AOI22_X1 port map( A1 => n3681, A2 => n3113, B1 => n3703, B2 => 
                           n3112, ZN => n3114);
   U1297 : OAI21_X1 port map( B1 => n3814, B2 => n3115, A => n3114, ZN => N448)
                           ;
   U1298 : CLKBUF_X1 port map( A => n3588, Z => n3818);
   U1299 : AOI22_X1 port map( A1 => n3659, A2 => REGISTERS_28_30_port, B1 => 
                           n3818, B2 => REGISTERS_20_30_port, ZN => n3119);
   U1300 : CLKBUF_X1 port map( A => n3815, Z => n3762);
   U1301 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_30_port, B1 => 
                           n3833, B2 => REGISTERS_31_30_port, ZN => n3118);
   U1302 : CLKBUF_X1 port map( A => n3734, Z => n3822);
   U1303 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_30_port, B1 => 
                           n3832, B2 => REGISTERS_19_30_port, ZN => n3117);
   U1304 : CLKBUF_X1 port map( A => n3761, Z => n3828);
   U1305 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_30_port, B1 => 
                           n3831, B2 => REGISTERS_30_30_port, ZN => n3116);
   U1306 : NAND4_X1 port map( A1 => n3119, A2 => n3118, A3 => n3117, A4 => 
                           n3116, ZN => n3125);
   U1307 : CLKBUF_X1 port map( A => n3786, Z => n3830);
   U1308 : CLKBUF_X1 port map( A => n3827, Z => n3616);
   U1309 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_30_port, B1 => 
                           n3616, B2 => REGISTERS_27_30_port, ZN => n3123);
   U1310 : CLKBUF_X1 port map( A => n3390, Z => n3819);
   U1311 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_30_port, B1 => 
                           n3819, B2 => REGISTERS_25_30_port, ZN => n3122);
   U1312 : CLKBUF_X1 port map( A => n3816, Z => n3611);
   U1313 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_30_port, B1 => 
                           n3817, B2 => REGISTERS_23_30_port, ZN => n3121);
   U1314 : CLKBUF_X1 port map( A => n3568, Z => n3829);
   U1315 : AOI22_X1 port map( A1 => n3664, A2 => REGISTERS_29_30_port, B1 => 
                           n3829, B2 => REGISTERS_18_30_port, ZN => n3120);
   U1316 : NAND4_X1 port map( A1 => n3123, A2 => n3122, A3 => n3121, A4 => 
                           n3120, ZN => n3124);
   U1317 : NOR2_X1 port map( A1 => n3125, A2 => n3124, ZN => n3140);
   U1318 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_5_30_port, B1 => 
                           n3855, B2 => REGISTERS_6_30_port, ZN => n3132);
   U1319 : CLKBUF_X1 port map( A => n3854, Z => n3842);
   U1320 : INV_X1 port map( A => n3126, ZN => n3627);
   U1321 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_30_port, B1 => 
                           n3627, B2 => REGISTERS_7_30_port, ZN => n3131);
   U1322 : INV_X1 port map( A => n3127, ZN => n3741);
   U1323 : INV_X1 port map( A => n3128, ZN => n3853);
   U1324 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_1_30_port, B1 => 
                           n3853, B2 => REGISTERS_3_30_port, ZN => n3130);
   U1325 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_30_port, B1 => 
                           n3851, B2 => REGISTERS_4_30_port, ZN => n3129);
   U1326 : NAND4_X1 port map( A1 => n3132, A2 => n3131, A3 => n3130, A4 => 
                           n3129, ZN => n3138);
   U1327 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_30_port, B1 => 
                           n3746, B2 => REGISTERS_10_30_port, ZN => n3136);
   U1328 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_9_30_port, B1 => 
                           n3843, B2 => REGISTERS_11_30_port, ZN => n3135);
   U1329 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_30_port, B1 => 
                           n3851, B2 => REGISTERS_12_30_port, ZN => n3134);
   U1330 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_30_port, B1 => 
                           n3852, B2 => REGISTERS_15_30_port, ZN => n3133);
   U1331 : NAND4_X1 port map( A1 => n3136, A2 => n3135, A3 => n3134, A4 => 
                           n3133, ZN => n3137);
   U1332 : AOI22_X1 port map( A1 => n3681, A2 => n3138, B1 => n3703, B2 => 
                           n3137, ZN => n3139);
   U1333 : OAI21_X1 port map( B1 => n3814, B2 => n3140, A => n3139, ZN => N447)
                           ;
   U1334 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_29_port, B1 => 
                           n3568, B2 => REGISTERS_18_29_port, ZN => n3144);
   U1335 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_29_port, B1 => 
                           n3390, B2 => REGISTERS_25_29_port, ZN => n3143);
   U1336 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_29_port, B1 => 
                           n3658, B2 => REGISTERS_30_29_port, ZN => n3142);
   U1337 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_29_port, B1 => 
                           n3588, B2 => REGISTERS_20_29_port, ZN => n3141);
   U1338 : NAND4_X1 port map( A1 => n3144, A2 => n3143, A3 => n3142, A4 => 
                           n3141, ZN => n3150);
   U1339 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_29_port, B1 => 
                           n3664, B2 => REGISTERS_29_29_port, ZN => n3148);
   U1340 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_29_port, B1 => 
                           n3616, B2 => REGISTERS_27_29_port, ZN => n3147);
   U1341 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_29_port, B1 => 
                           n3786, B2 => REGISTERS_26_29_port, ZN => n3146);
   U1342 : AOI22_X1 port map( A1 => n3659, A2 => REGISTERS_28_29_port, B1 => 
                           n3756, B2 => REGISTERS_23_29_port, ZN => n3145);
   U1343 : NAND4_X1 port map( A1 => n3148, A2 => n3147, A3 => n3146, A4 => 
                           n3145, ZN => n3149);
   U1344 : NOR2_X1 port map( A1 => n3150, A2 => n3149, ZN => n3163);
   U1345 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_29_port, B1 => 
                           n3843, B2 => REGISTERS_3_29_port, ZN => n3155);
   U1346 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_29_port, B1 => 
                           n3798, B2 => REGISTERS_5_29_port, ZN => n3154);
   U1347 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_29_port, B1 => 
                           n3746, B2 => REGISTERS_2_29_port, ZN => n3153);
   U1348 : INV_X1 port map( A => n3151, ZN => n3841);
   U1349 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_29_port, B1 => 
                           n3775, B2 => REGISTERS_7_29_port, ZN => n3152);
   U1350 : NAND4_X1 port map( A1 => n3155, A2 => n3154, A3 => n3153, A4 => 
                           n3152, ZN => n3161);
   U1351 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_29_port, B1 => 
                           n3627, B2 => REGISTERS_15_29_port, ZN => n3159);
   U1352 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_29_port, B1 => 
                           n3843, B2 => REGISTERS_11_29_port, ZN => n3158);
   U1353 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_29_port, B1 => 
                           n3746, B2 => REGISTERS_10_29_port, ZN => n3157);
   U1354 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_29_port, B1 => 
                           n3774, B2 => REGISTERS_9_29_port, ZN => n3156);
   U1355 : NAND4_X1 port map( A1 => n3159, A2 => n3158, A3 => n3157, A4 => 
                           n3156, ZN => n3160);
   U1356 : AOI22_X1 port map( A1 => n3681, A2 => n3161, B1 => n3703, B2 => 
                           n3160, ZN => n3162);
   U1357 : OAI21_X1 port map( B1 => n3814, B2 => n3163, A => n3162, ZN => N446)
                           ;
   U1358 : AOI22_X1 port map( A1 => n3734, A2 => REGISTERS_22_28_port, B1 => 
                           n3821, B2 => REGISTERS_17_28_port, ZN => n3167);
   U1359 : CLKBUF_X1 port map( A => n3659, Z => n3834);
   U1360 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_28_port, B1 => 
                           n3569, B2 => REGISTERS_19_28_port, ZN => n3166);
   U1361 : AOI22_X1 port map( A1 => n3664, A2 => REGISTERS_29_28_port, B1 => 
                           n3786, B2 => REGISTERS_26_28_port, ZN => n3165);
   U1362 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_28_port, B1 => 
                           n3390, B2 => REGISTERS_25_28_port, ZN => n3164);
   U1363 : NAND4_X1 port map( A1 => n3167, A2 => n3166, A3 => n3165, A4 => 
                           n3164, ZN => n3173);
   U1364 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_28_port, B1 => 
                           n3756, B2 => REGISTERS_23_28_port, ZN => n3171);
   U1365 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_28_port, B1 => 
                           n3616, B2 => REGISTERS_27_28_port, ZN => n3170);
   U1366 : AOI22_X1 port map( A1 => n3815, A2 => REGISTERS_16_28_port, B1 => 
                           n3833, B2 => REGISTERS_31_28_port, ZN => n3169);
   U1367 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_28_port, B1 => 
                           n3568, B2 => REGISTERS_18_28_port, ZN => n3168);
   U1368 : NAND4_X1 port map( A1 => n3171, A2 => n3170, A3 => n3169, A4 => 
                           n3168, ZN => n3172);
   U1369 : NOR2_X1 port map( A1 => n3173, A2 => n3172, ZN => n3185);
   U1370 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_28_port, B1 => 
                           n3843, B2 => REGISTERS_3_28_port, ZN => n3177);
   U1371 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_28_port, B1 => 
                           n3774, B2 => REGISTERS_1_28_port, ZN => n3176);
   U1372 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_28_port, B1 => 
                           n3848, B2 => REGISTERS_5_28_port, ZN => n3175);
   U1373 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_28_port, B1 => 
                           n3852, B2 => REGISTERS_7_28_port, ZN => n3174);
   U1374 : NAND4_X1 port map( A1 => n3177, A2 => n3176, A3 => n3175, A4 => 
                           n3174, ZN => n3183);
   U1375 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_28_port, B1 => 
                           n3775, B2 => REGISTERS_15_28_port, ZN => n3181);
   U1376 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_28_port, B1 => 
                           n3774, B2 => REGISTERS_9_28_port, ZN => n3180);
   U1377 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_28_port, B1 => 
                           n3853, B2 => REGISTERS_11_28_port, ZN => n3179);
   U1378 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_28_port, B1 => 
                           n3746, B2 => REGISTERS_10_28_port, ZN => n3178);
   U1379 : NAND4_X1 port map( A1 => n3181, A2 => n3180, A3 => n3179, A4 => 
                           n3178, ZN => n3182);
   U1380 : AOI22_X1 port map( A1 => n3681, A2 => n3183, B1 => n3703, B2 => 
                           n3182, ZN => n3184);
   U1381 : OAI21_X1 port map( B1 => n3814, B2 => n3185, A => n3184, ZN => N445)
                           ;
   U1382 : AOI22_X1 port map( A1 => n3664, A2 => REGISTERS_29_27_port, B1 => 
                           n3756, B2 => REGISTERS_23_27_port, ZN => n3189);
   U1383 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_27_port, B1 => 
                           n3390, B2 => REGISTERS_25_27_port, ZN => n3188);
   U1384 : AOI22_X1 port map( A1 => n3815, A2 => REGISTERS_16_27_port, B1 => 
                           n3786, B2 => REGISTERS_26_27_port, ZN => n3187);
   U1385 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_27_port, B1 => 
                           n3658, B2 => REGISTERS_30_27_port, ZN => n3186);
   U1386 : NAND4_X1 port map( A1 => n3189, A2 => n3188, A3 => n3187, A4 => 
                           n3186, ZN => n3195);
   U1387 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_27_port, B1 => 
                           n3616, B2 => REGISTERS_27_27_port, ZN => n3193);
   U1388 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_27_port, B1 => 
                           n3568, B2 => REGISTERS_18_27_port, ZN => n3192);
   U1389 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_27_port, B1 => 
                           n3569, B2 => REGISTERS_19_27_port, ZN => n3191);
   U1390 : AOI22_X1 port map( A1 => n3659, A2 => REGISTERS_28_27_port, B1 => 
                           n3821, B2 => REGISTERS_17_27_port, ZN => n3190);
   U1391 : NAND4_X1 port map( A1 => n3193, A2 => n3192, A3 => n3191, A4 => 
                           n3190, ZN => n3194);
   U1392 : NOR2_X1 port map( A1 => n3195, A2 => n3194, ZN => n3207);
   U1393 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_27_port, B1 => 
                           n3627, B2 => REGISTERS_7_27_port, ZN => n3199);
   U1394 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_5_27_port, B1 => 
                           n3853, B2 => REGISTERS_3_27_port, ZN => n3198);
   U1395 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_27_port, B1 => 
                           n3741, B2 => REGISTERS_1_27_port, ZN => n3197);
   U1396 : INV_X1 port map( A => n3222, ZN => n3799);
   U1397 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_27_port, B1 => 
                           n3799, B2 => REGISTERS_6_27_port, ZN => n3196);
   U1398 : NAND4_X1 port map( A1 => n3199, A2 => n3198, A3 => n3197, A4 => 
                           n3196, ZN => n3205);
   U1399 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_27_port, B1 => 
                           n3853, B2 => REGISTERS_11_27_port, ZN => n3203);
   U1400 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_27_port, B1 => 
                           n3741, B2 => REGISTERS_9_27_port, ZN => n3202);
   U1401 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_27_port, B1 => 
                           n3799, B2 => REGISTERS_14_27_port, ZN => n3201);
   U1402 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_10_27_port, B1 => 
                           n3852, B2 => REGISTERS_15_27_port, ZN => n3200);
   U1403 : NAND4_X1 port map( A1 => n3203, A2 => n3202, A3 => n3201, A4 => 
                           n3200, ZN => n3204);
   U1404 : AOI22_X1 port map( A1 => n3681, A2 => n3205, B1 => n3703, B2 => 
                           n3204, ZN => n3206);
   U1405 : OAI21_X1 port map( B1 => n3814, B2 => n3207, A => n3206, ZN => N444)
                           ;
   U1406 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_26_port, B1 => 
                           n3658, B2 => REGISTERS_30_26_port, ZN => n3211);
   U1407 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_26_port, B1 => 
                           n3756, B2 => REGISTERS_23_26_port, ZN => n3210);
   U1408 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_26_port, B1 => 
                           n3568, B2 => REGISTERS_18_26_port, ZN => n3209);
   U1409 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_26_port, B1 => 
                           n3390, B2 => REGISTERS_25_26_port, ZN => n3208);
   U1410 : NAND4_X1 port map( A1 => n3211, A2 => n3210, A3 => n3209, A4 => 
                           n3208, ZN => n3217);
   U1411 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_26_port, B1 => 
                           n3664, B2 => REGISTERS_29_26_port, ZN => n3215);
   U1412 : AOI22_X1 port map( A1 => n3659, A2 => REGISTERS_28_26_port, B1 => 
                           n3787, B2 => REGISTERS_31_26_port, ZN => n3214);
   U1413 : AOI22_X1 port map( A1 => n3815, A2 => REGISTERS_16_26_port, B1 => 
                           n3588, B2 => REGISTERS_20_26_port, ZN => n3213);
   U1414 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_26_port, B1 => 
                           n3616, B2 => REGISTERS_27_26_port, ZN => n3212);
   U1415 : NAND4_X1 port map( A1 => n3215, A2 => n3214, A3 => n3213, A4 => 
                           n3212, ZN => n3216);
   U1416 : NOR2_X1 port map( A1 => n3217, A2 => n3216, ZN => n3230);
   U1417 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_26_port, B1 => 
                           n3853, B2 => REGISTERS_3_26_port, ZN => n3221);
   U1418 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_26_port, B1 => 
                           n3775, B2 => REGISTERS_7_26_port, ZN => n3220);
   U1419 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_5_26_port, B1 => 
                           n3799, B2 => REGISTERS_6_26_port, ZN => n3219);
   U1420 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_26_port, B1 => 
                           n3854, B2 => REGISTERS_2_26_port, ZN => n3218);
   U1421 : NAND4_X1 port map( A1 => n3221, A2 => n3220, A3 => n3219, A4 => 
                           n3218, ZN => n3228);
   U1422 : AOI22_X1 port map( A1 => n3853, A2 => REGISTERS_11_26_port, B1 => 
                           n3627, B2 => REGISTERS_15_26_port, ZN => n3226);
   U1423 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_26_port, B1 => 
                           n3746, B2 => REGISTERS_10_26_port, ZN => n3225);
   U1424 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_26_port, B1 => 
                           n3741, B2 => REGISTERS_9_26_port, ZN => n3224);
   U1425 : INV_X1 port map( A => n3222, ZN => n3776);
   U1426 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_26_port, B1 => 
                           n3776, B2 => REGISTERS_14_26_port, ZN => n3223);
   U1427 : NAND4_X1 port map( A1 => n3226, A2 => n3225, A3 => n3224, A4 => 
                           n3223, ZN => n3227);
   U1428 : AOI22_X1 port map( A1 => n3681, A2 => n3228, B1 => n3703, B2 => 
                           n3227, ZN => n3229);
   U1429 : OAI21_X1 port map( B1 => n3814, B2 => n3230, A => n3229, ZN => N443)
                           ;
   U1430 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_25_port, B1 => 
                           n3588, B2 => REGISTERS_20_25_port, ZN => n3234);
   U1431 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_25_port, B1 => 
                           n3568, B2 => REGISTERS_18_25_port, ZN => n3233);
   U1432 : AOI22_X1 port map( A1 => n3664, A2 => REGISTERS_29_25_port, B1 => 
                           n3756, B2 => REGISTERS_23_25_port, ZN => n3232);
   U1433 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_25_port, B1 => 
                           n3390, B2 => REGISTERS_25_25_port, ZN => n3231);
   U1434 : NAND4_X1 port map( A1 => n3234, A2 => n3233, A3 => n3232, A4 => 
                           n3231, ZN => n3240);
   U1435 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_25_port, B1 => 
                           n3569, B2 => REGISTERS_19_25_port, ZN => n3238);
   U1436 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_25_port, B1 => 
                           n3787, B2 => REGISTERS_31_25_port, ZN => n3237);
   U1437 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_25_port, B1 => 
                           n3616, B2 => REGISTERS_27_25_port, ZN => n3236);
   U1438 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_25_port, B1 => 
                           n3786, B2 => REGISTERS_26_25_port, ZN => n3235);
   U1439 : NAND4_X1 port map( A1 => n3238, A2 => n3237, A3 => n3236, A4 => 
                           n3235, ZN => n3239);
   U1440 : NOR2_X1 port map( A1 => n3240, A2 => n3239, ZN => n3252);
   U1441 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_25_port, B1 => 
                           n3854, B2 => REGISTERS_2_25_port, ZN => n3244);
   U1442 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_1_25_port, B1 => 
                           n3852, B2 => REGISTERS_7_25_port, ZN => n3243);
   U1443 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_25_port, B1 => 
                           n3853, B2 => REGISTERS_3_25_port, ZN => n3242);
   U1444 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_25_port, B1 => 
                           n3798, B2 => REGISTERS_5_25_port, ZN => n3241);
   U1445 : NAND4_X1 port map( A1 => n3244, A2 => n3243, A3 => n3242, A4 => 
                           n3241, ZN => n3250);
   U1446 : CLKBUF_X1 port map( A => n3769, Z => n3849);
   U1447 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_25_port, B1 => 
                           n3853, B2 => REGISTERS_11_25_port, ZN => n3248);
   U1448 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_14_25_port, B1 => 
                           n3775, B2 => REGISTERS_15_25_port, ZN => n3247);
   U1449 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_25_port, B1 => 
                           n3741, B2 => REGISTERS_9_25_port, ZN => n3246);
   U1450 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_25_port, B1 => 
                           n3746, B2 => REGISTERS_10_25_port, ZN => n3245);
   U1451 : NAND4_X1 port map( A1 => n3248, A2 => n3247, A3 => n3246, A4 => 
                           n3245, ZN => n3249);
   U1452 : AOI22_X1 port map( A1 => n3681, A2 => n3250, B1 => n3703, B2 => 
                           n3249, ZN => n3251);
   U1453 : OAI21_X1 port map( B1 => n3814, B2 => n3252, A => n3251, ZN => N442)
                           ;
   U1454 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_24_port, B1 => 
                           n3756, B2 => REGISTERS_23_24_port, ZN => n3256);
   U1455 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_24_port, B1 => 
                           n3390, B2 => REGISTERS_25_24_port, ZN => n3255);
   U1456 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_24_port, B1 => 
                           n3830, B2 => REGISTERS_26_24_port, ZN => n3254);
   U1457 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_24_port, B1 => 
                           n3569, B2 => REGISTERS_19_24_port, ZN => n3253);
   U1458 : NAND4_X1 port map( A1 => n3256, A2 => n3255, A3 => n3254, A4 => 
                           n3253, ZN => n3262);
   U1459 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_24_port, B1 => 
                           n3616, B2 => REGISTERS_27_24_port, ZN => n3260);
   U1460 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_24_port, B1 => 
                           n3588, B2 => REGISTERS_20_24_port, ZN => n3259);
   U1461 : CLKBUF_X1 port map( A => n3664, Z => n3820);
   U1462 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_24_port, B1 => 
                           n3658, B2 => REGISTERS_30_24_port, ZN => n3258);
   U1463 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_24_port, B1 => 
                           n3568, B2 => REGISTERS_18_24_port, ZN => n3257);
   U1464 : NAND4_X1 port map( A1 => n3260, A2 => n3259, A3 => n3258, A4 => 
                           n3257, ZN => n3261);
   U1465 : NOR2_X1 port map( A1 => n3262, A2 => n3261, ZN => n3274);
   U1466 : AOI22_X1 port map( A1 => n3805, A2 => REGISTERS_3_24_port, B1 => 
                           n3627, B2 => REGISTERS_7_24_port, ZN => n3266);
   U1467 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_24_port, B1 => 
                           n3741, B2 => REGISTERS_1_24_port, ZN => n3265);
   U1468 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_24_port, B1 => 
                           n3776, B2 => REGISTERS_6_24_port, ZN => n3264);
   U1469 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_24_port, B1 => 
                           n3854, B2 => REGISTERS_2_24_port, ZN => n3263);
   U1470 : NAND4_X1 port map( A1 => n3266, A2 => n3265, A3 => n3264, A4 => 
                           n3263, ZN => n3272);
   U1471 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_24_port, B1 => 
                           n3741, B2 => REGISTERS_9_24_port, ZN => n3270);
   U1472 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_24_port, B1 => 
                           n3853, B2 => REGISTERS_11_24_port, ZN => n3269);
   U1473 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_24_port, B1 => 
                           n3746, B2 => REGISTERS_10_24_port, ZN => n3268);
   U1474 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_24_port, B1 => 
                           n3852, B2 => REGISTERS_15_24_port, ZN => n3267);
   U1475 : NAND4_X1 port map( A1 => n3270, A2 => n3269, A3 => n3268, A4 => 
                           n3267, ZN => n3271);
   U1476 : AOI22_X1 port map( A1 => n3681, A2 => n3272, B1 => n3703, B2 => 
                           n3271, ZN => n3273);
   U1477 : OAI21_X1 port map( B1 => n3814, B2 => n3274, A => n3273, ZN => N441)
                           ;
   U1478 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_23_port, B1 => 
                           n3568, B2 => REGISTERS_18_23_port, ZN => n3278);
   U1479 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_23_port, B1 => 
                           n3815, B2 => REGISTERS_16_23_port, ZN => n3277);
   U1480 : AOI22_X1 port map( A1 => n3831, A2 => REGISTERS_30_23_port, B1 => 
                           n3616, B2 => REGISTERS_27_23_port, ZN => n3276);
   U1481 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_23_port, B1 => 
                           n3787, B2 => REGISTERS_31_23_port, ZN => n3275);
   U1482 : NAND4_X1 port map( A1 => n3278, A2 => n3277, A3 => n3276, A4 => 
                           n3275, ZN => n3284);
   U1483 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_23_port, B1 => 
                           n3390, B2 => REGISTERS_25_23_port, ZN => n3282);
   U1484 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_23_port, B1 => 
                           n3569, B2 => REGISTERS_19_23_port, ZN => n3281);
   U1485 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_23_port, B1 => 
                           n3756, B2 => REGISTERS_23_23_port, ZN => n3280);
   U1486 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_23_port, B1 => 
                           n3734, B2 => REGISTERS_22_23_port, ZN => n3279);
   U1487 : NAND4_X1 port map( A1 => n3282, A2 => n3281, A3 => n3280, A4 => 
                           n3279, ZN => n3283);
   U1488 : NOR2_X1 port map( A1 => n3284, A2 => n3283, ZN => n3296);
   U1489 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_1_23_port, B1 => 
                           n3775, B2 => REGISTERS_7_23_port, ZN => n3288);
   U1490 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_0_23_port, B1 => 
                           n3854, B2 => REGISTERS_2_23_port, ZN => n3287);
   U1491 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_23_port, B1 => 
                           n3853, B2 => REGISTERS_3_23_port, ZN => n3286);
   U1492 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_23_port, B1 => 
                           n3776, B2 => REGISTERS_6_23_port, ZN => n3285);
   U1493 : NAND4_X1 port map( A1 => n3288, A2 => n3287, A3 => n3286, A4 => 
                           n3285, ZN => n3294);
   U1494 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_23_port, B1 => 
                           n3776, B2 => REGISTERS_14_23_port, ZN => n3292);
   U1495 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_8_23_port, B1 => 
                           n3853, B2 => REGISTERS_11_23_port, ZN => n3291);
   U1496 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_23_port, B1 => 
                           n3741, B2 => REGISTERS_9_23_port, ZN => n3290);
   U1497 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_10_23_port, B1 => 
                           n3775, B2 => REGISTERS_15_23_port, ZN => n3289);
   U1498 : NAND4_X1 port map( A1 => n3292, A2 => n3291, A3 => n3290, A4 => 
                           n3289, ZN => n3293);
   U1499 : AOI22_X1 port map( A1 => n3681, A2 => n3294, B1 => n3703, B2 => 
                           n3293, ZN => n3295);
   U1500 : OAI21_X1 port map( B1 => n3866, B2 => n3296, A => n3295, ZN => N440)
                           ;
   U1501 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_22_port, B1 => 
                           n3658, B2 => REGISTERS_30_22_port, ZN => n3300);
   U1502 : AOI22_X1 port map( A1 => n3786, A2 => REGISTERS_26_22_port, B1 => 
                           n3616, B2 => REGISTERS_27_22_port, ZN => n3299);
   U1503 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_22_port, B1 => 
                           n3821, B2 => REGISTERS_17_22_port, ZN => n3298);
   U1504 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_22_port, B1 => 
                           n3568, B2 => REGISTERS_18_22_port, ZN => n3297);
   U1505 : NAND4_X1 port map( A1 => n3300, A2 => n3299, A3 => n3298, A4 => 
                           n3297, ZN => n3306);
   U1506 : AOI22_X1 port map( A1 => n3833, A2 => REGISTERS_31_22_port, B1 => 
                           n3390, B2 => REGISTERS_25_22_port, ZN => n3304);
   U1507 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_22_port, B1 => 
                           n3761, B2 => REGISTERS_21_22_port, ZN => n3303);
   U1508 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_22_port, B1 => 
                           n3756, B2 => REGISTERS_23_22_port, ZN => n3302);
   U1509 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_22_port, B1 => 
                           n3569, B2 => REGISTERS_19_22_port, ZN => n3301);
   U1510 : NAND4_X1 port map( A1 => n3304, A2 => n3303, A3 => n3302, A4 => 
                           n3301, ZN => n3305);
   U1511 : NOR2_X1 port map( A1 => n3306, A2 => n3305, ZN => n3318);
   U1512 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_22_port, B1 => 
                           n3741, B2 => REGISTERS_1_22_port, ZN => n3310);
   U1513 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_22_port, B1 => 
                           n3776, B2 => REGISTERS_6_22_port, ZN => n3309);
   U1514 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_22_port, B1 => 
                           n3853, B2 => REGISTERS_3_22_port, ZN => n3308);
   U1515 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_22_port, B1 => 
                           n3627, B2 => REGISTERS_7_22_port, ZN => n3307);
   U1516 : NAND4_X1 port map( A1 => n3310, A2 => n3309, A3 => n3308, A4 => 
                           n3307, ZN => n3316);
   U1517 : AOI22_X1 port map( A1 => n3843, A2 => REGISTERS_11_22_port, B1 => 
                           n3852, B2 => REGISTERS_15_22_port, ZN => n3314);
   U1518 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_22_port, B1 => 
                           n3777, B2 => REGISTERS_12_22_port, ZN => n3313);
   U1519 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_9_22_port, B1 => 
                           n3746, B2 => REGISTERS_10_22_port, ZN => n3312);
   U1520 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_22_port, B1 => 
                           n3776, B2 => REGISTERS_14_22_port, ZN => n3311);
   U1521 : NAND4_X1 port map( A1 => n3314, A2 => n3313, A3 => n3312, A4 => 
                           n3311, ZN => n3315);
   U1522 : AOI22_X1 port map( A1 => n3681, A2 => n3316, B1 => n3703, B2 => 
                           n3315, ZN => n3317);
   U1523 : OAI21_X1 port map( B1 => n3866, B2 => n3318, A => n3317, ZN => N439)
                           ;
   U1524 : AOI22_X1 port map( A1 => n3819, A2 => REGISTERS_25_21_port, B1 => 
                           n3829, B2 => REGISTERS_18_21_port, ZN => n3322);
   U1525 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_21_port, B1 => 
                           n3827, B2 => REGISTERS_27_21_port, ZN => n3321);
   U1526 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_21_port, B1 => 
                           n3821, B2 => REGISTERS_17_21_port, ZN => n3320);
   U1527 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_21_port, B1 => 
                           n3588, B2 => REGISTERS_20_21_port, ZN => n3319);
   U1528 : NAND4_X1 port map( A1 => n3322, A2 => n3321, A3 => n3320, A4 => 
                           n3319, ZN => n3328);
   U1529 : AOI22_X1 port map( A1 => n3833, A2 => REGISTERS_31_21_port, B1 => 
                           n3658, B2 => REGISTERS_30_21_port, ZN => n3326);
   U1530 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_21_port, B1 => 
                           n3569, B2 => REGISTERS_19_21_port, ZN => n3325);
   U1531 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_21_port, B1 => 
                           n3817, B2 => REGISTERS_23_21_port, ZN => n3324);
   U1532 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_21_port, B1 => 
                           n3734, B2 => REGISTERS_22_21_port, ZN => n3323);
   U1533 : NAND4_X1 port map( A1 => n3326, A2 => n3325, A3 => n3324, A4 => 
                           n3323, ZN => n3327);
   U1534 : NOR2_X1 port map( A1 => n3328, A2 => n3327, ZN => n3341);
   U1535 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_21_port, B1 => 
                           n3854, B2 => REGISTERS_2_21_port, ZN => n3332);
   U1536 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_21_port, B1 => 
                           n3627, B2 => REGISTERS_7_21_port, ZN => n3331);
   U1537 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_21_port, B1 => 
                           n3841, B2 => REGISTERS_4_21_port, ZN => n3330);
   U1538 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_21_port, B1 => 
                           n3853, B2 => REGISTERS_3_21_port, ZN => n3329);
   U1539 : NAND4_X1 port map( A1 => n3332, A2 => n3331, A3 => n3330, A4 => 
                           n3329, ZN => n3339);
   U1540 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_21_port, B1 => 
                           n3776, B2 => REGISTERS_14_21_port, ZN => n3337);
   U1541 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_9_21_port, B1 => 
                           n3746, B2 => REGISTERS_10_21_port, ZN => n3336);
   U1542 : INV_X1 port map( A => n3333, ZN => n3804);
   U1543 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_21_port, B1 => 
                           n3775, B2 => REGISTERS_15_21_port, ZN => n3335);
   U1544 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_21_port, B1 => 
                           n3853, B2 => REGISTERS_11_21_port, ZN => n3334);
   U1545 : NAND4_X1 port map( A1 => n3337, A2 => n3336, A3 => n3335, A4 => 
                           n3334, ZN => n3338);
   U1546 : AOI22_X1 port map( A1 => n3681, A2 => n3339, B1 => n3703, B2 => 
                           n3338, ZN => n3340);
   U1547 : OAI21_X1 port map( B1 => n3866, B2 => n3341, A => n3340, ZN => N438)
                           ;
   U1548 : AOI22_X1 port map( A1 => n3831, A2 => REGISTERS_30_20_port, B1 => 
                           n3819, B2 => REGISTERS_25_20_port, ZN => n3345);
   U1549 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_20_port, B1 => 
                           n3588, B2 => REGISTERS_20_20_port, ZN => n3344);
   U1550 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_20_port, B1 => 
                           n3761, B2 => REGISTERS_21_20_port, ZN => n3343);
   U1551 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_20_port, B1 => 
                           n3830, B2 => REGISTERS_26_20_port, ZN => n3342);
   U1552 : NAND4_X1 port map( A1 => n3345, A2 => n3344, A3 => n3343, A4 => 
                           n3342, ZN => n3351);
   U1553 : AOI22_X1 port map( A1 => n3833, A2 => REGISTERS_31_20_port, B1 => 
                           n3829, B2 => REGISTERS_18_20_port, ZN => n3349);
   U1554 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_20_port, B1 => 
                           n3827, B2 => REGISTERS_27_20_port, ZN => n3348);
   U1555 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_20_port, B1 => 
                           n3821, B2 => REGISTERS_17_20_port, ZN => n3347);
   U1556 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_20_port, B1 => 
                           n3817, B2 => REGISTERS_23_20_port, ZN => n3346);
   U1557 : NAND4_X1 port map( A1 => n3349, A2 => n3348, A3 => n3347, A4 => 
                           n3346, ZN => n3350);
   U1558 : NOR2_X1 port map( A1 => n3351, A2 => n3350, ZN => n3363);
   U1559 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_0_20_port, B1 => 
                           n3776, B2 => REGISTERS_6_20_port, ZN => n3355);
   U1560 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_5_20_port, B1 => 
                           n3627, B2 => REGISTERS_7_20_port, ZN => n3354);
   U1561 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_20_port, B1 => 
                           n3854, B2 => REGISTERS_2_20_port, ZN => n3353);
   U1562 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_20_port, B1 => 
                           n3805, B2 => REGISTERS_3_20_port, ZN => n3352);
   U1563 : NAND4_X1 port map( A1 => n3355, A2 => n3354, A3 => n3353, A4 => 
                           n3352, ZN => n3361);
   U1564 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_9_20_port, B1 => 
                           n3852, B2 => REGISTERS_15_20_port, ZN => n3359);
   U1565 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_8_20_port, B1 => 
                           n3777, B2 => REGISTERS_12_20_port, ZN => n3358);
   U1566 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_20_port, B1 => 
                           n3805, B2 => REGISTERS_11_20_port, ZN => n3357);
   U1567 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_20_port, B1 => 
                           n3854, B2 => REGISTERS_10_20_port, ZN => n3356);
   U1568 : NAND4_X1 port map( A1 => n3359, A2 => n3358, A3 => n3357, A4 => 
                           n3356, ZN => n3360);
   U1569 : AOI22_X1 port map( A1 => n3681, A2 => n3361, B1 => n3861, B2 => 
                           n3360, ZN => n3362);
   U1570 : OAI21_X1 port map( B1 => n3866, B2 => n3363, A => n3362, ZN => N437)
                           ;
   U1571 : AOI22_X1 port map( A1 => n3831, A2 => REGISTERS_30_19_port, B1 => 
                           n3616, B2 => REGISTERS_27_19_port, ZN => n3367);
   U1572 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_19_port, B1 => 
                           n3829, B2 => REGISTERS_18_19_port, ZN => n3366);
   U1573 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_19_port, B1 => 
                           n3588, B2 => REGISTERS_20_19_port, ZN => n3365);
   U1574 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_19_port, B1 => 
                           n3815, B2 => REGISTERS_16_19_port, ZN => n3364);
   U1575 : NAND4_X1 port map( A1 => n3367, A2 => n3366, A3 => n3365, A4 => 
                           n3364, ZN => n3373);
   U1576 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_19_port, B1 => 
                           n3830, B2 => REGISTERS_26_19_port, ZN => n3371);
   U1577 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_19_port, B1 => 
                           n3755, B2 => REGISTERS_17_19_port, ZN => n3370);
   U1578 : AOI22_X1 port map( A1 => n3390, A2 => REGISTERS_25_19_port, B1 => 
                           n3817, B2 => REGISTERS_23_19_port, ZN => n3369);
   U1579 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_19_port, B1 => 
                           n3569, B2 => REGISTERS_19_19_port, ZN => n3368);
   U1580 : NAND4_X1 port map( A1 => n3371, A2 => n3370, A3 => n3369, A4 => 
                           n3368, ZN => n3372);
   U1581 : NOR2_X1 port map( A1 => n3373, A2 => n3372, ZN => n3385);
   U1582 : CLKBUF_X1 port map( A => n3863, Z => n3705);
   U1583 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_4_19_port, B1 => 
                           n3852, B2 => REGISTERS_7_19_port, ZN => n3377);
   U1584 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_19_port, B1 => 
                           n3746, B2 => REGISTERS_2_19_port, ZN => n3376);
   U1585 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_19_port, B1 => 
                           n3855, B2 => REGISTERS_6_19_port, ZN => n3375);
   U1586 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_1_19_port, B1 => 
                           n3805, B2 => REGISTERS_3_19_port, ZN => n3374);
   U1587 : NAND4_X1 port map( A1 => n3377, A2 => n3376, A3 => n3375, A4 => 
                           n3374, ZN => n3383);
   U1588 : AOI22_X1 port map( A1 => n3853, A2 => REGISTERS_11_19_port, B1 => 
                           n3775, B2 => REGISTERS_15_19_port, ZN => n3381);
   U1589 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_14_19_port, B1 => 
                           n3741, B2 => REGISTERS_9_19_port, ZN => n3380);
   U1590 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_19_port, B1 => 
                           n3777, B2 => REGISTERS_12_19_port, ZN => n3379);
   U1591 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_19_port, B1 => 
                           n3854, B2 => REGISTERS_10_19_port, ZN => n3378);
   U1592 : NAND4_X1 port map( A1 => n3381, A2 => n3380, A3 => n3379, A4 => 
                           n3378, ZN => n3382);
   U1593 : AOI22_X1 port map( A1 => n3705, A2 => n3383, B1 => n3703, B2 => 
                           n3382, ZN => n3384);
   U1594 : OAI21_X1 port map( B1 => n3866, B2 => n3385, A => n3384, ZN => N436)
                           ;
   U1595 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_18_port, B1 => 
                           n3787, B2 => REGISTERS_31_18_port, ZN => n3389);
   U1596 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_18_port, B1 => 
                           n3658, B2 => REGISTERS_30_18_port, ZN => n3388);
   U1597 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_18_port, B1 => 
                           n3828, B2 => REGISTERS_21_18_port, ZN => n3387);
   U1598 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_18_port, B1 => 
                           n3734, B2 => REGISTERS_22_18_port, ZN => n3386);
   U1599 : NAND4_X1 port map( A1 => n3389, A2 => n3388, A3 => n3387, A4 => 
                           n3386, ZN => n3396);
   U1600 : AOI22_X1 port map( A1 => n3569, A2 => REGISTERS_19_18_port, B1 => 
                           n3817, B2 => REGISTERS_23_18_port, ZN => n3394);
   U1601 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_18_port, B1 => 
                           n3755, B2 => REGISTERS_17_18_port, ZN => n3393);
   U1602 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_18_port, B1 => 
                           n3829, B2 => REGISTERS_18_18_port, ZN => n3392);
   U1603 : AOI22_X1 port map( A1 => n3390, A2 => REGISTERS_25_18_port, B1 => 
                           n3616, B2 => REGISTERS_27_18_port, ZN => n3391);
   U1604 : NAND4_X1 port map( A1 => n3394, A2 => n3393, A3 => n3392, A4 => 
                           n3391, ZN => n3395);
   U1605 : NOR2_X1 port map( A1 => n3396, A2 => n3395, ZN => n3408);
   U1606 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_18_port, B1 => 
                           n3848, B2 => REGISTERS_5_18_port, ZN => n3400);
   U1607 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_1_18_port, B1 => 
                           n3627, B2 => REGISTERS_7_18_port, ZN => n3399);
   U1608 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_6_18_port, B1 => 
                           n3805, B2 => REGISTERS_3_18_port, ZN => n3398);
   U1609 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_18_port, B1 => 
                           n3746, B2 => REGISTERS_2_18_port, ZN => n3397);
   U1610 : NAND4_X1 port map( A1 => n3400, A2 => n3399, A3 => n3398, A4 => 
                           n3397, ZN => n3406);
   U1611 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_9_18_port, B1 => 
                           n3852, B2 => REGISTERS_15_18_port, ZN => n3404);
   U1612 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_18_port, B1 => 
                           n3777, B2 => REGISTERS_12_18_port, ZN => n3403);
   U1613 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_14_18_port, B1 => 
                           n3854, B2 => REGISTERS_10_18_port, ZN => n3402);
   U1614 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_18_port, B1 => 
                           n3805, B2 => REGISTERS_11_18_port, ZN => n3401);
   U1615 : NAND4_X1 port map( A1 => n3404, A2 => n3403, A3 => n3402, A4 => 
                           n3401, ZN => n3405);
   U1616 : AOI22_X1 port map( A1 => n3705, A2 => n3406, B1 => n3703, B2 => 
                           n3405, ZN => n3407);
   U1617 : OAI21_X1 port map( B1 => n3866, B2 => n3408, A => n3407, ZN => N435)
                           ;
   U1618 : AOI22_X1 port map( A1 => n3569, A2 => REGISTERS_19_17_port, B1 => 
                           n3819, B2 => REGISTERS_25_17_port, ZN => n3412);
   U1619 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_17_port, B1 => 
                           n3588, B2 => REGISTERS_20_17_port, ZN => n3411);
   U1620 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_17_port, B1 => 
                           n3658, B2 => REGISTERS_30_17_port, ZN => n3410);
   U1621 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_17_port, B1 => 
                           n3616, B2 => REGISTERS_27_17_port, ZN => n3409);
   U1622 : NAND4_X1 port map( A1 => n3412, A2 => n3411, A3 => n3410, A4 => 
                           n3409, ZN => n3418);
   U1623 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_17_port, B1 => 
                           n3829, B2 => REGISTERS_18_17_port, ZN => n3416);
   U1624 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_17_port, B1 => 
                           n3830, B2 => REGISTERS_26_17_port, ZN => n3415);
   U1625 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_17_port, B1 => 
                           n3659, B2 => REGISTERS_28_17_port, ZN => n3414);
   U1626 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_17_port, B1 => 
                           n3817, B2 => REGISTERS_23_17_port, ZN => n3413);
   U1627 : NAND4_X1 port map( A1 => n3416, A2 => n3415, A3 => n3414, A4 => 
                           n3413, ZN => n3417);
   U1628 : NOR2_X1 port map( A1 => n3418, A2 => n3417, ZN => n3430);
   U1629 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_4_17_port, B1 => 
                           n3852, B2 => REGISTERS_7_17_port, ZN => n3422);
   U1630 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_17_port, B1 => 
                           n3799, B2 => REGISTERS_6_17_port, ZN => n3421);
   U1631 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_17_port, B1 => 
                           n3746, B2 => REGISTERS_2_17_port, ZN => n3420);
   U1632 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_17_port, B1 => 
                           n3805, B2 => REGISTERS_3_17_port, ZN => n3419);
   U1633 : NAND4_X1 port map( A1 => n3422, A2 => n3421, A3 => n3420, A4 => 
                           n3419, ZN => n3428);
   U1634 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_17_port, B1 => 
                           n3841, B2 => REGISTERS_12_17_port, ZN => n3426);
   U1635 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_17_port, B1 => 
                           n3805, B2 => REGISTERS_11_17_port, ZN => n3425);
   U1636 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_17_port, B1 => 
                           n3854, B2 => REGISTERS_10_17_port, ZN => n3424);
   U1637 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_9_17_port, B1 => 
                           n3852, B2 => REGISTERS_15_17_port, ZN => n3423);
   U1638 : NAND4_X1 port map( A1 => n3426, A2 => n3425, A3 => n3424, A4 => 
                           n3423, ZN => n3427);
   U1639 : AOI22_X1 port map( A1 => n3705, A2 => n3428, B1 => n3703, B2 => 
                           n3427, ZN => n3429);
   U1640 : OAI21_X1 port map( B1 => n3866, B2 => n3430, A => n3429, ZN => N434)
                           ;
   U1641 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_16_port, B1 => 
                           n3818, B2 => REGISTERS_20_16_port, ZN => n3434);
   U1642 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_16_port, B1 => 
                           n3829, B2 => REGISTERS_18_16_port, ZN => n3433);
   U1643 : AOI22_X1 port map( A1 => n3761, A2 => REGISTERS_21_16_port, B1 => 
                           n3819, B2 => REGISTERS_25_16_port, ZN => n3432);
   U1644 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_16_port, B1 => 
                           n3616, B2 => REGISTERS_27_16_port, ZN => n3431);
   U1645 : NAND4_X1 port map( A1 => n3434, A2 => n3433, A3 => n3432, A4 => 
                           n3431, ZN => n3440);
   U1646 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_16_port, B1 => 
                           n3817, B2 => REGISTERS_23_16_port, ZN => n3438);
   U1647 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_16_port, B1 => 
                           n3830, B2 => REGISTERS_26_16_port, ZN => n3437);
   U1648 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_16_port, B1 => 
                           n3787, B2 => REGISTERS_31_16_port, ZN => n3436);
   U1649 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_16_port, B1 => 
                           n3734, B2 => REGISTERS_22_16_port, ZN => n3435);
   U1650 : NAND4_X1 port map( A1 => n3438, A2 => n3437, A3 => n3436, A4 => 
                           n3435, ZN => n3439);
   U1651 : NOR2_X1 port map( A1 => n3440, A2 => n3439, ZN => n3452);
   U1652 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_16_port, B1 => 
                           n3805, B2 => REGISTERS_3_16_port, ZN => n3444);
   U1653 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_16_port, B1 => 
                           n3852, B2 => REGISTERS_7_16_port, ZN => n3443);
   U1654 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_4_16_port, B1 => 
                           n3854, B2 => REGISTERS_2_16_port, ZN => n3442);
   U1655 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_5_16_port, B1 => 
                           n3776, B2 => REGISTERS_6_16_port, ZN => n3441);
   U1656 : NAND4_X1 port map( A1 => n3444, A2 => n3443, A3 => n3442, A4 => 
                           n3441, ZN => n3450);
   U1657 : AOI22_X1 port map( A1 => n3843, A2 => REGISTERS_11_16_port, B1 => 
                           n3842, B2 => REGISTERS_10_16_port, ZN => n3448);
   U1658 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_16_port, B1 => 
                           n3776, B2 => REGISTERS_14_16_port, ZN => n3447);
   U1659 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_16_port, B1 => 
                           n3741, B2 => REGISTERS_9_16_port, ZN => n3446);
   U1660 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_16_port, B1 => 
                           n3852, B2 => REGISTERS_15_16_port, ZN => n3445);
   U1661 : NAND4_X1 port map( A1 => n3448, A2 => n3447, A3 => n3446, A4 => 
                           n3445, ZN => n3449);
   U1662 : AOI22_X1 port map( A1 => n3705, A2 => n3450, B1 => n3703, B2 => 
                           n3449, ZN => n3451);
   U1663 : OAI21_X1 port map( B1 => n3866, B2 => n3452, A => n3451, ZN => N433)
                           ;
   U1664 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_15_port, B1 => 
                           n3761, B2 => REGISTERS_21_15_port, ZN => n3456);
   U1665 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_15_port, B1 => 
                           n3817, B2 => REGISTERS_23_15_port, ZN => n3455);
   U1666 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_15_port, B1 => 
                           n3658, B2 => REGISTERS_30_15_port, ZN => n3454);
   U1667 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_15_port, B1 => 
                           n3819, B2 => REGISTERS_25_15_port, ZN => n3453);
   U1668 : NAND4_X1 port map( A1 => n3456, A2 => n3455, A3 => n3454, A4 => 
                           n3453, ZN => n3462);
   U1669 : AOI22_X1 port map( A1 => n3588, A2 => REGISTERS_20_15_port, B1 => 
                           n3616, B2 => REGISTERS_27_15_port, ZN => n3460);
   U1670 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_15_port, B1 => 
                           n3830, B2 => REGISTERS_26_15_port, ZN => n3459);
   U1671 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_15_port, B1 => 
                           n3829, B2 => REGISTERS_18_15_port, ZN => n3458);
   U1672 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_15_port, B1 => 
                           n3832, B2 => REGISTERS_19_15_port, ZN => n3457);
   U1673 : NAND4_X1 port map( A1 => n3460, A2 => n3459, A3 => n3458, A4 => 
                           n3457, ZN => n3461);
   U1674 : NOR2_X1 port map( A1 => n3462, A2 => n3461, ZN => n3474);
   U1675 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_15_port, B1 => 
                           n3741, B2 => REGISTERS_1_15_port, ZN => n3466);
   U1676 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_15_port, B1 => 
                           n3848, B2 => REGISTERS_5_15_port, ZN => n3465);
   U1677 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_6_15_port, B1 => 
                           n3854, B2 => REGISTERS_2_15_port, ZN => n3464);
   U1678 : AOI22_X1 port map( A1 => n3853, A2 => REGISTERS_3_15_port, B1 => 
                           n3852, B2 => REGISTERS_7_15_port, ZN => n3463);
   U1679 : NAND4_X1 port map( A1 => n3466, A2 => n3465, A3 => n3464, A4 => 
                           n3463, ZN => n3472);
   U1680 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_15_port, B1 => 
                           n3852, B2 => REGISTERS_15_15_port, ZN => n3470);
   U1681 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_15_port, B1 => 
                           n3741, B2 => REGISTERS_9_15_port, ZN => n3469);
   U1682 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_15_port, B1 => 
                           n3746, B2 => REGISTERS_10_15_port, ZN => n3468);
   U1683 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_14_15_port, B1 => 
                           n3805, B2 => REGISTERS_11_15_port, ZN => n3467);
   U1684 : NAND4_X1 port map( A1 => n3470, A2 => n3469, A3 => n3468, A4 => 
                           n3467, ZN => n3471);
   U1685 : AOI22_X1 port map( A1 => n3705, A2 => n3472, B1 => n3703, B2 => 
                           n3471, ZN => n3473);
   U1686 : OAI21_X1 port map( B1 => n3814, B2 => n3474, A => n3473, ZN => N432)
                           ;
   U1687 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_14_port, B1 => 
                           n3761, B2 => REGISTERS_21_14_port, ZN => n3478);
   U1688 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_14_port, B1 => 
                           n3830, B2 => REGISTERS_26_14_port, ZN => n3477);
   U1689 : AOI22_X1 port map( A1 => n3568, A2 => REGISTERS_18_14_port, B1 => 
                           n3616, B2 => REGISTERS_27_14_port, ZN => n3476);
   U1690 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_14_port, B1 => 
                           n3817, B2 => REGISTERS_23_14_port, ZN => n3475);
   U1691 : NAND4_X1 port map( A1 => n3478, A2 => n3477, A3 => n3476, A4 => 
                           n3475, ZN => n3484);
   U1692 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_14_port, B1 => 
                           n3832, B2 => REGISTERS_19_14_port, ZN => n3482);
   U1693 : AOI22_X1 port map( A1 => n3659, A2 => REGISTERS_28_14_port, B1 => 
                           n3819, B2 => REGISTERS_25_14_port, ZN => n3481);
   U1694 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_14_port, B1 => 
                           n3787, B2 => REGISTERS_31_14_port, ZN => n3480);
   U1695 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_14_port, B1 => 
                           n3818, B2 => REGISTERS_20_14_port, ZN => n3479);
   U1696 : NAND4_X1 port map( A1 => n3482, A2 => n3481, A3 => n3480, A4 => 
                           n3479, ZN => n3483);
   U1697 : NOR2_X1 port map( A1 => n3484, A2 => n3483, ZN => n3496);
   U1698 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_14_port, B1 => 
                           n3854, B2 => REGISTERS_2_14_port, ZN => n3488);
   U1699 : AOI22_X1 port map( A1 => n3843, A2 => REGISTERS_3_14_port, B1 => 
                           n3852, B2 => REGISTERS_7_14_port, ZN => n3487);
   U1700 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_14_port, B1 => 
                           n3848, B2 => REGISTERS_5_14_port, ZN => n3486);
   U1701 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_4_14_port, B1 => 
                           n3776, B2 => REGISTERS_6_14_port, ZN => n3485);
   U1702 : NAND4_X1 port map( A1 => n3488, A2 => n3487, A3 => n3486, A4 => 
                           n3485, ZN => n3494);
   U1703 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_8_14_port, B1 => 
                           n3842, B2 => REGISTERS_10_14_port, ZN => n3492);
   U1704 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_14_14_port, B1 => 
                           n3850, B2 => REGISTERS_9_14_port, ZN => n3491);
   U1705 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_14_port, B1 => 
                           n3777, B2 => REGISTERS_12_14_port, ZN => n3490);
   U1706 : AOI22_X1 port map( A1 => n3805, A2 => REGISTERS_11_14_port, B1 => 
                           n3852, B2 => REGISTERS_15_14_port, ZN => n3489);
   U1707 : NAND4_X1 port map( A1 => n3492, A2 => n3491, A3 => n3490, A4 => 
                           n3489, ZN => n3493);
   U1708 : AOI22_X1 port map( A1 => n3705, A2 => n3494, B1 => n3703, B2 => 
                           n3493, ZN => n3495);
   U1709 : OAI21_X1 port map( B1 => n3866, B2 => n3496, A => n3495, ZN => N431)
                           ;
   U1710 : AOI22_X1 port map( A1 => n3815, A2 => REGISTERS_16_13_port, B1 => 
                           n3755, B2 => REGISTERS_17_13_port, ZN => n3500);
   U1711 : AOI22_X1 port map( A1 => n3659, A2 => REGISTERS_28_13_port, B1 => 
                           n3832, B2 => REGISTERS_19_13_port, ZN => n3499);
   U1712 : AOI22_X1 port map( A1 => n3664, A2 => REGISTERS_29_13_port, B1 => 
                           n3818, B2 => REGISTERS_20_13_port, ZN => n3498);
   U1713 : AOI22_X1 port map( A1 => n3756, A2 => REGISTERS_23_13_port, B1 => 
                           n3616, B2 => REGISTERS_27_13_port, ZN => n3497);
   U1714 : NAND4_X1 port map( A1 => n3500, A2 => n3499, A3 => n3498, A4 => 
                           n3497, ZN => n3506);
   U1715 : AOI22_X1 port map( A1 => n3734, A2 => REGISTERS_22_13_port, B1 => 
                           n3787, B2 => REGISTERS_31_13_port, ZN => n3504);
   U1716 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_13_port, B1 => 
                           n3819, B2 => REGISTERS_25_13_port, ZN => n3503);
   U1717 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_13_port, B1 => 
                           n3830, B2 => REGISTERS_26_13_port, ZN => n3502);
   U1718 : AOI22_X1 port map( A1 => n3761, A2 => REGISTERS_21_13_port, B1 => 
                           n3829, B2 => REGISTERS_18_13_port, ZN => n3501);
   U1719 : NAND4_X1 port map( A1 => n3504, A2 => n3503, A3 => n3502, A4 => 
                           n3501, ZN => n3505);
   U1720 : NOR2_X1 port map( A1 => n3506, A2 => n3505, ZN => n3518);
   U1721 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_0_13_port, B1 => 
                           n3805, B2 => REGISTERS_3_13_port, ZN => n3510);
   U1722 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_13_port, B1 => 
                           n3776, B2 => REGISTERS_6_13_port, ZN => n3509);
   U1723 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_13_port, B1 => 
                           n3627, B2 => REGISTERS_7_13_port, ZN => n3508);
   U1724 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_13_port, B1 => 
                           n3746, B2 => REGISTERS_2_13_port, ZN => n3507);
   U1725 : NAND4_X1 port map( A1 => n3510, A2 => n3509, A3 => n3508, A4 => 
                           n3507, ZN => n3516);
   U1726 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_13_port, B1 => 
                           n3627, B2 => REGISTERS_15_13_port, ZN => n3514);
   U1727 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_13_port, B1 => 
                           n3842, B2 => REGISTERS_10_13_port, ZN => n3513);
   U1728 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_13_port, B1 => 
                           n3776, B2 => REGISTERS_14_13_port, ZN => n3512);
   U1729 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_9_13_port, B1 => 
                           n3805, B2 => REGISTERS_11_13_port, ZN => n3511);
   U1730 : NAND4_X1 port map( A1 => n3514, A2 => n3513, A3 => n3512, A4 => 
                           n3511, ZN => n3515);
   U1731 : AOI22_X1 port map( A1 => n3705, A2 => n3516, B1 => n3703, B2 => 
                           n3515, ZN => n3517);
   U1732 : OAI21_X1 port map( B1 => n3814, B2 => n3518, A => n3517, ZN => N430)
                           ;
   U1733 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_12_port, B1 => 
                           n3817, B2 => REGISTERS_23_12_port, ZN => n3522);
   U1734 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_12_port, B1 => 
                           n3734, B2 => REGISTERS_22_12_port, ZN => n3521);
   U1735 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_12_port, B1 => 
                           n3818, B2 => REGISTERS_20_12_port, ZN => n3520);
   U1736 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_12_port, B1 => 
                           n3829, B2 => REGISTERS_18_12_port, ZN => n3519);
   U1737 : NAND4_X1 port map( A1 => n3522, A2 => n3521, A3 => n3520, A4 => 
                           n3519, ZN => n3528);
   U1738 : AOI22_X1 port map( A1 => n3664, A2 => REGISTERS_29_12_port, B1 => 
                           n3761, B2 => REGISTERS_21_12_port, ZN => n3526);
   U1739 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_12_port, B1 => 
                           n3819, B2 => REGISTERS_25_12_port, ZN => n3525);
   U1740 : AOI22_X1 port map( A1 => n3815, A2 => REGISTERS_16_12_port, B1 => 
                           n3832, B2 => REGISTERS_19_12_port, ZN => n3524);
   U1741 : AOI22_X1 port map( A1 => n3659, A2 => REGISTERS_28_12_port, B1 => 
                           n3616, B2 => REGISTERS_27_12_port, ZN => n3523);
   U1742 : NAND4_X1 port map( A1 => n3526, A2 => n3525, A3 => n3524, A4 => 
                           n3523, ZN => n3527);
   U1743 : NOR2_X1 port map( A1 => n3528, A2 => n3527, ZN => n3540);
   U1744 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_12_port, B1 => 
                           n3850, B2 => REGISTERS_1_12_port, ZN => n3532);
   U1745 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_12_port, B1 => 
                           n3627, B2 => REGISTERS_7_12_port, ZN => n3531);
   U1746 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_12_port, B1 => 
                           n3854, B2 => REGISTERS_2_12_port, ZN => n3530);
   U1747 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_12_port, B1 => 
                           n3843, B2 => REGISTERS_3_12_port, ZN => n3529);
   U1748 : NAND4_X1 port map( A1 => n3532, A2 => n3531, A3 => n3530, A4 => 
                           n3529, ZN => n3538);
   U1749 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_14_12_port, B1 => 
                           n3843, B2 => REGISTERS_11_12_port, ZN => n3536);
   U1750 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_8_12_port, B1 => 
                           n3627, B2 => REGISTERS_15_12_port, ZN => n3535);
   U1751 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_12_port, B1 => 
                           n3850, B2 => REGISTERS_9_12_port, ZN => n3534);
   U1752 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_12_12_port, B1 => 
                           n3842, B2 => REGISTERS_10_12_port, ZN => n3533);
   U1753 : NAND4_X1 port map( A1 => n3536, A2 => n3535, A3 => n3534, A4 => 
                           n3533, ZN => n3537);
   U1754 : AOI22_X1 port map( A1 => n3705, A2 => n3538, B1 => n3703, B2 => 
                           n3537, ZN => n3539);
   U1755 : OAI21_X1 port map( B1 => n3866, B2 => n3540, A => n3539, ZN => N429)
                           ;
   U1756 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_11_port, B1 => 
                           n3817, B2 => REGISTERS_23_11_port, ZN => n3544);
   U1757 : AOI22_X1 port map( A1 => n3664, A2 => REGISTERS_29_11_port, B1 => 
                           n3818, B2 => REGISTERS_20_11_port, ZN => n3543);
   U1758 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_11_port, B1 => 
                           n3616, B2 => REGISTERS_27_11_port, ZN => n3542);
   U1759 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_11_port, B1 => 
                           n3832, B2 => REGISTERS_19_11_port, ZN => n3541);
   U1760 : NAND4_X1 port map( A1 => n3544, A2 => n3543, A3 => n3542, A4 => 
                           n3541, ZN => n3550);
   U1761 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_11_port, B1 => 
                           n3819, B2 => REGISTERS_25_11_port, ZN => n3548);
   U1762 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_11_port, B1 => 
                           n3658, B2 => REGISTERS_30_11_port, ZN => n3547);
   U1763 : AOI22_X1 port map( A1 => n3734, A2 => REGISTERS_22_11_port, B1 => 
                           n3787, B2 => REGISTERS_31_11_port, ZN => n3546);
   U1764 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_11_port, B1 => 
                           n3829, B2 => REGISTERS_18_11_port, ZN => n3545);
   U1765 : NAND4_X1 port map( A1 => n3548, A2 => n3547, A3 => n3546, A4 => 
                           n3545, ZN => n3549);
   U1766 : NOR2_X1 port map( A1 => n3550, A2 => n3549, ZN => n3563);
   U1767 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_6_11_port, B1 => 
                           n3843, B2 => REGISTERS_3_11_port, ZN => n3554);
   U1768 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_11_port, B1 => 
                           n3850, B2 => REGISTERS_1_11_port, ZN => n3553);
   U1769 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_11_port, B1 => 
                           n3627, B2 => REGISTERS_7_11_port, ZN => n3552);
   U1770 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_11_port, B1 => 
                           n3777, B2 => REGISTERS_4_11_port, ZN => n3551);
   U1771 : NAND4_X1 port map( A1 => n3554, A2 => n3553, A3 => n3552, A4 => 
                           n3551, ZN => n3561);
   U1772 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_11_port, B1 => 
                           n3627, B2 => REGISTERS_15_11_port, ZN => n3559);
   U1773 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_11_port, B1 => 
                           n3776, B2 => REGISTERS_14_11_port, ZN => n3558);
   U1774 : AOI22_X1 port map( A1 => n3805, A2 => REGISTERS_11_11_port, B1 => 
                           n3746, B2 => REGISTERS_10_11_port, ZN => n3557);
   U1775 : AOI22_X1 port map( A1 => n3555, A2 => REGISTERS_8_11_port, B1 => 
                           n3850, B2 => REGISTERS_9_11_port, ZN => n3556);
   U1776 : NAND4_X1 port map( A1 => n3559, A2 => n3558, A3 => n3557, A4 => 
                           n3556, ZN => n3560);
   U1777 : AOI22_X1 port map( A1 => n3705, A2 => n3561, B1 => n3703, B2 => 
                           n3560, ZN => n3562);
   U1778 : OAI21_X1 port map( B1 => n3866, B2 => n3563, A => n3562, ZN => N428)
                           ;
   U1779 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_10_port, B1 => 
                           n3761, B2 => REGISTERS_21_10_port, ZN => n3567);
   U1780 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_10_port, B1 => 
                           n3819, B2 => REGISTERS_25_10_port, ZN => n3566);
   U1781 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_10_port, B1 => 
                           n3815, B2 => REGISTERS_16_10_port, ZN => n3565);
   U1782 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_10_port, B1 => 
                           n3817, B2 => REGISTERS_23_10_port, ZN => n3564);
   U1783 : NAND4_X1 port map( A1 => n3567, A2 => n3566, A3 => n3565, A4 => 
                           n3564, ZN => n3575);
   U1784 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_10_port, B1 => 
                           n3616, B2 => REGISTERS_27_10_port, ZN => n3573);
   U1785 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_10_port, B1 => 
                           n3755, B2 => REGISTERS_17_10_port, ZN => n3572);
   U1786 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_10_port, B1 => 
                           n3830, B2 => REGISTERS_26_10_port, ZN => n3571);
   U1787 : AOI22_X1 port map( A1 => n3569, A2 => REGISTERS_19_10_port, B1 => 
                           n3568, B2 => REGISTERS_18_10_port, ZN => n3570);
   U1788 : NAND4_X1 port map( A1 => n3573, A2 => n3572, A3 => n3571, A4 => 
                           n3570, ZN => n3574);
   U1789 : NOR2_X1 port map( A1 => n3575, A2 => n3574, ZN => n3587);
   U1790 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_10_port, B1 => 
                           n3746, B2 => REGISTERS_2_10_port, ZN => n3579);
   U1791 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_10_port, B1 => 
                           n3850, B2 => REGISTERS_1_10_port, ZN => n3578);
   U1792 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_0_10_port, B1 => 
                           n3799, B2 => REGISTERS_6_10_port, ZN => n3577);
   U1793 : AOI22_X1 port map( A1 => n3843, A2 => REGISTERS_3_10_port, B1 => 
                           n3627, B2 => REGISTERS_7_10_port, ZN => n3576);
   U1794 : NAND4_X1 port map( A1 => n3579, A2 => n3578, A3 => n3577, A4 => 
                           n3576, ZN => n3585);
   U1795 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_14_10_port, B1 => 
                           n3854, B2 => REGISTERS_10_10_port, ZN => n3583);
   U1796 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_10_port, B1 => 
                           n3777, B2 => REGISTERS_12_10_port, ZN => n3582);
   U1797 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_9_10_port, B1 => 
                           n3843, B2 => REGISTERS_11_10_port, ZN => n3581);
   U1798 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_8_10_port, B1 => 
                           n3627, B2 => REGISTERS_15_10_port, ZN => n3580);
   U1799 : NAND4_X1 port map( A1 => n3583, A2 => n3582, A3 => n3581, A4 => 
                           n3580, ZN => n3584);
   U1800 : AOI22_X1 port map( A1 => n3705, A2 => n3585, B1 => n3703, B2 => 
                           n3584, ZN => n3586);
   U1801 : OAI21_X1 port map( B1 => n3866, B2 => n3587, A => n3586, ZN => N427)
                           ;
   U1802 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_9_port, B1 => 
                           n3659, B2 => REGISTERS_28_9_port, ZN => n3592);
   U1803 : AOI22_X1 port map( A1 => n3588, A2 => REGISTERS_20_9_port, B1 => 
                           n3616, B2 => REGISTERS_27_9_port, ZN => n3591);
   U1804 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_9_port, B1 => 
                           n3819, B2 => REGISTERS_25_9_port, ZN => n3590);
   U1805 : AOI22_X1 port map( A1 => n3821, A2 => REGISTERS_17_9_port, B1 => 
                           n3817, B2 => REGISTERS_23_9_port, ZN => n3589);
   U1806 : NAND4_X1 port map( A1 => n3592, A2 => n3591, A3 => n3590, A4 => 
                           n3589, ZN => n3598);
   U1807 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_9_port, B1 => 
                           n3832, B2 => REGISTERS_19_9_port, ZN => n3596);
   U1808 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_9_port, B1 => 
                           n3787, B2 => REGISTERS_31_9_port, ZN => n3595);
   U1809 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_9_port, B1 => 
                           n3658, B2 => REGISTERS_30_9_port, ZN => n3594);
   U1810 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_9_port, B1 => 
                           n3829, B2 => REGISTERS_18_9_port, ZN => n3593);
   U1811 : NAND4_X1 port map( A1 => n3596, A2 => n3595, A3 => n3594, A4 => 
                           n3593, ZN => n3597);
   U1812 : NOR2_X1 port map( A1 => n3598, A2 => n3597, ZN => n3610);
   U1813 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_1_9_port, B1 => 
                           n3842, B2 => REGISTERS_2_9_port, ZN => n3602);
   U1814 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_9_port, B1 => 
                           n3799, B2 => REGISTERS_6_9_port, ZN => n3601);
   U1815 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_4_9_port, B1 => 
                           n3843, B2 => REGISTERS_3_9_port, ZN => n3600);
   U1816 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_0_9_port, B1 => 
                           n3627, B2 => REGISTERS_7_9_port, ZN => n3599);
   U1817 : NAND4_X1 port map( A1 => n3602, A2 => n3601, A3 => n3600, A4 => 
                           n3599, ZN => n3608);
   U1818 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_9_9_port, B1 => 
                           n3746, B2 => REGISTERS_10_9_port, ZN => n3606);
   U1819 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_9_port, B1 => 
                           n3627, B2 => REGISTERS_15_9_port, ZN => n3605);
   U1820 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_9_port, B1 => 
                           n3843, B2 => REGISTERS_11_9_port, ZN => n3604);
   U1821 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_8_9_port, B1 => 
                           n3777, B2 => REGISTERS_12_9_port, ZN => n3603);
   U1822 : NAND4_X1 port map( A1 => n3606, A2 => n3605, A3 => n3604, A4 => 
                           n3603, ZN => n3607);
   U1823 : AOI22_X1 port map( A1 => n3705, A2 => n3608, B1 => n3703, B2 => 
                           n3607, ZN => n3609);
   U1824 : OAI21_X1 port map( B1 => n3814, B2 => n3610, A => n3609, ZN => N426)
                           ;
   U1825 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_8_port, B1 => 
                           n3786, B2 => REGISTERS_26_8_port, ZN => n3615);
   U1826 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_8_port, B1 => 
                           n3658, B2 => REGISTERS_30_8_port, ZN => n3614);
   U1827 : AOI22_X1 port map( A1 => n3611, A2 => REGISTERS_24_8_port, B1 => 
                           n3832, B2 => REGISTERS_19_8_port, ZN => n3613);
   U1828 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_8_port, B1 => 
                           n3829, B2 => REGISTERS_18_8_port, ZN => n3612);
   U1829 : NAND4_X1 port map( A1 => n3615, A2 => n3614, A3 => n3613, A4 => 
                           n3612, ZN => n3622);
   U1830 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_8_port, B1 => 
                           n3616, B2 => REGISTERS_27_8_port, ZN => n3620);
   U1831 : AOI22_X1 port map( A1 => n3819, A2 => REGISTERS_25_8_port, B1 => 
                           n3817, B2 => REGISTERS_23_8_port, ZN => n3619);
   U1832 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_8_port, B1 => 
                           n3755, B2 => REGISTERS_17_8_port, ZN => n3618);
   U1833 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_8_port, B1 => 
                           n3818, B2 => REGISTERS_20_8_port, ZN => n3617);
   U1834 : NAND4_X1 port map( A1 => n3620, A2 => n3619, A3 => n3618, A4 => 
                           n3617, ZN => n3621);
   U1835 : NOR2_X1 port map( A1 => n3622, A2 => n3621, ZN => n3635);
   U1836 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_8_port, B1 => 
                           n3627, B2 => REGISTERS_7_8_port, ZN => n3626);
   U1837 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_6_8_port, B1 => 
                           n3854, B2 => REGISTERS_2_8_port, ZN => n3625);
   U1838 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_0_8_port, B1 => 
                           n3850, B2 => REGISTERS_1_8_port, ZN => n3624);
   U1839 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_8_port, B1 => 
                           n3843, B2 => REGISTERS_3_8_port, ZN => n3623);
   U1840 : NAND4_X1 port map( A1 => n3626, A2 => n3625, A3 => n3624, A4 => 
                           n3623, ZN => n3633);
   U1841 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_8_port, B1 => 
                           n3627, B2 => REGISTERS_15_8_port, ZN => n3631);
   U1842 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_14_8_port, B1 => 
                           n3842, B2 => REGISTERS_10_8_port, ZN => n3630);
   U1843 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_9_8_port, B1 => 
                           n3805, B2 => REGISTERS_11_8_port, ZN => n3629);
   U1844 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_8_8_port, B1 => 
                           n3851, B2 => REGISTERS_12_8_port, ZN => n3628);
   U1845 : NAND4_X1 port map( A1 => n3631, A2 => n3630, A3 => n3629, A4 => 
                           n3628, ZN => n3632);
   U1846 : AOI22_X1 port map( A1 => n3705, A2 => n3633, B1 => n3703, B2 => 
                           n3632, ZN => n3634);
   U1847 : OAI21_X1 port map( B1 => n3866, B2 => n3635, A => n3634, ZN => N425)
                           ;
   U1848 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_7_port, B1 => 
                           n3819, B2 => REGISTERS_25_7_port, ZN => n3639);
   U1849 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_7_port, B1 => 
                           n3829, B2 => REGISTERS_18_7_port, ZN => n3638);
   U1850 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_7_port, B1 => 
                           n3833, B2 => REGISTERS_31_7_port, ZN => n3637);
   U1851 : AOI22_X1 port map( A1 => n3821, A2 => REGISTERS_17_7_port, B1 => 
                           n3831, B2 => REGISTERS_30_7_port, ZN => n3636);
   U1852 : NAND4_X1 port map( A1 => n3639, A2 => n3638, A3 => n3637, A4 => 
                           n3636, ZN => n3645);
   U1853 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_7_port, B1 => 
                           n3761, B2 => REGISTERS_21_7_port, ZN => n3643);
   U1854 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_7_port, B1 => 
                           n3817, B2 => REGISTERS_23_7_port, ZN => n3642);
   U1855 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_7_port, B1 => 
                           n3832, B2 => REGISTERS_19_7_port, ZN => n3641);
   U1856 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_7_port, B1 => 
                           n3827, B2 => REGISTERS_27_7_port, ZN => n3640);
   U1857 : NAND4_X1 port map( A1 => n3643, A2 => n3642, A3 => n3641, A4 => 
                           n3640, ZN => n3644);
   U1858 : NOR2_X1 port map( A1 => n3645, A2 => n3644, ZN => n3657);
   U1859 : AOI22_X1 port map( A1 => n3805, A2 => REGISTERS_3_7_port, B1 => 
                           n3775, B2 => REGISTERS_7_7_port, ZN => n3649);
   U1860 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_7_port, B1 => 
                           n3799, B2 => REGISTERS_6_7_port, ZN => n3648);
   U1861 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_7_port, B1 => 
                           n3746, B2 => REGISTERS_2_7_port, ZN => n3647);
   U1862 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_7_port, B1 => 
                           n3850, B2 => REGISTERS_1_7_port, ZN => n3646);
   U1863 : NAND4_X1 port map( A1 => n3649, A2 => n3648, A3 => n3647, A4 => 
                           n3646, ZN => n3655);
   U1864 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_7_port, B1 => 
                           n3843, B2 => REGISTERS_11_7_port, ZN => n3653);
   U1865 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_9_7_port, B1 => 
                           n3775, B2 => REGISTERS_15_7_port, ZN => n3652);
   U1866 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_12_7_port, B1 => 
                           n3854, B2 => REGISTERS_10_7_port, ZN => n3651);
   U1867 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_7_port, B1 => 
                           n3799, B2 => REGISTERS_14_7_port, ZN => n3650);
   U1868 : NAND4_X1 port map( A1 => n3653, A2 => n3652, A3 => n3651, A4 => 
                           n3650, ZN => n3654);
   U1869 : AOI22_X1 port map( A1 => n3705, A2 => n3655, B1 => n3703, B2 => 
                           n3654, ZN => n3656);
   U1870 : OAI21_X1 port map( B1 => n3814, B2 => n3657, A => n3656, ZN => N424)
                           ;
   U1871 : AOI22_X1 port map( A1 => n3658, A2 => REGISTERS_30_6_port, B1 => 
                           n3829, B2 => REGISTERS_18_6_port, ZN => n3663);
   U1872 : AOI22_X1 port map( A1 => n3821, A2 => REGISTERS_17_6_port, B1 => 
                           n3818, B2 => REGISTERS_20_6_port, ZN => n3662);
   U1873 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_6_port, B1 => 
                           n3659, B2 => REGISTERS_28_6_port, ZN => n3661);
   U1874 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_6_port, B1 => 
                           n3832, B2 => REGISTERS_19_6_port, ZN => n3660);
   U1875 : NAND4_X1 port map( A1 => n3663, A2 => n3662, A3 => n3661, A4 => 
                           n3660, ZN => n3670);
   U1876 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_6_port, B1 => 
                           n3833, B2 => REGISTERS_31_6_port, ZN => n3668);
   U1877 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_6_port, B1 => 
                           n3819, B2 => REGISTERS_25_6_port, ZN => n3667);
   U1878 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_6_port, B1 => 
                           n3664, B2 => REGISTERS_29_6_port, ZN => n3666);
   U1879 : AOI22_X1 port map( A1 => n3756, A2 => REGISTERS_23_6_port, B1 => 
                           n3827, B2 => REGISTERS_27_6_port, ZN => n3665);
   U1880 : NAND4_X1 port map( A1 => n3668, A2 => n3667, A3 => n3666, A4 => 
                           n3665, ZN => n3669);
   U1881 : NOR2_X1 port map( A1 => n3670, A2 => n3669, ZN => n3683);
   U1882 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_4_6_port, B1 => 
                           n3842, B2 => REGISTERS_2_6_port, ZN => n3674);
   U1883 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_6_port, B1 => 
                           n3848, B2 => REGISTERS_5_6_port, ZN => n3673);
   U1884 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_6_port, B1 => 
                           n3805, B2 => REGISTERS_3_6_port, ZN => n3672);
   U1885 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_1_6_port, B1 => 
                           n3775, B2 => REGISTERS_7_6_port, ZN => n3671);
   U1886 : NAND4_X1 port map( A1 => n3674, A2 => n3673, A3 => n3672, A4 => 
                           n3671, ZN => n3680);
   U1887 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_6_port, B1 => 
                           n3853, B2 => REGISTERS_11_6_port, ZN => n3678);
   U1888 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_9_6_port, B1 => 
                           n3746, B2 => REGISTERS_10_6_port, ZN => n3677);
   U1889 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_6_port, B1 => 
                           n3775, B2 => REGISTERS_15_6_port, ZN => n3676);
   U1890 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_12_6_port, B1 => 
                           n3799, B2 => REGISTERS_14_6_port, ZN => n3675);
   U1891 : NAND4_X1 port map( A1 => n3678, A2 => n3677, A3 => n3676, A4 => 
                           n3675, ZN => n3679);
   U1892 : AOI22_X1 port map( A1 => n3681, A2 => n3680, B1 => n3703, B2 => 
                           n3679, ZN => n3682);
   U1893 : OAI21_X1 port map( B1 => n3866, B2 => n3683, A => n3682, ZN => N423)
                           ;
   U1894 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_5_port, B1 => 
                           n3786, B2 => REGISTERS_26_5_port, ZN => n3687);
   U1895 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_5_port, B1 => 
                           n3817, B2 => REGISTERS_23_5_port, ZN => n3686);
   U1896 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_5_port, B1 => 
                           n3734, B2 => REGISTERS_22_5_port, ZN => n3685);
   U1897 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_5_port, B1 => 
                           n3833, B2 => REGISTERS_31_5_port, ZN => n3684);
   U1898 : NAND4_X1 port map( A1 => n3687, A2 => n3686, A3 => n3685, A4 => 
                           n3684, ZN => n3693);
   U1899 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_5_port, B1 => 
                           n3819, B2 => REGISTERS_25_5_port, ZN => n3691);
   U1900 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_5_port, B1 => 
                           n3827, B2 => REGISTERS_27_5_port, ZN => n3690);
   U1901 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_5_port, B1 => 
                           n3831, B2 => REGISTERS_30_5_port, ZN => n3689);
   U1902 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_5_port, B1 => 
                           n3829, B2 => REGISTERS_18_5_port, ZN => n3688);
   U1903 : NAND4_X1 port map( A1 => n3691, A2 => n3690, A3 => n3689, A4 => 
                           n3688, ZN => n3692);
   U1904 : NOR2_X1 port map( A1 => n3693, A2 => n3692, ZN => n3707);
   U1905 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_1_5_port, B1 => 
                           n3843, B2 => REGISTERS_3_5_port, ZN => n3697);
   U1906 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_5_port, B1 => 
                           n3775, B2 => REGISTERS_7_5_port, ZN => n3696);
   U1907 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_5_port, B1 => 
                           n3799, B2 => REGISTERS_6_5_port, ZN => n3695);
   U1908 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_5_5_port, B1 => 
                           n3777, B2 => REGISTERS_4_5_port, ZN => n3694);
   U1909 : NAND4_X1 port map( A1 => n3697, A2 => n3696, A3 => n3695, A4 => 
                           n3694, ZN => n3704);
   U1910 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_5_port, B1 => 
                           n3777, B2 => REGISTERS_12_5_port, ZN => n3701);
   U1911 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_14_5_port, B1 => 
                           n3775, B2 => REGISTERS_15_5_port, ZN => n3700);
   U1912 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_13_5_port, B1 => 
                           n3854, B2 => REGISTERS_10_5_port, ZN => n3699);
   U1913 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_9_5_port, B1 => 
                           n3805, B2 => REGISTERS_11_5_port, ZN => n3698);
   U1914 : NAND4_X1 port map( A1 => n3701, A2 => n3700, A3 => n3699, A4 => 
                           n3698, ZN => n3702);
   U1915 : AOI22_X1 port map( A1 => n3705, A2 => n3704, B1 => n3703, B2 => 
                           n3702, ZN => n3706);
   U1916 : OAI21_X1 port map( B1 => n3814, B2 => n3707, A => n3706, ZN => N422)
                           ;
   U1917 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_4_port, B1 => 
                           n3832, B2 => REGISTERS_19_4_port, ZN => n3711);
   U1918 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_4_port, B1 => 
                           n3818, B2 => REGISTERS_20_4_port, ZN => n3710);
   U1919 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_4_port, B1 => 
                           n3817, B2 => REGISTERS_23_4_port, ZN => n3709);
   U1920 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_4_port, B1 => 
                           n3829, B2 => REGISTERS_18_4_port, ZN => n3708);
   U1921 : NAND4_X1 port map( A1 => n3711, A2 => n3710, A3 => n3709, A4 => 
                           n3708, ZN => n3717);
   U1922 : AOI22_X1 port map( A1 => n3786, A2 => REGISTERS_26_4_port, B1 => 
                           n3831, B2 => REGISTERS_30_4_port, ZN => n3715);
   U1923 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_4_port, B1 => 
                           n3819, B2 => REGISTERS_25_4_port, ZN => n3714);
   U1924 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_4_port, B1 => 
                           n3827, B2 => REGISTERS_27_4_port, ZN => n3713);
   U1925 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_4_port, B1 => 
                           n3833, B2 => REGISTERS_31_4_port, ZN => n3712);
   U1926 : NAND4_X1 port map( A1 => n3715, A2 => n3714, A3 => n3713, A4 => 
                           n3712, ZN => n3716);
   U1927 : NOR2_X1 port map( A1 => n3717, A2 => n3716, ZN => n3729);
   U1928 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_4_4_port, B1 => 
                           n3850, B2 => REGISTERS_1_4_port, ZN => n3721);
   U1929 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_4_port, B1 => 
                           n3775, B2 => REGISTERS_7_4_port, ZN => n3720);
   U1930 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_4_port, B1 => 
                           n3799, B2 => REGISTERS_6_4_port, ZN => n3719);
   U1931 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_4_port, B1 => 
                           n3853, B2 => REGISTERS_3_4_port, ZN => n3718);
   U1932 : NAND4_X1 port map( A1 => n3721, A2 => n3720, A3 => n3719, A4 => 
                           n3718, ZN => n3727);
   U1933 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_9_4_port, B1 => 
                           n3843, B2 => REGISTERS_11_4_port, ZN => n3725);
   U1934 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_4_port, B1 => 
                           n3775, B2 => REGISTERS_15_4_port, ZN => n3724);
   U1935 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_4_port, B1 => 
                           n3799, B2 => REGISTERS_14_4_port, ZN => n3723);
   U1936 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_4_port, B1 => 
                           n3842, B2 => REGISTERS_10_4_port, ZN => n3722);
   U1937 : NAND4_X1 port map( A1 => n3725, A2 => n3724, A3 => n3723, A4 => 
                           n3722, ZN => n3726);
   U1938 : AOI22_X1 port map( A1 => n3863, A2 => n3727, B1 => n3861, B2 => 
                           n3726, ZN => n3728);
   U1939 : OAI21_X1 port map( B1 => n3866, B2 => n3729, A => n3728, ZN => N421)
                           ;
   U1940 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_3_port, B1 => 
                           n3829, B2 => REGISTERS_18_3_port, ZN => n3733);
   U1941 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_3_port, B1 => 
                           n3819, B2 => REGISTERS_25_3_port, ZN => n3732);
   U1942 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_3_port, B1 => 
                           n3831, B2 => REGISTERS_30_3_port, ZN => n3731);
   U1943 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_3_port, B1 => 
                           n3827, B2 => REGISTERS_27_3_port, ZN => n3730);
   U1944 : NAND4_X1 port map( A1 => n3733, A2 => n3732, A3 => n3731, A4 => 
                           n3730, ZN => n3740);
   U1945 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_3_port, B1 => 
                           n3821, B2 => REGISTERS_17_3_port, ZN => n3738);
   U1946 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_3_port, B1 => 
                           n3786, B2 => REGISTERS_26_3_port, ZN => n3737);
   U1947 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_3_port, B1 => 
                           n3734, B2 => REGISTERS_22_3_port, ZN => n3736);
   U1948 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_3_port, B1 => 
                           n3817, B2 => REGISTERS_23_3_port, ZN => n3735);
   U1949 : NAND4_X1 port map( A1 => n3738, A2 => n3737, A3 => n3736, A4 => 
                           n3735, ZN => n3739);
   U1950 : NOR2_X1 port map( A1 => n3740, A2 => n3739, ZN => n3754);
   U1951 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_3_port, B1 => 
                           n3853, B2 => REGISTERS_3_3_port, ZN => n3745);
   U1952 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_3_port, B1 => 
                           n3854, B2 => REGISTERS_2_3_port, ZN => n3744);
   U1953 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_3_port, B1 => 
                           n3799, B2 => REGISTERS_6_3_port, ZN => n3743);
   U1954 : AOI22_X1 port map( A1 => n3741, A2 => REGISTERS_1_3_port, B1 => 
                           n3775, B2 => REGISTERS_7_3_port, ZN => n3742);
   U1955 : NAND4_X1 port map( A1 => n3745, A2 => n3744, A3 => n3743, A4 => 
                           n3742, ZN => n3752);
   U1956 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_3_port, B1 => 
                           n3798, B2 => REGISTERS_13_3_port, ZN => n3750);
   U1957 : AOI22_X1 port map( A1 => n3777, A2 => REGISTERS_12_3_port, B1 => 
                           n3775, B2 => REGISTERS_15_3_port, ZN => n3749);
   U1958 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_14_3_port, B1 => 
                           n3746, B2 => REGISTERS_10_3_port, ZN => n3748);
   U1959 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_9_3_port, B1 => 
                           n3805, B2 => REGISTERS_11_3_port, ZN => n3747);
   U1960 : NAND4_X1 port map( A1 => n3750, A2 => n3749, A3 => n3748, A4 => 
                           n3747, ZN => n3751);
   U1961 : AOI22_X1 port map( A1 => n3863, A2 => n3752, B1 => n3861, B2 => 
                           n3751, ZN => n3753);
   U1962 : OAI21_X1 port map( B1 => n3814, B2 => n3754, A => n3753, ZN => N420)
                           ;
   U1963 : AOI22_X1 port map( A1 => n3755, A2 => REGISTERS_17_2_port, B1 => 
                           n3831, B2 => REGISTERS_30_2_port, ZN => n3760);
   U1964 : AOI22_X1 port map( A1 => n3756, A2 => REGISTERS_23_2_port, B1 => 
                           n3829, B2 => REGISTERS_18_2_port, ZN => n3759);
   U1965 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_2_port, B1 => 
                           n3818, B2 => REGISTERS_20_2_port, ZN => n3758);
   U1966 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_2_port, B1 => 
                           n3832, B2 => REGISTERS_19_2_port, ZN => n3757);
   U1967 : NAND4_X1 port map( A1 => n3760, A2 => n3759, A3 => n3758, A4 => 
                           n3757, ZN => n3768);
   U1968 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_2_port, B1 => 
                           n3761, B2 => REGISTERS_21_2_port, ZN => n3766);
   U1969 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_2_port, B1 => 
                           n3819, B2 => REGISTERS_25_2_port, ZN => n3765);
   U1970 : AOI22_X1 port map( A1 => n3762, A2 => REGISTERS_16_2_port, B1 => 
                           n3827, B2 => REGISTERS_27_2_port, ZN => n3764);
   U1971 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_2_port, B1 => 
                           n3833, B2 => REGISTERS_31_2_port, ZN => n3763);
   U1972 : NAND4_X1 port map( A1 => n3766, A2 => n3765, A3 => n3764, A4 => 
                           n3763, ZN => n3767);
   U1973 : NOR2_X1 port map( A1 => n3768, A2 => n3767, ZN => n3785);
   U1974 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_2_port, B1 => 
                           n3775, B2 => REGISTERS_7_2_port, ZN => n3773);
   U1975 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_5_2_port, B1 => 
                           n3853, B2 => REGISTERS_3_2_port, ZN => n3772);
   U1976 : AOI22_X1 port map( A1 => n3769, A2 => REGISTERS_0_2_port, B1 => 
                           n3777, B2 => REGISTERS_4_2_port, ZN => n3771);
   U1977 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_6_2_port, B1 => 
                           n3774, B2 => REGISTERS_1_2_port, ZN => n3770);
   U1978 : NAND4_X1 port map( A1 => n3773, A2 => n3772, A3 => n3771, A4 => 
                           n3770, ZN => n3783);
   U1979 : AOI22_X1 port map( A1 => n3774, A2 => REGISTERS_9_2_port, B1 => 
                           n3854, B2 => REGISTERS_10_2_port, ZN => n3781);
   U1980 : AOI22_X1 port map( A1 => n3776, A2 => REGISTERS_14_2_port, B1 => 
                           n3775, B2 => REGISTERS_15_2_port, ZN => n3780);
   U1981 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_2_port, B1 => 
                           n3853, B2 => REGISTERS_11_2_port, ZN => n3779);
   U1982 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_13_2_port, B1 => 
                           n3777, B2 => REGISTERS_12_2_port, ZN => n3778);
   U1983 : NAND4_X1 port map( A1 => n3781, A2 => n3780, A3 => n3779, A4 => 
                           n3778, ZN => n3782);
   U1984 : AOI22_X1 port map( A1 => n3863, A2 => n3783, B1 => n3861, B2 => 
                           n3782, ZN => n3784);
   U1985 : OAI21_X1 port map( B1 => n3866, B2 => n3785, A => n3784, ZN => N419)
                           ;
   U1986 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_1_port, B1 => 
                           n3821, B2 => REGISTERS_17_1_port, ZN => n3791);
   U1987 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_1_port, B1 => 
                           n3786, B2 => REGISTERS_26_1_port, ZN => n3790);
   U1988 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_1_port, B1 => 
                           n3815, B2 => REGISTERS_16_1_port, ZN => n3789);
   U1989 : AOI22_X1 port map( A1 => n3787, A2 => REGISTERS_31_1_port, B1 => 
                           n3817, B2 => REGISTERS_23_1_port, ZN => n3788);
   U1990 : NAND4_X1 port map( A1 => n3791, A2 => n3790, A3 => n3789, A4 => 
                           n3788, ZN => n3797);
   U1991 : AOI22_X1 port map( A1 => n3819, A2 => REGISTERS_25_1_port, B1 => 
                           n3827, B2 => REGISTERS_27_1_port, ZN => n3795);
   U1992 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_1_port, B1 => 
                           n3831, B2 => REGISTERS_30_1_port, ZN => n3794);
   U1993 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_1_port, B1 => 
                           n3818, B2 => REGISTERS_20_1_port, ZN => n3793);
   U1994 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_1_port, B1 => 
                           n3829, B2 => REGISTERS_18_1_port, ZN => n3792);
   U1995 : NAND4_X1 port map( A1 => n3795, A2 => n3794, A3 => n3793, A4 => 
                           n3792, ZN => n3796);
   U1996 : NOR2_X1 port map( A1 => n3797, A2 => n3796, ZN => n3813);
   U1997 : AOI22_X1 port map( A1 => n3798, A2 => REGISTERS_5_1_port, B1 => 
                           n3852, B2 => REGISTERS_7_1_port, ZN => n3803);
   U1998 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_0_1_port, B1 => 
                           n3851, B2 => REGISTERS_4_1_port, ZN => n3802);
   U1999 : AOI22_X1 port map( A1 => n3799, A2 => REGISTERS_6_1_port, B1 => 
                           n3843, B2 => REGISTERS_3_1_port, ZN => n3801);
   U2000 : AOI22_X1 port map( A1 => n3850, A2 => REGISTERS_1_1_port, B1 => 
                           n3842, B2 => REGISTERS_2_1_port, ZN => n3800);
   U2001 : NAND4_X1 port map( A1 => n3803, A2 => n3802, A3 => n3801, A4 => 
                           n3800, ZN => n3811);
   U2002 : AOI22_X1 port map( A1 => n3804, A2 => REGISTERS_13_1_port, B1 => 
                           n3850, B2 => REGISTERS_9_1_port, ZN => n3809);
   U2003 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_10_1_port, B1 => 
                           n3852, B2 => REGISTERS_15_1_port, ZN => n3808);
   U2004 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_1_port, B1 => 
                           n3855, B2 => REGISTERS_14_1_port, ZN => n3807);
   U2005 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_1_port, B1 => 
                           n3805, B2 => REGISTERS_11_1_port, ZN => n3806);
   U2006 : NAND4_X1 port map( A1 => n3809, A2 => n3808, A3 => n3807, A4 => 
                           n3806, ZN => n3810);
   U2007 : AOI22_X1 port map( A1 => n3863, A2 => n3811, B1 => n3861, B2 => 
                           n3810, ZN => n3812);
   U2008 : OAI21_X1 port map( B1 => n3814, B2 => n3813, A => n3812, ZN => N418)
                           ;
   U2009 : AOI22_X1 port map( A1 => n3816, A2 => REGISTERS_24_0_port, B1 => 
                           n3815, B2 => REGISTERS_16_0_port, ZN => n3826);
   U2010 : AOI22_X1 port map( A1 => n3818, A2 => REGISTERS_20_0_port, B1 => 
                           n3817, B2 => REGISTERS_23_0_port, ZN => n3825);
   U2011 : AOI22_X1 port map( A1 => n3820, A2 => REGISTERS_29_0_port, B1 => 
                           n3819, B2 => REGISTERS_25_0_port, ZN => n3824);
   U2012 : AOI22_X1 port map( A1 => n3822, A2 => REGISTERS_22_0_port, B1 => 
                           n3821, B2 => REGISTERS_17_0_port, ZN => n3823);
   U2013 : NAND4_X1 port map( A1 => n3826, A2 => n3825, A3 => n3824, A4 => 
                           n3823, ZN => n3840);
   U2014 : AOI22_X1 port map( A1 => n3828, A2 => REGISTERS_21_0_port, B1 => 
                           n3827, B2 => REGISTERS_27_0_port, ZN => n3838);
   U2015 : AOI22_X1 port map( A1 => n3830, A2 => REGISTERS_26_0_port, B1 => 
                           n3829, B2 => REGISTERS_18_0_port, ZN => n3837);
   U2016 : AOI22_X1 port map( A1 => n3832, A2 => REGISTERS_19_0_port, B1 => 
                           n3831, B2 => REGISTERS_30_0_port, ZN => n3836);
   U2017 : AOI22_X1 port map( A1 => n3834, A2 => REGISTERS_28_0_port, B1 => 
                           n3833, B2 => REGISTERS_31_0_port, ZN => n3835);
   U2018 : NAND4_X1 port map( A1 => n3838, A2 => n3837, A3 => n3836, A4 => 
                           n3835, ZN => n3839);
   U2019 : NOR2_X1 port map( A1 => n3840, A2 => n3839, ZN => n3865);
   U2020 : AOI22_X1 port map( A1 => n3848, A2 => REGISTERS_5_0_port, B1 => 
                           n3855, B2 => REGISTERS_6_0_port, ZN => n3847);
   U2021 : AOI22_X1 port map( A1 => n3841, A2 => REGISTERS_4_0_port, B1 => 
                           n3850, B2 => REGISTERS_1_0_port, ZN => n3846);
   U2022 : AOI22_X1 port map( A1 => n3842, A2 => REGISTERS_2_0_port, B1 => 
                           n3852, B2 => REGISTERS_7_0_port, ZN => n3845);
   U2023 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_0_0_port, B1 => 
                           n3843, B2 => REGISTERS_3_0_port, ZN => n3844);
   U2024 : NAND4_X1 port map( A1 => n3847, A2 => n3846, A3 => n3845, A4 => 
                           n3844, ZN => n3862);
   U2025 : AOI22_X1 port map( A1 => n3849, A2 => REGISTERS_8_0_port, B1 => 
                           n3848, B2 => REGISTERS_13_0_port, ZN => n3859);
   U2026 : AOI22_X1 port map( A1 => n3851, A2 => REGISTERS_12_0_port, B1 => 
                           n3850, B2 => REGISTERS_9_0_port, ZN => n3858);
   U2027 : AOI22_X1 port map( A1 => n3853, A2 => REGISTERS_11_0_port, B1 => 
                           n3852, B2 => REGISTERS_15_0_port, ZN => n3857);
   U2028 : AOI22_X1 port map( A1 => n3855, A2 => REGISTERS_14_0_port, B1 => 
                           n3854, B2 => REGISTERS_10_0_port, ZN => n3856);
   U2029 : NAND4_X1 port map( A1 => n3859, A2 => n3858, A3 => n3857, A4 => 
                           n3856, ZN => n3860);
   U2030 : AOI22_X1 port map( A1 => n3863, A2 => n3862, B1 => n3861, B2 => 
                           n3860, ZN => n3864);
   U2031 : OAI21_X1 port map( B1 => n3866, B2 => n3865, A => n3864, ZN => N417)
                           ;
   U2032 : NAND3_X1 port map( A1 => n2898, A2 => ENABLE, A3 => RD1, ZN => n4647
                           );
   U2033 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n3875);
   U2034 : NOR2_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), ZN => n3867);
   U2035 : INV_X1 port map( A => ADD_RD1(1), ZN => n3873);
   U2036 : NAND2_X1 port map( A1 => n3867, A2 => n3873, ZN => n3883);
   U2037 : NOR2_X1 port map( A1 => n3875, A2 => n3883, ZN => n4396);
   U2038 : CLKBUF_X1 port map( A => n4396, Z => n4612);
   U2039 : INV_X1 port map( A => ADD_RD1(3), ZN => n3892);
   U2040 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n3892, ZN => n3874);
   U2041 : INV_X1 port map( A => ADD_RD1(2), ZN => n3872);
   U2042 : OR3_X1 port map( A1 => n3872, A2 => ADD_RD1(1), A3 => ADD_RD1(0), ZN
                           => n3911);
   U2043 : NOR2_X1 port map( A1 => n3874, A2 => n3911, ZN => n4415);
   U2044 : CLKBUF_X1 port map( A => n4415, Z => n4596);
   U2045 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n4612, B1 => 
                           REGISTERS_20_31_port, B2 => n4596, ZN => n3871);
   U2046 : NOR2_X1 port map( A1 => n3874, A2 => n3883, ZN => n4395);
   U2047 : CLKBUF_X1 port map( A => n4395, Z => n4613);
   U2048 : NAND2_X1 port map( A1 => ADD_RD1(1), A2 => n3867, ZN => n3885);
   U2049 : NOR2_X1 port map( A1 => n3875, A2 => n3885, ZN => n4390);
   U2050 : CLKBUF_X1 port map( A => n4390, Z => n4601);
   U2051 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n4613, B1 => 
                           REGISTERS_26_31_port, B2 => n4601, ZN => n3870);
   U2052 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n3873, 
                           ZN => n3886);
   U2053 : NOR2_X1 port map( A1 => n3874, A2 => n3886, ZN => n4600);
   U2054 : CLKBUF_X1 port map( A => n4600, Z => n4570);
   U2055 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => 
                           ADD_RD1(2), ZN => n3887);
   U2056 : NOR2_X1 port map( A1 => n3874, A2 => n3887, ZN => n4420);
   U2057 : CLKBUF_X1 port map( A => n4420, Z => n4610);
   U2058 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n4570, B1 => 
                           REGISTERS_23_31_port, B2 => n4610, ZN => n3869);
   U2059 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => n3872, 
                           ZN => n3884);
   U2060 : NOR2_X1 port map( A1 => n3874, A2 => n3884, ZN => n4541);
   U2061 : NOR2_X1 port map( A1 => n3874, A2 => n3885, ZN => n4540);
   U2062 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n4541, B1 => 
                           REGISTERS_18_31_port, B2 => n4540, ZN => n3868);
   U2063 : NAND4_X1 port map( A1 => n3871, A2 => n3870, A3 => n3869, A4 => 
                           n3868, ZN => n3881);
   U2064 : NOR2_X1 port map( A1 => n3875, A2 => n3911, ZN => n4539);
   U2065 : CLKBUF_X1 port map( A => n4539, Z => n4595);
   U2066 : NOR2_X1 port map( A1 => n3875, A2 => n3887, ZN => n4571);
   U2067 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n4595, B1 => 
                           REGISTERS_31_31_port, B2 => n4571, ZN => n3879);
   U2068 : OR3_X1 port map( A1 => n3873, A2 => n3872, A3 => ADD_RD1(0), ZN => 
                           n4004);
   U2069 : NOR2_X1 port map( A1 => n4004, A2 => n3874, ZN => n4594);
   U2070 : NOR2_X1 port map( A1 => n4004, A2 => n3875, ZN => n4326);
   U2071 : CLKBUF_X1 port map( A => n4326, Z => n4609);
   U2072 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n4594, B1 => 
                           REGISTERS_30_31_port, B2 => n4609, ZN => n3878);
   U2073 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n3873, A3 => n3872, ZN =>
                           n3882);
   U2074 : NOR2_X1 port map( A1 => n3874, A2 => n3882, ZN => n4486);
   U2075 : CLKBUF_X1 port map( A => n4486, Z => n4608);
   U2076 : NOR2_X1 port map( A1 => n3875, A2 => n3884, ZN => n4349);
   U2077 : CLKBUF_X1 port map( A => n4349, Z => n4607);
   U2078 : AOI22_X1 port map( A1 => REGISTERS_17_31_port, A2 => n4608, B1 => 
                           REGISTERS_27_31_port, B2 => n4607, ZN => n3877);
   U2079 : NOR2_X1 port map( A1 => n3875, A2 => n3886, ZN => n4598);
   U2080 : NOR2_X1 port map( A1 => n3875, A2 => n3882, ZN => n4321);
   U2081 : CLKBUF_X1 port map( A => n4321, Z => n4606);
   U2082 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n4598, B1 => 
                           REGISTERS_25_31_port, B2 => n4606, ZN => n3876);
   U2083 : NAND4_X1 port map( A1 => n3879, A2 => n3878, A3 => n3877, A4 => 
                           n3876, ZN => n3880);
   U2084 : NOR2_X1 port map( A1 => n3881, A2 => n3880, ZN => n3900);
   U2085 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n4593, 
                           ZN => n4644);
   U2086 : CLKBUF_X1 port map( A => n4644, Z => n4459);
   U2087 : INV_X1 port map( A => n3882, ZN => n4633);
   U2088 : CLKBUF_X1 port map( A => n4633, Z => n4556);
   U2089 : INV_X1 port map( A => n3883, ZN => n4634);
   U2090 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n4556, B1 => 
                           REGISTERS_0_31_port, B2 => n4634, ZN => n3891);
   U2091 : INV_X1 port map( A => n3884, ZN => n4630);
   U2092 : CLKBUF_X1 port map( A => n4630, Z => n4548);
   U2093 : INV_X1 port map( A => n3885, ZN => n4579);
   U2094 : CLKBUF_X1 port map( A => n4579, Z => n4501);
   U2095 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n4548, B1 => 
                           REGISTERS_2_31_port, B2 => n4501, ZN => n3890);
   U2096 : INV_X1 port map( A => n3911, ZN => n4636);
   U2097 : INV_X1 port map( A => n3886, ZN => n4557);
   U2098 : CLKBUF_X1 port map( A => n4557, Z => n4550);
   U2099 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n4636, B1 => 
                           REGISTERS_5_31_port, B2 => n4550, ZN => n3889);
   U2100 : INV_X1 port map( A => n3887, ZN => n4635);
   U2101 : CLKBUF_X1 port map( A => n4635, Z => n4624);
   U2102 : INV_X1 port map( A => n4004, ZN => n4629);
   U2103 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n4624, B1 => 
                           REGISTERS_6_31_port, B2 => n4629, ZN => n3888);
   U2104 : NAND4_X1 port map( A1 => n3891, A2 => n3890, A3 => n3889, A4 => 
                           n3888, ZN => n3898);
   U2105 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n3892, A3 => n4593, ZN => 
                           n4642);
   U2106 : CLKBUF_X1 port map( A => n4642, Z => n4481);
   U2107 : CLKBUF_X1 port map( A => n4557, Z => n4632);
   U2108 : AOI22_X1 port map( A1 => REGISTERS_13_31_port, A2 => n4632, B1 => 
                           REGISTERS_10_31_port, B2 => n4501, ZN => n3896);
   U2109 : CLKBUF_X1 port map( A => n4634, Z => n4580);
   U2110 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n4580, B1 => 
                           REGISTERS_14_31_port, B2 => n4629, ZN => n3895);
   U2111 : INV_X1 port map( A => n3911, ZN => n4555);
   U2112 : CLKBUF_X1 port map( A => n4633, Z => n4621);
   U2113 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n4555, B1 => 
                           REGISTERS_9_31_port, B2 => n4621, ZN => n3894);
   U2114 : CLKBUF_X1 port map( A => n4630, Z => n4623);
   U2115 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n4624, B1 => 
                           REGISTERS_11_31_port, B2 => n4623, ZN => n3893);
   U2116 : NAND4_X1 port map( A1 => n3896, A2 => n3895, A3 => n3894, A4 => 
                           n3893, ZN => n3897);
   U2117 : AOI22_X1 port map( A1 => n4459, A2 => n3898, B1 => n4481, B2 => 
                           n3897, ZN => n3899);
   U2118 : OAI21_X1 port map( B1 => n4593, B2 => n3900, A => n3899, ZN => N416)
                           ;
   U2119 : AOI22_X1 port map( A1 => REGISTERS_25_30_port, A2 => n4606, B1 => 
                           REGISTERS_31_30_port, B2 => n4571, ZN => n3904);
   U2120 : CLKBUF_X1 port map( A => n4598, Z => n4572);
   U2121 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n4572, B1 => 
                           REGISTERS_19_30_port, B2 => n4541, ZN => n3903);
   U2122 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n4607, B1 => 
                           REGISTERS_21_30_port, B2 => n4600, ZN => n3902);
   U2123 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n4612, B1 => 
                           REGISTERS_22_30_port, B2 => n4594, ZN => n3901);
   U2124 : NAND4_X1 port map( A1 => n3904, A2 => n3903, A3 => n3902, A4 => 
                           n3901, ZN => n3910);
   U2125 : AOI22_X1 port map( A1 => REGISTERS_17_30_port, A2 => n4608, B1 => 
                           REGISTERS_28_30_port, B2 => n4539, ZN => n3908);
   U2126 : AOI22_X1 port map( A1 => REGISTERS_26_30_port, A2 => n4601, B1 => 
                           REGISTERS_16_30_port, B2 => n4613, ZN => n3907);
   U2127 : AOI22_X1 port map( A1 => REGISTERS_23_30_port, A2 => n4610, B1 => 
                           REGISTERS_20_30_port, B2 => n4415, ZN => n3906);
   U2128 : CLKBUF_X1 port map( A => n4540, Z => n4597);
   U2129 : AOI22_X1 port map( A1 => REGISTERS_18_30_port, A2 => n4597, B1 => 
                           REGISTERS_30_30_port, B2 => n4609, ZN => n3905);
   U2130 : NAND4_X1 port map( A1 => n3908, A2 => n3907, A3 => n3906, A4 => 
                           n3905, ZN => n3909);
   U2131 : NOR2_X1 port map( A1 => n3910, A2 => n3909, ZN => n3923);
   U2132 : INV_X1 port map( A => n4004, ZN => n4622);
   U2133 : CLKBUF_X1 port map( A => n4635, Z => n4522);
   U2134 : AOI22_X1 port map( A1 => REGISTERS_6_30_port, A2 => n4622, B1 => 
                           REGISTERS_7_30_port, B2 => n4522, ZN => n3915);
   U2135 : CLKBUF_X1 port map( A => n4579, Z => n4631);
   U2136 : AOI22_X1 port map( A1 => REGISTERS_2_30_port, A2 => n4631, B1 => 
                           REGISTERS_3_30_port, B2 => n4630, ZN => n3914);
   U2137 : INV_X1 port map( A => n3911, ZN => n4549);
   U2138 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n4633, B1 => 
                           REGISTERS_4_30_port, B2 => n4549, ZN => n3913);
   U2139 : CLKBUF_X1 port map( A => n4634, Z => n4620);
   U2140 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n4632, B1 => 
                           REGISTERS_0_30_port, B2 => n4620, ZN => n3912);
   U2141 : NAND4_X1 port map( A1 => n3915, A2 => n3914, A3 => n3913, A4 => 
                           n3912, ZN => n3921);
   U2142 : AOI22_X1 port map( A1 => REGISTERS_14_30_port, A2 => n4622, B1 => 
                           REGISTERS_13_30_port, B2 => n4557, ZN => n3919);
   U2143 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n4556, B1 => 
                           REGISTERS_12_30_port, B2 => n4636, ZN => n3918);
   U2144 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n4580, B1 => 
                           REGISTERS_15_30_port, B2 => n4522, ZN => n3917);
   U2145 : AOI22_X1 port map( A1 => REGISTERS_10_30_port, A2 => n4631, B1 => 
                           REGISTERS_11_30_port, B2 => n4623, ZN => n3916);
   U2146 : NAND4_X1 port map( A1 => n3919, A2 => n3918, A3 => n3917, A4 => 
                           n3916, ZN => n3920);
   U2147 : AOI22_X1 port map( A1 => n4459, A2 => n3921, B1 => n4481, B2 => 
                           n3920, ZN => n3922);
   U2148 : OAI21_X1 port map( B1 => n4593, B2 => n3923, A => n3922, ZN => N415)
                           ;
   U2149 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n4595, B1 => 
                           REGISTERS_21_29_port, B2 => n4600, ZN => n3927);
   U2150 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n4572, B1 => 
                           REGISTERS_25_29_port, B2 => n4321, ZN => n3926);
   U2151 : CLKBUF_X1 port map( A => n4541, Z => n4599);
   U2152 : AOI22_X1 port map( A1 => REGISTERS_19_29_port, A2 => n4599, B1 => 
                           REGISTERS_17_29_port, B2 => n4608, ZN => n3925);
   U2153 : AOI22_X1 port map( A1 => REGISTERS_18_29_port, A2 => n4597, B1 => 
                           REGISTERS_20_29_port, B2 => n4415, ZN => n3924);
   U2154 : NAND4_X1 port map( A1 => n3927, A2 => n3926, A3 => n3925, A4 => 
                           n3924, ZN => n3933);
   U2155 : CLKBUF_X1 port map( A => n4594, Z => n4510);
   U2156 : AOI22_X1 port map( A1 => REGISTERS_22_29_port, A2 => n4510, B1 => 
                           REGISTERS_26_29_port, B2 => n4601, ZN => n3931);
   U2157 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n4607, B1 => 
                           REGISTERS_24_29_port, B2 => n4612, ZN => n3930);
   U2158 : CLKBUF_X1 port map( A => n4571, Z => n4611);
   U2159 : AOI22_X1 port map( A1 => REGISTERS_31_29_port, A2 => n4611, B1 => 
                           REGISTERS_30_29_port, B2 => n4326, ZN => n3929);
   U2160 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n4610, B1 => 
                           REGISTERS_16_29_port, B2 => n4395, ZN => n3928);
   U2161 : NAND4_X1 port map( A1 => n3931, A2 => n3930, A3 => n3929, A4 => 
                           n3928, ZN => n3932);
   U2162 : NOR2_X1 port map( A1 => n3933, A2 => n3932, ZN => n3945);
   U2163 : AOI22_X1 port map( A1 => REGISTERS_2_29_port, A2 => n4631, B1 => 
                           REGISTERS_7_29_port, B2 => n4522, ZN => n3937);
   U2164 : AOI22_X1 port map( A1 => REGISTERS_6_29_port, A2 => n4622, B1 => 
                           REGISTERS_5_29_port, B2 => n4550, ZN => n3936);
   U2165 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n4630, B1 => 
                           REGISTERS_4_29_port, B2 => n4636, ZN => n3935);
   U2166 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n4580, B1 => 
                           REGISTERS_1_29_port, B2 => n4621, ZN => n3934);
   U2167 : NAND4_X1 port map( A1 => n3937, A2 => n3936, A3 => n3935, A4 => 
                           n3934, ZN => n3943);
   U2168 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n4623, B1 => 
                           REGISTERS_10_29_port, B2 => n4501, ZN => n3941);
   U2169 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n4555, B1 => 
                           REGISTERS_8_29_port, B2 => n4620, ZN => n3940);
   U2170 : AOI22_X1 port map( A1 => REGISTERS_14_29_port, A2 => n4622, B1 => 
                           REGISTERS_9_29_port, B2 => n4633, ZN => n3939);
   U2171 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n4635, B1 => 
                           REGISTERS_13_29_port, B2 => n4550, ZN => n3938);
   U2172 : NAND4_X1 port map( A1 => n3941, A2 => n3940, A3 => n3939, A4 => 
                           n3938, ZN => n3942);
   U2173 : AOI22_X1 port map( A1 => n4459, A2 => n3943, B1 => n4481, B2 => 
                           n3942, ZN => n3944);
   U2174 : OAI21_X1 port map( B1 => n4593, B2 => n3945, A => n3944, ZN => N414)
                           ;
   U2175 : AOI22_X1 port map( A1 => REGISTERS_17_28_port, A2 => n4608, B1 => 
                           REGISTERS_25_28_port, B2 => n4321, ZN => n3949);
   U2176 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n4613, B1 => 
                           REGISTERS_28_28_port, B2 => n4539, ZN => n3948);
   U2177 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n4607, B1 => 
                           REGISTERS_21_28_port, B2 => n4600, ZN => n3947);
   U2178 : AOI22_X1 port map( A1 => REGISTERS_18_28_port, A2 => n4597, B1 => 
                           REGISTERS_19_28_port, B2 => n4599, ZN => n3946);
   U2179 : NAND4_X1 port map( A1 => n3949, A2 => n3948, A3 => n3947, A4 => 
                           n3946, ZN => n3955);
   U2180 : AOI22_X1 port map( A1 => REGISTERS_30_28_port, A2 => n4609, B1 => 
                           REGISTERS_31_28_port, B2 => n4571, ZN => n3953);
   U2181 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n4612, B1 => 
                           REGISTERS_26_28_port, B2 => n4390, ZN => n3952);
   U2182 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n4596, B1 => 
                           REGISTERS_29_28_port, B2 => n4598, ZN => n3951);
   U2183 : AOI22_X1 port map( A1 => REGISTERS_23_28_port, A2 => n4610, B1 => 
                           REGISTERS_22_28_port, B2 => n4594, ZN => n3950);
   U2184 : NAND4_X1 port map( A1 => n3953, A2 => n3952, A3 => n3951, A4 => 
                           n3950, ZN => n3954);
   U2185 : NOR2_X1 port map( A1 => n3955, A2 => n3954, ZN => n3967);
   U2186 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n4549, B1 => 
                           REGISTERS_0_28_port, B2 => n4620, ZN => n3959);
   U2187 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n4632, B1 => 
                           REGISTERS_2_28_port, B2 => n4501, ZN => n3958);
   U2188 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n4630, B1 => 
                           REGISTERS_1_28_port, B2 => n4633, ZN => n3957);
   U2189 : AOI22_X1 port map( A1 => REGISTERS_6_28_port, A2 => n4622, B1 => 
                           REGISTERS_7_28_port, B2 => n4522, ZN => n3956);
   U2190 : NAND4_X1 port map( A1 => n3959, A2 => n3958, A3 => n3957, A4 => 
                           n3956, ZN => n3965);
   U2191 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n4632, B1 => 
                           REGISTERS_14_28_port, B2 => n4629, ZN => n3963);
   U2192 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n4630, B1 => 
                           REGISTERS_10_28_port, B2 => n4501, ZN => n3962);
   U2193 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n4635, B1 => 
                           REGISTERS_8_28_port, B2 => n4620, ZN => n3961);
   U2194 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n4621, B1 => 
                           REGISTERS_12_28_port, B2 => n4636, ZN => n3960);
   U2195 : NAND4_X1 port map( A1 => n3963, A2 => n3962, A3 => n3961, A4 => 
                           n3960, ZN => n3964);
   U2196 : AOI22_X1 port map( A1 => n4459, A2 => n3965, B1 => n4481, B2 => 
                           n3964, ZN => n3966);
   U2197 : OAI21_X1 port map( B1 => n4593, B2 => n3967, A => n3966, ZN => N413)
                           ;
   U2198 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n4612, B1 => 
                           REGISTERS_19_27_port, B2 => n4599, ZN => n3971);
   U2199 : AOI22_X1 port map( A1 => REGISTERS_21_27_port, A2 => n4570, B1 => 
                           REGISTERS_17_27_port, B2 => n4486, ZN => n3970);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_25_27_port, A2 => n4606, B1 => 
                           REGISTERS_20_27_port, B2 => n4415, ZN => n3969);
   U2201 : AOI22_X1 port map( A1 => REGISTERS_18_27_port, A2 => n4597, B1 => 
                           REGISTERS_16_27_port, B2 => n4395, ZN => n3968);
   U2202 : NAND4_X1 port map( A1 => n3971, A2 => n3970, A3 => n3969, A4 => 
                           n3968, ZN => n3977);
   U2203 : AOI22_X1 port map( A1 => REGISTERS_23_27_port, A2 => n4610, B1 => 
                           REGISTERS_30_27_port, B2 => n4326, ZN => n3975);
   U2204 : AOI22_X1 port map( A1 => REGISTERS_31_27_port, A2 => n4611, B1 => 
                           REGISTERS_28_27_port, B2 => n4539, ZN => n3974);
   U2205 : AOI22_X1 port map( A1 => REGISTERS_22_27_port, A2 => n4510, B1 => 
                           REGISTERS_29_27_port, B2 => n4572, ZN => n3973);
   U2206 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n4607, B1 => 
                           REGISTERS_26_27_port, B2 => n4390, ZN => n3972);
   U2207 : NAND4_X1 port map( A1 => n3975, A2 => n3974, A3 => n3973, A4 => 
                           n3972, ZN => n3976);
   U2208 : NOR2_X1 port map( A1 => n3977, A2 => n3976, ZN => n3989);
   U2209 : AOI22_X1 port map( A1 => REGISTERS_1_27_port, A2 => n4633, B1 => 
                           REGISTERS_6_27_port, B2 => n4629, ZN => n3981);
   U2210 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n4624, B1 => 
                           REGISTERS_3_27_port, B2 => n4623, ZN => n3980);
   U2211 : AOI22_X1 port map( A1 => REGISTERS_2_27_port, A2 => n4631, B1 => 
                           REGISTERS_5_27_port, B2 => n4550, ZN => n3979);
   U2212 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n4580, B1 => 
                           REGISTERS_4_27_port, B2 => n4636, ZN => n3978);
   U2213 : NAND4_X1 port map( A1 => n3981, A2 => n3980, A3 => n3979, A4 => 
                           n3978, ZN => n3987);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n4548, B1 => 
                           REGISTERS_15_27_port, B2 => n4635, ZN => n3985);
   U2215 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n4580, B1 => 
                           REGISTERS_12_27_port, B2 => n4555, ZN => n3984);
   U2216 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n4633, B1 => 
                           REGISTERS_13_27_port, B2 => n4550, ZN => n3983);
   U2217 : AOI22_X1 port map( A1 => REGISTERS_14_27_port, A2 => n4622, B1 => 
                           REGISTERS_10_27_port, B2 => n4501, ZN => n3982);
   U2218 : NAND4_X1 port map( A1 => n3985, A2 => n3984, A3 => n3983, A4 => 
                           n3982, ZN => n3986);
   U2219 : AOI22_X1 port map( A1 => n4459, A2 => n3987, B1 => n4481, B2 => 
                           n3986, ZN => n3988);
   U2220 : OAI21_X1 port map( B1 => n4593, B2 => n3989, A => n3988, ZN => N412)
                           ;
   U2221 : AOI22_X1 port map( A1 => REGISTERS_31_26_port, A2 => n4611, B1 => 
                           REGISTERS_16_26_port, B2 => n4395, ZN => n3993);
   U2222 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n4607, B1 => 
                           REGISTERS_21_26_port, B2 => n4600, ZN => n3992);
   U2223 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n4612, B1 => 
                           REGISTERS_26_26_port, B2 => n4390, ZN => n3991);
   U2224 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n4572, B1 => 
                           REGISTERS_23_26_port, B2 => n4420, ZN => n3990);
   U2225 : NAND4_X1 port map( A1 => n3993, A2 => n3992, A3 => n3991, A4 => 
                           n3990, ZN => n3999);
   U2226 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n4595, B1 => 
                           REGISTERS_18_26_port, B2 => n4540, ZN => n3997);
   U2227 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n4608, B1 => 
                           REGISTERS_20_26_port, B2 => n4415, ZN => n3996);
   U2228 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n4599, B1 => 
                           REGISTERS_25_26_port, B2 => n4321, ZN => n3995);
   U2229 : AOI22_X1 port map( A1 => REGISTERS_30_26_port, A2 => n4609, B1 => 
                           REGISTERS_22_26_port, B2 => n4510, ZN => n3994);
   U2230 : NAND4_X1 port map( A1 => n3997, A2 => n3996, A3 => n3995, A4 => 
                           n3994, ZN => n3998);
   U2231 : NOR2_X1 port map( A1 => n3999, A2 => n3998, ZN => n4012);
   U2232 : AOI22_X1 port map( A1 => REGISTERS_1_26_port, A2 => n4556, B1 => 
                           REGISTERS_6_26_port, B2 => n4629, ZN => n4003);
   U2233 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n4548, B1 => 
                           REGISTERS_5_26_port, B2 => n4550, ZN => n4002);
   U2234 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n4580, B1 => 
                           REGISTERS_2_26_port, B2 => n4579, ZN => n4001);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n4635, B1 => 
                           REGISTERS_4_26_port, B2 => n4555, ZN => n4000);
   U2236 : NAND4_X1 port map( A1 => n4003, A2 => n4002, A3 => n4001, A4 => 
                           n4000, ZN => n4010);
   U2237 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n4630, B1 => 
                           REGISTERS_10_26_port, B2 => n4501, ZN => n4008);
   U2238 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n4635, B1 => 
                           REGISTERS_9_26_port, B2 => n4633, ZN => n4007);
   U2239 : AOI22_X1 port map( A1 => REGISTERS_13_26_port, A2 => n4632, B1 => 
                           REGISTERS_8_26_port, B2 => n4620, ZN => n4006);
   U2240 : INV_X1 port map( A => n4004, ZN => n4521);
   U2241 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n4549, B1 => 
                           REGISTERS_14_26_port, B2 => n4521, ZN => n4005);
   U2242 : NAND4_X1 port map( A1 => n4008, A2 => n4007, A3 => n4006, A4 => 
                           n4005, ZN => n4009);
   U2243 : AOI22_X1 port map( A1 => n4459, A2 => n4010, B1 => n4481, B2 => 
                           n4009, ZN => n4011);
   U2244 : OAI21_X1 port map( B1 => n4593, B2 => n4012, A => n4011, ZN => N411)
                           ;
   U2245 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n4595, B1 => 
                           REGISTERS_27_25_port, B2 => n4607, ZN => n4016);
   U2246 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n4570, B1 => 
                           REGISTERS_20_25_port, B2 => n4415, ZN => n4015);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n4599, B1 => 
                           REGISTERS_29_25_port, B2 => n4572, ZN => n4014);
   U2248 : AOI22_X1 port map( A1 => REGISTERS_31_25_port, A2 => n4611, B1 => 
                           REGISTERS_22_25_port, B2 => n4510, ZN => n4013);
   U2249 : NAND4_X1 port map( A1 => n4016, A2 => n4015, A3 => n4014, A4 => 
                           n4013, ZN => n4022);
   U2250 : AOI22_X1 port map( A1 => REGISTERS_18_25_port, A2 => n4597, B1 => 
                           REGISTERS_23_25_port, B2 => n4420, ZN => n4020);
   U2251 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n4608, B1 => 
                           REGISTERS_25_25_port, B2 => n4321, ZN => n4019);
   U2252 : AOI22_X1 port map( A1 => REGISTERS_30_25_port, A2 => n4609, B1 => 
                           REGISTERS_24_25_port, B2 => n4396, ZN => n4018);
   U2253 : AOI22_X1 port map( A1 => REGISTERS_26_25_port, A2 => n4601, B1 => 
                           REGISTERS_16_25_port, B2 => n4395, ZN => n4017);
   U2254 : NAND4_X1 port map( A1 => n4020, A2 => n4019, A3 => n4018, A4 => 
                           n4017, ZN => n4021);
   U2255 : NOR2_X1 port map( A1 => n4022, A2 => n4021, ZN => n4034);
   U2256 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n4556, B1 => 
                           REGISTERS_4_25_port, B2 => n4555, ZN => n4026);
   U2257 : AOI22_X1 port map( A1 => REGISTERS_3_25_port, A2 => n4548, B1 => 
                           REGISTERS_5_25_port, B2 => n4557, ZN => n4025);
   U2258 : AOI22_X1 port map( A1 => REGISTERS_2_25_port, A2 => n4631, B1 => 
                           REGISTERS_7_25_port, B2 => n4635, ZN => n4024);
   U2259 : AOI22_X1 port map( A1 => REGISTERS_6_25_port, A2 => n4622, B1 => 
                           REGISTERS_0_25_port, B2 => n4634, ZN => n4023);
   U2260 : NAND4_X1 port map( A1 => n4026, A2 => n4025, A3 => n4024, A4 => 
                           n4023, ZN => n4032);
   U2261 : AOI22_X1 port map( A1 => REGISTERS_14_25_port, A2 => n4622, B1 => 
                           REGISTERS_9_25_port, B2 => n4633, ZN => n4030);
   U2262 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n4624, B1 => 
                           REGISTERS_12_25_port, B2 => n4555, ZN => n4029);
   U2263 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n4630, B1 => 
                           REGISTERS_13_25_port, B2 => n4550, ZN => n4028);
   U2264 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n4580, B1 => 
                           REGISTERS_10_25_port, B2 => n4579, ZN => n4027);
   U2265 : NAND4_X1 port map( A1 => n4030, A2 => n4029, A3 => n4028, A4 => 
                           n4027, ZN => n4031);
   U2266 : AOI22_X1 port map( A1 => n4459, A2 => n4032, B1 => n4481, B2 => 
                           n4031, ZN => n4033);
   U2267 : OAI21_X1 port map( B1 => n4593, B2 => n4034, A => n4033, ZN => N410)
                           ;
   U2268 : AOI22_X1 port map( A1 => REGISTERS_30_24_port, A2 => n4609, B1 => 
                           REGISTERS_19_24_port, B2 => n4599, ZN => n4038);
   U2269 : AOI22_X1 port map( A1 => REGISTERS_18_24_port, A2 => n4597, B1 => 
                           REGISTERS_23_24_port, B2 => n4420, ZN => n4037);
   U2270 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n4596, B1 => 
                           REGISTERS_28_24_port, B2 => n4539, ZN => n4036);
   U2271 : AOI22_X1 port map( A1 => REGISTERS_22_24_port, A2 => n4510, B1 => 
                           REGISTERS_31_24_port, B2 => n4571, ZN => n4035);
   U2272 : NAND4_X1 port map( A1 => n4038, A2 => n4037, A3 => n4036, A4 => 
                           n4035, ZN => n4044);
   U2273 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n4613, B1 => 
                           REGISTERS_25_24_port, B2 => n4321, ZN => n4042);
   U2274 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n4570, B1 => 
                           REGISTERS_26_24_port, B2 => n4390, ZN => n4041);
   U2275 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n4607, B1 => 
                           REGISTERS_17_24_port, B2 => n4486, ZN => n4040);
   U2276 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n4572, B1 => 
                           REGISTERS_24_24_port, B2 => n4396, ZN => n4039);
   U2277 : NAND4_X1 port map( A1 => n4042, A2 => n4041, A3 => n4040, A4 => 
                           n4039, ZN => n4043);
   U2278 : NOR2_X1 port map( A1 => n4044, A2 => n4043, ZN => n4056);
   U2279 : AOI22_X1 port map( A1 => REGISTERS_1_24_port, A2 => n4556, B1 => 
                           REGISTERS_6_24_port, B2 => n4521, ZN => n4048);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n4623, B1 => 
                           REGISTERS_5_24_port, B2 => n4557, ZN => n4047);
   U2281 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n4635, B1 => 
                           REGISTERS_2_24_port, B2 => n4501, ZN => n4046);
   U2282 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n4549, B1 => 
                           REGISTERS_0_24_port, B2 => n4620, ZN => n4045);
   U2283 : NAND4_X1 port map( A1 => n4048, A2 => n4047, A3 => n4046, A4 => 
                           n4045, ZN => n4054);
   U2284 : AOI22_X1 port map( A1 => REGISTERS_10_24_port, A2 => n4631, B1 => 
                           REGISTERS_8_24_port, B2 => n4634, ZN => n4052);
   U2285 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n4548, B1 => 
                           REGISTERS_13_24_port, B2 => n4550, ZN => n4051);
   U2286 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n4636, B1 => 
                           REGISTERS_15_24_port, B2 => n4635, ZN => n4050);
   U2287 : AOI22_X1 port map( A1 => REGISTERS_9_24_port, A2 => n4633, B1 => 
                           REGISTERS_14_24_port, B2 => n4521, ZN => n4049);
   U2288 : NAND4_X1 port map( A1 => n4052, A2 => n4051, A3 => n4050, A4 => 
                           n4049, ZN => n4053);
   U2289 : AOI22_X1 port map( A1 => n4459, A2 => n4054, B1 => n4481, B2 => 
                           n4053, ZN => n4055);
   U2290 : OAI21_X1 port map( B1 => n4593, B2 => n4056, A => n4055, ZN => N409)
                           ;
   U2291 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n4572, B1 => 
                           REGISTERS_31_23_port, B2 => n4611, ZN => n4060);
   U2292 : AOI22_X1 port map( A1 => REGISTERS_22_23_port, A2 => n4510, B1 => 
                           REGISTERS_23_23_port, B2 => n4420, ZN => n4059);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_18_23_port, A2 => n4540, B1 => 
                           REGISTERS_27_23_port, B2 => n4349, ZN => n4058);
   U2294 : AOI22_X1 port map( A1 => REGISTERS_19_23_port, A2 => n4599, B1 => 
                           REGISTERS_30_23_port, B2 => n4326, ZN => n4057);
   U2295 : NAND4_X1 port map( A1 => n4060, A2 => n4059, A3 => n4058, A4 => 
                           n4057, ZN => n4066);
   U2296 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n4596, B1 => 
                           REGISTERS_25_23_port, B2 => n4321, ZN => n4064);
   U2297 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n4570, B1 => 
                           REGISTERS_26_23_port, B2 => n4390, ZN => n4063);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n4608, B1 => 
                           REGISTERS_24_23_port, B2 => n4396, ZN => n4062);
   U2299 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n4595, B1 => 
                           REGISTERS_16_23_port, B2 => n4613, ZN => n4061);
   U2300 : NAND4_X1 port map( A1 => n4064, A2 => n4063, A3 => n4062, A4 => 
                           n4061, ZN => n4065);
   U2301 : NOR2_X1 port map( A1 => n4066, A2 => n4065, ZN => n4078);
   U2302 : AOI22_X1 port map( A1 => REGISTERS_1_23_port, A2 => n4633, B1 => 
                           REGISTERS_0_23_port, B2 => n4620, ZN => n4070);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n4557, B1 => 
                           REGISTERS_4_23_port, B2 => n4549, ZN => n4069);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n4522, B1 => 
                           REGISTERS_3_23_port, B2 => n4630, ZN => n4068);
   U2305 : AOI22_X1 port map( A1 => REGISTERS_2_23_port, A2 => n4579, B1 => 
                           REGISTERS_6_23_port, B2 => n4521, ZN => n4067);
   U2306 : NAND4_X1 port map( A1 => n4070, A2 => n4069, A3 => n4068, A4 => 
                           n4067, ZN => n4076);
   U2307 : AOI22_X1 port map( A1 => REGISTERS_14_23_port, A2 => n4622, B1 => 
                           REGISTERS_8_23_port, B2 => n4634, ZN => n4074);
   U2308 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n4632, B1 => 
                           REGISTERS_12_23_port, B2 => n4555, ZN => n4073);
   U2309 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n4623, B1 => 
                           REGISTERS_15_23_port, B2 => n4522, ZN => n4072);
   U2310 : AOI22_X1 port map( A1 => REGISTERS_9_23_port, A2 => n4621, B1 => 
                           REGISTERS_10_23_port, B2 => n4579, ZN => n4071);
   U2311 : NAND4_X1 port map( A1 => n4074, A2 => n4073, A3 => n4072, A4 => 
                           n4071, ZN => n4075);
   U2312 : AOI22_X1 port map( A1 => n4459, A2 => n4076, B1 => n4481, B2 => 
                           n4075, ZN => n4077);
   U2313 : OAI21_X1 port map( B1 => n4647, B2 => n4078, A => n4077, ZN => N408)
                           ;
   U2314 : AOI22_X1 port map( A1 => REGISTERS_21_22_port, A2 => n4570, B1 => 
                           REGISTERS_28_22_port, B2 => n4595, ZN => n4082);
   U2315 : AOI22_X1 port map( A1 => REGISTERS_31_22_port, A2 => n4611, B1 => 
                           REGISTERS_30_22_port, B2 => n4326, ZN => n4081);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n4613, B1 => 
                           REGISTERS_27_22_port, B2 => n4349, ZN => n4080);
   U2317 : AOI22_X1 port map( A1 => REGISTERS_25_22_port, A2 => n4606, B1 => 
                           REGISTERS_22_22_port, B2 => n4594, ZN => n4079);
   U2318 : NAND4_X1 port map( A1 => n4082, A2 => n4081, A3 => n4080, A4 => 
                           n4079, ZN => n4088);
   U2319 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n4612, B1 => 
                           REGISTERS_26_22_port, B2 => n4390, ZN => n4086);
   U2320 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n4596, B1 => 
                           REGISTERS_18_22_port, B2 => n4597, ZN => n4085);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n4598, B1 => 
                           REGISTERS_17_22_port, B2 => n4486, ZN => n4084);
   U2322 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n4599, B1 => 
                           REGISTERS_23_22_port, B2 => n4420, ZN => n4083);
   U2323 : NAND4_X1 port map( A1 => n4086, A2 => n4085, A3 => n4084, A4 => 
                           n4083, ZN => n4087);
   U2324 : NOR2_X1 port map( A1 => n4088, A2 => n4087, ZN => n4100);
   U2325 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n4548, B1 => 
                           REGISTERS_0_22_port, B2 => n4620, ZN => n4092);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n4636, B1 => 
                           REGISTERS_5_22_port, B2 => n4557, ZN => n4091);
   U2327 : AOI22_X1 port map( A1 => REGISTERS_6_22_port, A2 => n4622, B1 => 
                           REGISTERS_2_22_port, B2 => n4501, ZN => n4090);
   U2328 : AOI22_X1 port map( A1 => REGISTERS_1_22_port, A2 => n4621, B1 => 
                           REGISTERS_7_22_port, B2 => n4522, ZN => n4089);
   U2329 : NAND4_X1 port map( A1 => n4092, A2 => n4091, A3 => n4090, A4 => 
                           n4089, ZN => n4098);
   U2330 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n4555, B1 => 
                           REGISTERS_8_22_port, B2 => n4634, ZN => n4096);
   U2331 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n4522, B1 => 
                           REGISTERS_9_22_port, B2 => n4621, ZN => n4095);
   U2332 : AOI22_X1 port map( A1 => REGISTERS_13_22_port, A2 => n4557, B1 => 
                           REGISTERS_10_22_port, B2 => n4579, ZN => n4094);
   U2333 : AOI22_X1 port map( A1 => REGISTERS_11_22_port, A2 => n4623, B1 => 
                           REGISTERS_14_22_port, B2 => n4521, ZN => n4093);
   U2334 : NAND4_X1 port map( A1 => n4096, A2 => n4095, A3 => n4094, A4 => 
                           n4093, ZN => n4097);
   U2335 : AOI22_X1 port map( A1 => n4459, A2 => n4098, B1 => n4481, B2 => 
                           n4097, ZN => n4099);
   U2336 : OAI21_X1 port map( B1 => n4647, B2 => n4100, A => n4099, ZN => N407)
                           ;
   U2337 : AOI22_X1 port map( A1 => REGISTERS_27_21_port, A2 => n4607, B1 => 
                           REGISTERS_20_21_port, B2 => n4415, ZN => n4104);
   U2338 : AOI22_X1 port map( A1 => REGISTERS_23_21_port, A2 => n4610, B1 => 
                           REGISTERS_18_21_port, B2 => n4597, ZN => n4103);
   U2339 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n4599, B1 => 
                           REGISTERS_30_21_port, B2 => n4326, ZN => n4102);
   U2340 : AOI22_X1 port map( A1 => REGISTERS_21_21_port, A2 => n4570, B1 => 
                           REGISTERS_17_21_port, B2 => n4486, ZN => n4101);
   U2341 : NAND4_X1 port map( A1 => n4104, A2 => n4103, A3 => n4102, A4 => 
                           n4101, ZN => n4110);
   U2342 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n4510, B1 => 
                           REGISTERS_26_21_port, B2 => n4390, ZN => n4108);
   U2343 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n4598, B1 => 
                           REGISTERS_25_21_port, B2 => n4321, ZN => n4107);
   U2344 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n4595, B1 => 
                           REGISTERS_31_21_port, B2 => n4611, ZN => n4106);
   U2345 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n4612, B1 => 
                           REGISTERS_16_21_port, B2 => n4395, ZN => n4105);
   U2346 : NAND4_X1 port map( A1 => n4108, A2 => n4107, A3 => n4106, A4 => 
                           n4105, ZN => n4109);
   U2347 : NOR2_X1 port map( A1 => n4110, A2 => n4109, ZN => n4122);
   U2348 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n4635, B1 => 
                           REGISTERS_5_21_port, B2 => n4550, ZN => n4114);
   U2349 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n4580, B1 => 
                           REGISTERS_3_21_port, B2 => n4630, ZN => n4113);
   U2350 : AOI22_X1 port map( A1 => REGISTERS_6_21_port, A2 => n4622, B1 => 
                           REGISTERS_4_21_port, B2 => n4555, ZN => n4112);
   U2351 : AOI22_X1 port map( A1 => REGISTERS_2_21_port, A2 => n4501, B1 => 
                           REGISTERS_1_21_port, B2 => n4633, ZN => n4111);
   U2352 : NAND4_X1 port map( A1 => n4114, A2 => n4113, A3 => n4112, A4 => 
                           n4111, ZN => n4120);
   U2353 : AOI22_X1 port map( A1 => REGISTERS_14_21_port, A2 => n4521, B1 => 
                           REGISTERS_13_21_port, B2 => n4557, ZN => n4118);
   U2354 : AOI22_X1 port map( A1 => REGISTERS_10_21_port, A2 => n4501, B1 => 
                           REGISTERS_15_21_port, B2 => n4522, ZN => n4117);
   U2355 : AOI22_X1 port map( A1 => REGISTERS_9_21_port, A2 => n4621, B1 => 
                           REGISTERS_11_21_port, B2 => n4623, ZN => n4116);
   U2356 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n4580, B1 => 
                           REGISTERS_12_21_port, B2 => n4555, ZN => n4115);
   U2357 : NAND4_X1 port map( A1 => n4118, A2 => n4117, A3 => n4116, A4 => 
                           n4115, ZN => n4119);
   U2358 : AOI22_X1 port map( A1 => n4459, A2 => n4120, B1 => n4481, B2 => 
                           n4119, ZN => n4121);
   U2359 : OAI21_X1 port map( B1 => n4647, B2 => n4122, A => n4121, ZN => N406)
                           ;
   U2360 : AOI22_X1 port map( A1 => REGISTERS_31_20_port, A2 => n4611, B1 => 
                           REGISTERS_23_20_port, B2 => n4420, ZN => n4126);
   U2361 : AOI22_X1 port map( A1 => REGISTERS_22_20_port, A2 => n4510, B1 => 
                           REGISTERS_17_20_port, B2 => n4486, ZN => n4125);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n4595, B1 => 
                           REGISTERS_24_20_port, B2 => n4396, ZN => n4124);
   U2363 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n4349, B1 => 
                           REGISTERS_25_20_port, B2 => n4321, ZN => n4123);
   U2364 : NAND4_X1 port map( A1 => n4126, A2 => n4125, A3 => n4124, A4 => 
                           n4123, ZN => n4132);
   U2365 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n4572, B1 => 
                           REGISTERS_30_20_port, B2 => n4326, ZN => n4130);
   U2366 : AOI22_X1 port map( A1 => REGISTERS_18_20_port, A2 => n4540, B1 => 
                           REGISTERS_21_20_port, B2 => n4600, ZN => n4129);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_19_20_port, A2 => n4541, B1 => 
                           REGISTERS_26_20_port, B2 => n4390, ZN => n4128);
   U2368 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n4596, B1 => 
                           REGISTERS_16_20_port, B2 => n4395, ZN => n4127);
   U2369 : NAND4_X1 port map( A1 => n4130, A2 => n4129, A3 => n4128, A4 => 
                           n4127, ZN => n4131);
   U2370 : NOR2_X1 port map( A1 => n4132, A2 => n4131, ZN => n4144);
   U2371 : AOI22_X1 port map( A1 => REGISTERS_6_20_port, A2 => n4629, B1 => 
                           REGISTERS_2_20_port, B2 => n4501, ZN => n4136);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n4522, B1 => 
                           REGISTERS_3_20_port, B2 => n4548, ZN => n4135);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n4556, B1 => 
                           REGISTERS_4_20_port, B2 => n4555, ZN => n4134);
   U2374 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n4620, B1 => 
                           REGISTERS_5_20_port, B2 => n4550, ZN => n4133);
   U2375 : NAND4_X1 port map( A1 => n4136, A2 => n4135, A3 => n4134, A4 => 
                           n4133, ZN => n4142);
   U2376 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n4580, B1 => 
                           REGISTERS_12_20_port, B2 => n4555, ZN => n4140);
   U2377 : AOI22_X1 port map( A1 => REGISTERS_15_20_port, A2 => n4522, B1 => 
                           REGISTERS_14_20_port, B2 => n4521, ZN => n4139);
   U2378 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n4633, B1 => 
                           REGISTERS_10_20_port, B2 => n4579, ZN => n4138);
   U2379 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n4548, B1 => 
                           REGISTERS_13_20_port, B2 => n4557, ZN => n4137);
   U2380 : NAND4_X1 port map( A1 => n4140, A2 => n4139, A3 => n4138, A4 => 
                           n4137, ZN => n4141);
   U2381 : AOI22_X1 port map( A1 => n4459, A2 => n4142, B1 => n4642, B2 => 
                           n4141, ZN => n4143);
   U2382 : OAI21_X1 port map( B1 => n4647, B2 => n4144, A => n4143, ZN => N405)
                           ;
   U2383 : AOI22_X1 port map( A1 => REGISTERS_22_19_port, A2 => n4594, B1 => 
                           REGISTERS_31_19_port, B2 => n4611, ZN => n4148);
   U2384 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n4610, B1 => 
                           REGISTERS_18_19_port, B2 => n4597, ZN => n4147);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_19_19_port, A2 => n4541, B1 => 
                           REGISTERS_27_19_port, B2 => n4349, ZN => n4146);
   U2386 : AOI22_X1 port map( A1 => REGISTERS_21_19_port, A2 => n4570, B1 => 
                           REGISTERS_16_19_port, B2 => n4395, ZN => n4145);
   U2387 : NAND4_X1 port map( A1 => n4148, A2 => n4147, A3 => n4146, A4 => 
                           n4145, ZN => n4154);
   U2388 : AOI22_X1 port map( A1 => REGISTERS_30_19_port, A2 => n4609, B1 => 
                           REGISTERS_29_19_port, B2 => n4572, ZN => n4152);
   U2389 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n4608, B1 => 
                           REGISTERS_25_19_port, B2 => n4606, ZN => n4151);
   U2390 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n4595, B1 => 
                           REGISTERS_20_19_port, B2 => n4415, ZN => n4150);
   U2391 : AOI22_X1 port map( A1 => REGISTERS_26_19_port, A2 => n4390, B1 => 
                           REGISTERS_24_19_port, B2 => n4396, ZN => n4149);
   U2392 : NAND4_X1 port map( A1 => n4152, A2 => n4151, A3 => n4150, A4 => 
                           n4149, ZN => n4153);
   U2393 : NOR2_X1 port map( A1 => n4154, A2 => n4153, ZN => n4166);
   U2394 : CLKBUF_X1 port map( A => n4644, Z => n4483);
   U2395 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n4635, B1 => 
                           REGISTERS_1_19_port, B2 => n4556, ZN => n4158);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n4550, B1 => 
                           REGISTERS_6_19_port, B2 => n4521, ZN => n4157);
   U2397 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n4580, B1 => 
                           REGISTERS_2_19_port, B2 => n4501, ZN => n4156);
   U2398 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n4549, B1 => 
                           REGISTERS_3_19_port, B2 => n4548, ZN => n4155);
   U2399 : NAND4_X1 port map( A1 => n4158, A2 => n4157, A3 => n4156, A4 => 
                           n4155, ZN => n4164);
   U2400 : AOI22_X1 port map( A1 => REGISTERS_14_19_port, A2 => n4622, B1 => 
                           REGISTERS_8_19_port, B2 => n4620, ZN => n4162);
   U2401 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n4549, B1 => 
                           REGISTERS_13_19_port, B2 => n4550, ZN => n4161);
   U2402 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n4522, B1 => 
                           REGISTERS_10_19_port, B2 => n4579, ZN => n4160);
   U2403 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n4630, B1 => 
                           REGISTERS_9_19_port, B2 => n4633, ZN => n4159);
   U2404 : NAND4_X1 port map( A1 => n4162, A2 => n4161, A3 => n4160, A4 => 
                           n4159, ZN => n4163);
   U2405 : AOI22_X1 port map( A1 => n4483, A2 => n4164, B1 => n4481, B2 => 
                           n4163, ZN => n4165);
   U2406 : OAI21_X1 port map( B1 => n4647, B2 => n4166, A => n4165, ZN => N404)
                           ;
   U2407 : AOI22_X1 port map( A1 => REGISTERS_19_18_port, A2 => n4599, B1 => 
                           REGISTERS_22_18_port, B2 => n4510, ZN => n4170);
   U2408 : AOI22_X1 port map( A1 => REGISTERS_26_18_port, A2 => n4390, B1 => 
                           REGISTERS_24_18_port, B2 => n4396, ZN => n4169);
   U2409 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n4539, B1 => 
                           REGISTERS_18_18_port, B2 => n4597, ZN => n4168);
   U2410 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n4420, B1 => 
                           REGISTERS_20_18_port, B2 => n4415, ZN => n4167);
   U2411 : NAND4_X1 port map( A1 => n4170, A2 => n4169, A3 => n4168, A4 => 
                           n4167, ZN => n4176);
   U2412 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n4349, B1 => 
                           REGISTERS_25_18_port, B2 => n4606, ZN => n4174);
   U2413 : AOI22_X1 port map( A1 => REGISTERS_30_18_port, A2 => n4326, B1 => 
                           REGISTERS_31_18_port, B2 => n4611, ZN => n4173);
   U2414 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n4395, B1 => 
                           REGISTERS_21_18_port, B2 => n4570, ZN => n4172);
   U2415 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n4486, B1 => 
                           REGISTERS_29_18_port, B2 => n4572, ZN => n4171);
   U2416 : NAND4_X1 port map( A1 => n4174, A2 => n4173, A3 => n4172, A4 => 
                           n4171, ZN => n4175);
   U2417 : NOR2_X1 port map( A1 => n4176, A2 => n4175, ZN => n4188);
   U2418 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n4621, B1 => 
                           REGISTERS_2_18_port, B2 => n4579, ZN => n4180);
   U2419 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n4620, B1 => 
                           REGISTERS_7_18_port, B2 => n4624, ZN => n4179);
   U2420 : AOI22_X1 port map( A1 => REGISTERS_6_18_port, A2 => n4521, B1 => 
                           REGISTERS_4_18_port, B2 => n4555, ZN => n4178);
   U2421 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n4632, B1 => 
                           REGISTERS_3_18_port, B2 => n4623, ZN => n4177);
   U2422 : NAND4_X1 port map( A1 => n4180, A2 => n4179, A3 => n4178, A4 => 
                           n4177, ZN => n4186);
   U2423 : AOI22_X1 port map( A1 => REGISTERS_14_18_port, A2 => n4521, B1 => 
                           REGISTERS_10_18_port, B2 => n4501, ZN => n4184);
   U2424 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n4624, B1 => 
                           REGISTERS_11_18_port, B2 => n4623, ZN => n4183);
   U2425 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n4556, B1 => 
                           REGISTERS_12_18_port, B2 => n4555, ZN => n4182);
   U2426 : AOI22_X1 port map( A1 => REGISTERS_13_18_port, A2 => n4550, B1 => 
                           REGISTERS_8_18_port, B2 => n4634, ZN => n4181);
   U2427 : NAND4_X1 port map( A1 => n4184, A2 => n4183, A3 => n4182, A4 => 
                           n4181, ZN => n4185);
   U2428 : AOI22_X1 port map( A1 => n4483, A2 => n4186, B1 => n4481, B2 => 
                           n4185, ZN => n4187);
   U2429 : OAI21_X1 port map( B1 => n4647, B2 => n4188, A => n4187, ZN => N403)
                           ;
   U2430 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n4571, B1 => 
                           REGISTERS_30_17_port, B2 => n4326, ZN => n4192);
   U2431 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n4420, B1 => 
                           REGISTERS_28_17_port, B2 => n4595, ZN => n4191);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_22_17_port, A2 => n4594, B1 => 
                           REGISTERS_27_17_port, B2 => n4349, ZN => n4190);
   U2433 : AOI22_X1 port map( A1 => REGISTERS_18_17_port, A2 => n4540, B1 => 
                           REGISTERS_25_17_port, B2 => n4606, ZN => n4189);
   U2434 : NAND4_X1 port map( A1 => n4192, A2 => n4191, A3 => n4190, A4 => 
                           n4189, ZN => n4198);
   U2435 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n4600, B1 => 
                           REGISTERS_17_17_port, B2 => n4486, ZN => n4196);
   U2436 : AOI22_X1 port map( A1 => REGISTERS_26_17_port, A2 => n4601, B1 => 
                           REGISTERS_16_17_port, B2 => n4395, ZN => n4195);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n4572, B1 => 
                           REGISTERS_19_17_port, B2 => n4599, ZN => n4194);
   U2438 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n4415, B1 => 
                           REGISTERS_24_17_port, B2 => n4396, ZN => n4193);
   U2439 : NAND4_X1 port map( A1 => n4196, A2 => n4195, A3 => n4194, A4 => 
                           n4193, ZN => n4197);
   U2440 : NOR2_X1 port map( A1 => n4198, A2 => n4197, ZN => n4210);
   U2441 : AOI22_X1 port map( A1 => REGISTERS_6_17_port, A2 => n4622, B1 => 
                           REGISTERS_1_17_port, B2 => n4621, ZN => n4202);
   U2442 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n4635, B1 => 
                           REGISTERS_5_17_port, B2 => n4557, ZN => n4201);
   U2443 : AOI22_X1 port map( A1 => REGISTERS_2_17_port, A2 => n4501, B1 => 
                           REGISTERS_3_17_port, B2 => n4630, ZN => n4200);
   U2444 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n4636, B1 => 
                           REGISTERS_0_17_port, B2 => n4620, ZN => n4199);
   U2445 : NAND4_X1 port map( A1 => n4202, A2 => n4201, A3 => n4200, A4 => 
                           n4199, ZN => n4208);
   U2446 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n4555, B1 => 
                           REGISTERS_8_17_port, B2 => n4634, ZN => n4206);
   U2447 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n4623, B1 => 
                           REGISTERS_9_17_port, B2 => n4556, ZN => n4205);
   U2448 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n4632, B1 => 
                           REGISTERS_14_17_port, B2 => n4521, ZN => n4204);
   U2449 : AOI22_X1 port map( A1 => REGISTERS_10_17_port, A2 => n4579, B1 => 
                           REGISTERS_15_17_port, B2 => n4522, ZN => n4203);
   U2450 : NAND4_X1 port map( A1 => n4206, A2 => n4205, A3 => n4204, A4 => 
                           n4203, ZN => n4207);
   U2451 : AOI22_X1 port map( A1 => n4483, A2 => n4208, B1 => n4481, B2 => 
                           n4207, ZN => n4209);
   U2452 : OAI21_X1 port map( B1 => n4647, B2 => n4210, A => n4209, ZN => N402)
                           ;
   U2453 : AOI22_X1 port map( A1 => REGISTERS_26_16_port, A2 => n4601, B1 => 
                           REGISTERS_23_16_port, B2 => n4420, ZN => n4214);
   U2454 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n4539, B1 => 
                           REGISTERS_27_16_port, B2 => n4349, ZN => n4213);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n4572, B1 => 
                           REGISTERS_25_16_port, B2 => n4606, ZN => n4212);
   U2456 : AOI22_X1 port map( A1 => REGISTERS_22_16_port, A2 => n4510, B1 => 
                           REGISTERS_30_16_port, B2 => n4326, ZN => n4211);
   U2457 : NAND4_X1 port map( A1 => n4214, A2 => n4213, A3 => n4212, A4 => 
                           n4211, ZN => n4220);
   U2458 : AOI22_X1 port map( A1 => REGISTERS_17_16_port, A2 => n4608, B1 => 
                           REGISTERS_24_16_port, B2 => n4396, ZN => n4218);
   U2459 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n4395, B1 => 
                           REGISTERS_31_16_port, B2 => n4611, ZN => n4217);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_18_16_port, A2 => n4597, B1 => 
                           REGISTERS_21_16_port, B2 => n4570, ZN => n4216);
   U2461 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n4599, B1 => 
                           REGISTERS_20_16_port, B2 => n4596, ZN => n4215);
   U2462 : NAND4_X1 port map( A1 => n4218, A2 => n4217, A3 => n4216, A4 => 
                           n4215, ZN => n4219);
   U2463 : NOR2_X1 port map( A1 => n4220, A2 => n4219, ZN => n4232);
   U2464 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n4620, B1 => 
                           REGISTERS_6_16_port, B2 => n4521, ZN => n4224);
   U2465 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n4522, B1 => 
                           REGISTERS_2_16_port, B2 => n4579, ZN => n4223);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_1_16_port, A2 => n4633, B1 => 
                           REGISTERS_4_16_port, B2 => n4555, ZN => n4222);
   U2467 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n4548, B1 => 
                           REGISTERS_5_16_port, B2 => n4557, ZN => n4221);
   U2468 : NAND4_X1 port map( A1 => n4224, A2 => n4223, A3 => n4222, A4 => 
                           n4221, ZN => n4230);
   U2469 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n4630, B1 => 
                           REGISTERS_13_16_port, B2 => n4550, ZN => n4228);
   U2470 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n4549, B1 => 
                           REGISTERS_8_16_port, B2 => n4634, ZN => n4227);
   U2471 : AOI22_X1 port map( A1 => REGISTERS_14_16_port, A2 => n4521, B1 => 
                           REGISTERS_15_16_port, B2 => n4635, ZN => n4226);
   U2472 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n4501, B1 => 
                           REGISTERS_9_16_port, B2 => n4621, ZN => n4225);
   U2473 : NAND4_X1 port map( A1 => n4228, A2 => n4227, A3 => n4226, A4 => 
                           n4225, ZN => n4229);
   U2474 : AOI22_X1 port map( A1 => n4483, A2 => n4230, B1 => n4481, B2 => 
                           n4229, ZN => n4231);
   U2475 : OAI21_X1 port map( B1 => n4647, B2 => n4232, A => n4231, ZN => N401)
                           ;
   U2476 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n4600, B1 => 
                           REGISTERS_24_15_port, B2 => n4612, ZN => n4236);
   U2477 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n4596, B1 => 
                           REGISTERS_29_15_port, B2 => n4572, ZN => n4235);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_18_15_port, A2 => n4597, B1 => 
                           REGISTERS_22_15_port, B2 => n4510, ZN => n4234);
   U2479 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n4571, B1 => 
                           REGISTERS_17_15_port, B2 => n4486, ZN => n4233);
   U2480 : NAND4_X1 port map( A1 => n4236, A2 => n4235, A3 => n4234, A4 => 
                           n4233, ZN => n4242);
   U2481 : AOI22_X1 port map( A1 => REGISTERS_27_15_port, A2 => n4607, B1 => 
                           REGISTERS_23_15_port, B2 => n4420, ZN => n4240);
   U2482 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n4613, B1 => 
                           REGISTERS_25_15_port, B2 => n4606, ZN => n4239);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_26_15_port, A2 => n4601, B1 => 
                           REGISTERS_28_15_port, B2 => n4595, ZN => n4238);
   U2484 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n4599, B1 => 
                           REGISTERS_30_15_port, B2 => n4609, ZN => n4237);
   U2485 : NAND4_X1 port map( A1 => n4240, A2 => n4239, A3 => n4238, A4 => 
                           n4237, ZN => n4241);
   U2486 : NOR2_X1 port map( A1 => n4242, A2 => n4241, ZN => n4254);
   U2487 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n4636, B1 => 
                           REGISTERS_3_15_port, B2 => n4623, ZN => n4246);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_1_15_port, A2 => n4621, B1 => 
                           REGISTERS_0_15_port, B2 => n4620, ZN => n4245);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_5_15_port, A2 => n4632, B1 => 
                           REGISTERS_6_15_port, B2 => n4521, ZN => n4244);
   U2490 : AOI22_X1 port map( A1 => REGISTERS_2_15_port, A2 => n4579, B1 => 
                           REGISTERS_7_15_port, B2 => n4635, ZN => n4243);
   U2491 : NAND4_X1 port map( A1 => n4246, A2 => n4245, A3 => n4244, A4 => 
                           n4243, ZN => n4252);
   U2492 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n4620, B1 => 
                           REGISTERS_14_15_port, B2 => n4521, ZN => n4250);
   U2493 : AOI22_X1 port map( A1 => REGISTERS_13_15_port, A2 => n4557, B1 => 
                           REGISTERS_12_15_port, B2 => n4549, ZN => n4249);
   U2494 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n4624, B1 => 
                           REGISTERS_10_15_port, B2 => n4501, ZN => n4248);
   U2495 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n4556, B1 => 
                           REGISTERS_11_15_port, B2 => n4548, ZN => n4247);
   U2496 : NAND4_X1 port map( A1 => n4250, A2 => n4249, A3 => n4248, A4 => 
                           n4247, ZN => n4251);
   U2497 : AOI22_X1 port map( A1 => n4483, A2 => n4252, B1 => n4481, B2 => 
                           n4251, ZN => n4253);
   U2498 : OAI21_X1 port map( B1 => n4593, B2 => n4254, A => n4253, ZN => N400)
                           ;
   U2499 : AOI22_X1 port map( A1 => REGISTERS_22_14_port, A2 => n4510, B1 => 
                           REGISTERS_23_14_port, B2 => n4610, ZN => n4258);
   U2500 : AOI22_X1 port map( A1 => REGISTERS_31_14_port, A2 => n4611, B1 => 
                           REGISTERS_26_14_port, B2 => n4601, ZN => n4257);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_17_14_port, A2 => n4608, B1 => 
                           REGISTERS_21_14_port, B2 => n4570, ZN => n4256);
   U2502 : AOI22_X1 port map( A1 => REGISTERS_19_14_port, A2 => n4599, B1 => 
                           REGISTERS_18_14_port, B2 => n4597, ZN => n4255);
   U2503 : NAND4_X1 port map( A1 => n4258, A2 => n4257, A3 => n4256, A4 => 
                           n4255, ZN => n4264);
   U2504 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n4415, B1 => 
                           REGISTERS_16_14_port, B2 => n4613, ZN => n4262);
   U2505 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n4539, B1 => 
                           REGISTERS_25_14_port, B2 => n4606, ZN => n4261);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n4572, B1 => 
                           REGISTERS_24_14_port, B2 => n4612, ZN => n4260);
   U2507 : AOI22_X1 port map( A1 => REGISTERS_30_14_port, A2 => n4326, B1 => 
                           REGISTERS_27_14_port, B2 => n4349, ZN => n4259);
   U2508 : NAND4_X1 port map( A1 => n4262, A2 => n4261, A3 => n4260, A4 => 
                           n4259, ZN => n4263);
   U2509 : NOR2_X1 port map( A1 => n4264, A2 => n4263, ZN => n4276);
   U2510 : AOI22_X1 port map( A1 => REGISTERS_3_14_port, A2 => n4548, B1 => 
                           REGISTERS_0_14_port, B2 => n4634, ZN => n4268);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n4633, B1 => 
                           REGISTERS_7_14_port, B2 => n4635, ZN => n4267);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_6_14_port, A2 => n4622, B1 => 
                           REGISTERS_4_14_port, B2 => n4549, ZN => n4266);
   U2513 : AOI22_X1 port map( A1 => REGISTERS_2_14_port, A2 => n4631, B1 => 
                           REGISTERS_5_14_port, B2 => n4557, ZN => n4265);
   U2514 : NAND4_X1 port map( A1 => n4268, A2 => n4267, A3 => n4266, A4 => 
                           n4265, ZN => n4274);
   U2515 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n4634, B1 => 
                           REGISTERS_11_14_port, B2 => n4630, ZN => n4272);
   U2516 : AOI22_X1 port map( A1 => REGISTERS_14_14_port, A2 => n4622, B1 => 
                           REGISTERS_12_14_port, B2 => n4549, ZN => n4271);
   U2517 : AOI22_X1 port map( A1 => REGISTERS_10_14_port, A2 => n4631, B1 => 
                           REGISTERS_9_14_port, B2 => n4621, ZN => n4270);
   U2518 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n4632, B1 => 
                           REGISTERS_15_14_port, B2 => n4624, ZN => n4269);
   U2519 : NAND4_X1 port map( A1 => n4272, A2 => n4271, A3 => n4270, A4 => 
                           n4269, ZN => n4273);
   U2520 : AOI22_X1 port map( A1 => n4483, A2 => n4274, B1 => n4481, B2 => 
                           n4273, ZN => n4275);
   U2521 : OAI21_X1 port map( B1 => n4647, B2 => n4276, A => n4275, ZN => N399)
                           ;
   U2522 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n4600, B1 => 
                           REGISTERS_27_13_port, B2 => n4349, ZN => n4280);
   U2523 : AOI22_X1 port map( A1 => REGISTERS_30_13_port, A2 => n4609, B1 => 
                           REGISTERS_22_13_port, B2 => n4510, ZN => n4279);
   U2524 : AOI22_X1 port map( A1 => REGISTERS_31_13_port, A2 => n4611, B1 => 
                           REGISTERS_19_13_port, B2 => n4599, ZN => n4278);
   U2525 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n4612, B1 => 
                           REGISTERS_20_13_port, B2 => n4596, ZN => n4277);
   U2526 : NAND4_X1 port map( A1 => n4280, A2 => n4279, A3 => n4278, A4 => 
                           n4277, ZN => n4286);
   U2527 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n4613, B1 => 
                           REGISTERS_17_13_port, B2 => n4486, ZN => n4284);
   U2528 : AOI22_X1 port map( A1 => REGISTERS_18_13_port, A2 => n4597, B1 => 
                           REGISTERS_28_13_port, B2 => n4595, ZN => n4283);
   U2529 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n4610, B1 => 
                           REGISTERS_29_13_port, B2 => n4572, ZN => n4282);
   U2530 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n4321, B1 => 
                           REGISTERS_26_13_port, B2 => n4601, ZN => n4281);
   U2531 : NAND4_X1 port map( A1 => n4284, A2 => n4283, A3 => n4282, A4 => 
                           n4281, ZN => n4285);
   U2532 : NOR2_X1 port map( A1 => n4286, A2 => n4285, ZN => n4298);
   U2533 : AOI22_X1 port map( A1 => REGISTERS_6_13_port, A2 => n4629, B1 => 
                           REGISTERS_1_13_port, B2 => n4621, ZN => n4290);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n4635, B1 => 
                           REGISTERS_2_13_port, B2 => n4579, ZN => n4289);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_5_13_port, A2 => n4632, B1 => 
                           REGISTERS_4_13_port, B2 => n4549, ZN => n4288);
   U2536 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n4580, B1 => 
                           REGISTERS_3_13_port, B2 => n4623, ZN => n4287);
   U2537 : NAND4_X1 port map( A1 => n4290, A2 => n4289, A3 => n4288, A4 => 
                           n4287, ZN => n4296);
   U2538 : AOI22_X1 port map( A1 => REGISTERS_14_13_port, A2 => n4521, B1 => 
                           REGISTERS_9_13_port, B2 => n4556, ZN => n4294);
   U2539 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n4557, B1 => 
                           REGISTERS_11_13_port, B2 => n4623, ZN => n4293);
   U2540 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n4522, B1 => 
                           REGISTERS_12_13_port, B2 => n4549, ZN => n4292);
   U2541 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n4580, B1 => 
                           REGISTERS_10_13_port, B2 => n4501, ZN => n4291);
   U2542 : NAND4_X1 port map( A1 => n4294, A2 => n4293, A3 => n4292, A4 => 
                           n4291, ZN => n4295);
   U2543 : AOI22_X1 port map( A1 => n4483, A2 => n4296, B1 => n4481, B2 => 
                           n4295, ZN => n4297);
   U2544 : OAI21_X1 port map( B1 => n4593, B2 => n4298, A => n4297, ZN => N398)
                           ;
   U2545 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n4396, B1 => 
                           REGISTERS_20_12_port, B2 => n4596, ZN => n4302);
   U2546 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n4321, B1 => 
                           REGISTERS_17_12_port, B2 => n4608, ZN => n4301);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n4570, B1 => 
                           REGISTERS_30_12_port, B2 => n4609, ZN => n4300);
   U2548 : AOI22_X1 port map( A1 => REGISTERS_31_12_port, A2 => n4571, B1 => 
                           REGISTERS_27_12_port, B2 => n4349, ZN => n4299);
   U2549 : NAND4_X1 port map( A1 => n4302, A2 => n4301, A3 => n4300, A4 => 
                           n4299, ZN => n4308);
   U2550 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n4572, B1 => 
                           REGISTERS_26_12_port, B2 => n4601, ZN => n4306);
   U2551 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n4595, B1 => 
                           REGISTERS_16_12_port, B2 => n4613, ZN => n4305);
   U2552 : AOI22_X1 port map( A1 => REGISTERS_19_12_port, A2 => n4599, B1 => 
                           REGISTERS_23_12_port, B2 => n4610, ZN => n4304);
   U2553 : AOI22_X1 port map( A1 => REGISTERS_22_12_port, A2 => n4510, B1 => 
                           REGISTERS_18_12_port, B2 => n4540, ZN => n4303);
   U2554 : NAND4_X1 port map( A1 => n4306, A2 => n4305, A3 => n4304, A4 => 
                           n4303, ZN => n4307);
   U2555 : NOR2_X1 port map( A1 => n4308, A2 => n4307, ZN => n4320);
   U2556 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n4636, B1 => 
                           REGISTERS_7_12_port, B2 => n4624, ZN => n4312);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_1_12_port, A2 => n4556, B1 => 
                           REGISTERS_3_12_port, B2 => n4630, ZN => n4311);
   U2558 : AOI22_X1 port map( A1 => REGISTERS_5_12_port, A2 => n4632, B1 => 
                           REGISTERS_6_12_port, B2 => n4521, ZN => n4310);
   U2559 : AOI22_X1 port map( A1 => REGISTERS_2_12_port, A2 => n4579, B1 => 
                           REGISTERS_0_12_port, B2 => n4620, ZN => n4309);
   U2560 : NAND4_X1 port map( A1 => n4312, A2 => n4311, A3 => n4310, A4 => 
                           n4309, ZN => n4318);
   U2561 : AOI22_X1 port map( A1 => REGISTERS_9_12_port, A2 => n4556, B1 => 
                           REGISTERS_12_12_port, B2 => n4549, ZN => n4316);
   U2562 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n4634, B1 => 
                           REGISTERS_13_12_port, B2 => n4550, ZN => n4315);
   U2563 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n4548, B1 => 
                           REGISTERS_15_12_port, B2 => n4522, ZN => n4314);
   U2564 : AOI22_X1 port map( A1 => REGISTERS_14_12_port, A2 => n4521, B1 => 
                           REGISTERS_10_12_port, B2 => n4631, ZN => n4313);
   U2565 : NAND4_X1 port map( A1 => n4316, A2 => n4315, A3 => n4314, A4 => 
                           n4313, ZN => n4317);
   U2566 : AOI22_X1 port map( A1 => n4483, A2 => n4318, B1 => n4481, B2 => 
                           n4317, ZN => n4319);
   U2567 : OAI21_X1 port map( B1 => n4647, B2 => n4320, A => n4319, ZN => N397)
                           ;
   U2568 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n4599, B1 => 
                           REGISTERS_17_11_port, B2 => n4608, ZN => n4325);
   U2569 : AOI22_X1 port map( A1 => REGISTERS_25_11_port, A2 => n4321, B1 => 
                           REGISTERS_29_11_port, B2 => n4572, ZN => n4324);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_22_11_port, A2 => n4510, B1 => 
                           REGISTERS_31_11_port, B2 => n4611, ZN => n4323);
   U2571 : AOI22_X1 port map( A1 => REGISTERS_26_11_port, A2 => n4601, B1 => 
                           REGISTERS_20_11_port, B2 => n4596, ZN => n4322);
   U2572 : NAND4_X1 port map( A1 => n4325, A2 => n4324, A3 => n4323, A4 => 
                           n4322, ZN => n4332);
   U2573 : AOI22_X1 port map( A1 => REGISTERS_30_11_port, A2 => n4326, B1 => 
                           REGISTERS_28_11_port, B2 => n4539, ZN => n4330);
   U2574 : AOI22_X1 port map( A1 => REGISTERS_18_11_port, A2 => n4597, B1 => 
                           REGISTERS_24_11_port, B2 => n4612, ZN => n4329);
   U2575 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n4613, B1 => 
                           REGISTERS_23_11_port, B2 => n4610, ZN => n4328);
   U2576 : AOI22_X1 port map( A1 => REGISTERS_21_11_port, A2 => n4570, B1 => 
                           REGISTERS_27_11_port, B2 => n4607, ZN => n4327);
   U2577 : NAND4_X1 port map( A1 => n4330, A2 => n4329, A3 => n4328, A4 => 
                           n4327, ZN => n4331);
   U2578 : NOR2_X1 port map( A1 => n4332, A2 => n4331, ZN => n4344);
   U2579 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n4634, B1 => 
                           REGISTERS_2_11_port, B2 => n4579, ZN => n4336);
   U2580 : AOI22_X1 port map( A1 => REGISTERS_3_11_port, A2 => n4548, B1 => 
                           REGISTERS_7_11_port, B2 => n4522, ZN => n4335);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n4556, B1 => 
                           REGISTERS_4_11_port, B2 => n4549, ZN => n4334);
   U2582 : AOI22_X1 port map( A1 => REGISTERS_6_11_port, A2 => n4622, B1 => 
                           REGISTERS_5_11_port, B2 => n4557, ZN => n4333);
   U2583 : NAND4_X1 port map( A1 => n4336, A2 => n4335, A3 => n4334, A4 => 
                           n4333, ZN => n4342);
   U2584 : AOI22_X1 port map( A1 => REGISTERS_15_11_port, A2 => n4624, B1 => 
                           REGISTERS_12_11_port, B2 => n4549, ZN => n4340);
   U2585 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n4632, B1 => 
                           REGISTERS_11_11_port, B2 => n4623, ZN => n4339);
   U2586 : AOI22_X1 port map( A1 => REGISTERS_14_11_port, A2 => n4629, B1 => 
                           REGISTERS_9_11_port, B2 => n4633, ZN => n4338);
   U2587 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n4579, B1 => 
                           REGISTERS_8_11_port, B2 => n4634, ZN => n4337);
   U2588 : NAND4_X1 port map( A1 => n4340, A2 => n4339, A3 => n4338, A4 => 
                           n4337, ZN => n4341);
   U2589 : AOI22_X1 port map( A1 => n4483, A2 => n4342, B1 => n4481, B2 => 
                           n4341, ZN => n4343);
   U2590 : OAI21_X1 port map( B1 => n4647, B2 => n4344, A => n4343, ZN => N396)
                           ;
   U2591 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n4608, B1 => 
                           REGISTERS_22_10_port, B2 => n4510, ZN => n4348);
   U2592 : AOI22_X1 port map( A1 => REGISTERS_26_10_port, A2 => n4601, B1 => 
                           REGISTERS_25_10_port, B2 => n4606, ZN => n4347);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_31_10_port, A2 => n4611, B1 => 
                           REGISTERS_23_10_port, B2 => n4610, ZN => n4346);
   U2594 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n4396, B1 => 
                           REGISTERS_30_10_port, B2 => n4609, ZN => n4345);
   U2595 : NAND4_X1 port map( A1 => n4348, A2 => n4347, A3 => n4346, A4 => 
                           n4345, ZN => n4355);
   U2596 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n4599, B1 => 
                           REGISTERS_21_10_port, B2 => n4570, ZN => n4353);
   U2597 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n4595, B1 => 
                           REGISTERS_18_10_port, B2 => n4540, ZN => n4352);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n4572, B1 => 
                           REGISTERS_16_10_port, B2 => n4613, ZN => n4351);
   U2599 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n4349, B1 => 
                           REGISTERS_20_10_port, B2 => n4596, ZN => n4350);
   U2600 : NAND4_X1 port map( A1 => n4353, A2 => n4352, A3 => n4351, A4 => 
                           n4350, ZN => n4354);
   U2601 : NOR2_X1 port map( A1 => n4355, A2 => n4354, ZN => n4367);
   U2602 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n4557, B1 => 
                           REGISTERS_1_10_port, B2 => n4621, ZN => n4359);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_6_10_port, A2 => n4521, B1 => 
                           REGISTERS_7_10_port, B2 => n4522, ZN => n4358);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_2_10_port, A2 => n4579, B1 => 
                           REGISTERS_0_10_port, B2 => n4634, ZN => n4357);
   U2605 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n4636, B1 => 
                           REGISTERS_3_10_port, B2 => n4630, ZN => n4356);
   U2606 : NAND4_X1 port map( A1 => n4359, A2 => n4358, A3 => n4357, A4 => 
                           n4356, ZN => n4365);
   U2607 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n4556, B1 => 
                           REGISTERS_11_10_port, B2 => n4623, ZN => n4363);
   U2608 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n4555, B1 => 
                           REGISTERS_8_10_port, B2 => n4580, ZN => n4362);
   U2609 : AOI22_X1 port map( A1 => REGISTERS_14_10_port, A2 => n4629, B1 => 
                           REGISTERS_13_10_port, B2 => n4632, ZN => n4361);
   U2610 : AOI22_X1 port map( A1 => REGISTERS_10_10_port, A2 => n4631, B1 => 
                           REGISTERS_15_10_port, B2 => n4635, ZN => n4360);
   U2611 : NAND4_X1 port map( A1 => n4363, A2 => n4362, A3 => n4361, A4 => 
                           n4360, ZN => n4364);
   U2612 : AOI22_X1 port map( A1 => n4483, A2 => n4365, B1 => n4481, B2 => 
                           n4364, ZN => n4366);
   U2613 : OAI21_X1 port map( B1 => n4647, B2 => n4367, A => n4366, ZN => N395)
                           ;
   U2614 : AOI22_X1 port map( A1 => REGISTERS_18_9_port, A2 => n4597, B1 => 
                           REGISTERS_24_9_port, B2 => n4612, ZN => n4371);
   U2615 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n4610, B1 => 
                           REGISTERS_29_9_port, B2 => n4598, ZN => n4370);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n4570, B1 => 
                           REGISTERS_30_9_port, B2 => n4609, ZN => n4369);
   U2617 : AOI22_X1 port map( A1 => REGISTERS_31_9_port, A2 => n4611, B1 => 
                           REGISTERS_20_9_port, B2 => n4596, ZN => n4368);
   U2618 : NAND4_X1 port map( A1 => n4371, A2 => n4370, A3 => n4369, A4 => 
                           n4368, ZN => n4377);
   U2619 : AOI22_X1 port map( A1 => REGISTERS_22_9_port, A2 => n4510, B1 => 
                           REGISTERS_27_9_port, B2 => n4607, ZN => n4375);
   U2620 : AOI22_X1 port map( A1 => REGISTERS_26_9_port, A2 => n4601, B1 => 
                           REGISTERS_19_9_port, B2 => n4599, ZN => n4374);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n4595, B1 => 
                           REGISTERS_17_9_port, B2 => n4608, ZN => n4373);
   U2622 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n4613, B1 => 
                           REGISTERS_25_9_port, B2 => n4606, ZN => n4372);
   U2623 : NAND4_X1 port map( A1 => n4375, A2 => n4374, A3 => n4373, A4 => 
                           n4372, ZN => n4376);
   U2624 : NOR2_X1 port map( A1 => n4377, A2 => n4376, ZN => n4389);
   U2625 : AOI22_X1 port map( A1 => REGISTERS_6_9_port, A2 => n4629, B1 => 
                           REGISTERS_4_9_port, B2 => n4549, ZN => n4381);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n4635, B1 => 
                           REGISTERS_0_9_port, B2 => n4634, ZN => n4380);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n4556, B1 => 
                           REGISTERS_5_9_port, B2 => n4550, ZN => n4379);
   U2628 : AOI22_X1 port map( A1 => REGISTERS_2_9_port, A2 => n4501, B1 => 
                           REGISTERS_3_9_port, B2 => n4630, ZN => n4378);
   U2629 : NAND4_X1 port map( A1 => n4381, A2 => n4380, A3 => n4379, A4 => 
                           n4378, ZN => n4387);
   U2630 : AOI22_X1 port map( A1 => REGISTERS_13_9_port, A2 => n4550, B1 => 
                           REGISTERS_11_9_port, B2 => n4630, ZN => n4385);
   U2631 : AOI22_X1 port map( A1 => REGISTERS_10_9_port, A2 => n4579, B1 => 
                           REGISTERS_12_9_port, B2 => n4549, ZN => n4384);
   U2632 : AOI22_X1 port map( A1 => REGISTERS_9_9_port, A2 => n4556, B1 => 
                           REGISTERS_14_9_port, B2 => n4629, ZN => n4383);
   U2633 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n4522, B1 => 
                           REGISTERS_8_9_port, B2 => n4634, ZN => n4382);
   U2634 : NAND4_X1 port map( A1 => n4385, A2 => n4384, A3 => n4383, A4 => 
                           n4382, ZN => n4386);
   U2635 : AOI22_X1 port map( A1 => n4483, A2 => n4387, B1 => n4481, B2 => 
                           n4386, ZN => n4388);
   U2636 : OAI21_X1 port map( B1 => n4593, B2 => n4389, A => n4388, ZN => N394)
                           ;
   U2637 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n4595, B1 => 
                           REGISTERS_30_8_port, B2 => n4609, ZN => n4394);
   U2638 : AOI22_X1 port map( A1 => REGISTERS_21_8_port, A2 => n4570, B1 => 
                           REGISTERS_17_8_port, B2 => n4608, ZN => n4393);
   U2639 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n4607, B1 => 
                           REGISTERS_22_8_port, B2 => n4594, ZN => n4392);
   U2640 : AOI22_X1 port map( A1 => REGISTERS_26_8_port, A2 => n4390, B1 => 
                           REGISTERS_18_8_port, B2 => n4540, ZN => n4391);
   U2641 : NAND4_X1 port map( A1 => n4394, A2 => n4393, A3 => n4392, A4 => 
                           n4391, ZN => n4402);
   U2642 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n4395, B1 => 
                           REGISTERS_29_8_port, B2 => n4598, ZN => n4400);
   U2643 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n4396, B1 => 
                           REGISTERS_19_8_port, B2 => n4541, ZN => n4399);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n4610, B1 => 
                           REGISTERS_25_8_port, B2 => n4606, ZN => n4398);
   U2645 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n4596, B1 => 
                           REGISTERS_31_8_port, B2 => n4571, ZN => n4397);
   U2646 : NAND4_X1 port map( A1 => n4400, A2 => n4399, A3 => n4398, A4 => 
                           n4397, ZN => n4401);
   U2647 : NOR2_X1 port map( A1 => n4402, A2 => n4401, ZN => n4414);
   U2648 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n4634, B1 => 
                           REGISTERS_4_8_port, B2 => n4549, ZN => n4406);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_5_8_port, A2 => n4557, B1 => 
                           REGISTERS_1_8_port, B2 => n4633, ZN => n4405);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n4624, B1 => 
                           REGISTERS_2_8_port, B2 => n4501, ZN => n4404);
   U2651 : AOI22_X1 port map( A1 => REGISTERS_6_8_port, A2 => n4521, B1 => 
                           REGISTERS_3_8_port, B2 => n4623, ZN => n4403);
   U2652 : NAND4_X1 port map( A1 => n4406, A2 => n4405, A3 => n4404, A4 => 
                           n4403, ZN => n4412);
   U2653 : AOI22_X1 port map( A1 => REGISTERS_13_8_port, A2 => n4557, B1 => 
                           REGISTERS_10_8_port, B2 => n4501, ZN => n4410);
   U2654 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n4624, B1 => 
                           REGISTERS_8_8_port, B2 => n4620, ZN => n4409);
   U2655 : AOI22_X1 port map( A1 => REGISTERS_14_8_port, A2 => n4629, B1 => 
                           REGISTERS_11_8_port, B2 => n4630, ZN => n4408);
   U2656 : AOI22_X1 port map( A1 => REGISTERS_9_8_port, A2 => n4633, B1 => 
                           REGISTERS_12_8_port, B2 => n4636, ZN => n4407);
   U2657 : NAND4_X1 port map( A1 => n4410, A2 => n4409, A3 => n4408, A4 => 
                           n4407, ZN => n4411);
   U2658 : AOI22_X1 port map( A1 => n4483, A2 => n4412, B1 => n4481, B2 => 
                           n4411, ZN => n4413);
   U2659 : OAI21_X1 port map( B1 => n4647, B2 => n4414, A => n4413, ZN => N393)
                           ;
   U2660 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n4570, B1 => 
                           REGISTERS_27_7_port, B2 => n4607, ZN => n4419);
   U2661 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n4415, B1 => 
                           REGISTERS_25_7_port, B2 => n4606, ZN => n4418);
   U2662 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n4613, B1 => 
                           REGISTERS_30_7_port, B2 => n4609, ZN => n4417);
   U2663 : AOI22_X1 port map( A1 => REGISTERS_26_7_port, A2 => n4601, B1 => 
                           REGISTERS_18_7_port, B2 => n4540, ZN => n4416);
   U2664 : NAND4_X1 port map( A1 => n4419, A2 => n4418, A3 => n4417, A4 => 
                           n4416, ZN => n4426);
   U2665 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n4595, B1 => 
                           REGISTERS_24_7_port, B2 => n4612, ZN => n4424);
   U2666 : AOI22_X1 port map( A1 => REGISTERS_17_7_port, A2 => n4486, B1 => 
                           REGISTERS_31_7_port, B2 => n4571, ZN => n4423);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_23_7_port, A2 => n4420, B1 => 
                           REGISTERS_19_7_port, B2 => n4541, ZN => n4422);
   U2668 : AOI22_X1 port map( A1 => REGISTERS_22_7_port, A2 => n4510, B1 => 
                           REGISTERS_29_7_port, B2 => n4598, ZN => n4421);
   U2669 : NAND4_X1 port map( A1 => n4424, A2 => n4423, A3 => n4422, A4 => 
                           n4421, ZN => n4425);
   U2670 : NOR2_X1 port map( A1 => n4426, A2 => n4425, ZN => n4438);
   U2671 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n4548, B1 => 
                           REGISTERS_7_7_port, B2 => n4522, ZN => n4430);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_5_7_port, A2 => n4632, B1 => 
                           REGISTERS_4_7_port, B2 => n4636, ZN => n4429);
   U2673 : AOI22_X1 port map( A1 => REGISTERS_2_7_port, A2 => n4631, B1 => 
                           REGISTERS_1_7_port, B2 => n4621, ZN => n4428);
   U2674 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n4580, B1 => 
                           REGISTERS_6_7_port, B2 => n4629, ZN => n4427);
   U2675 : NAND4_X1 port map( A1 => n4430, A2 => n4429, A3 => n4428, A4 => 
                           n4427, ZN => n4436);
   U2676 : AOI22_X1 port map( A1 => REGISTERS_9_7_port, A2 => n4556, B1 => 
                           REGISTERS_14_7_port, B2 => n4629, ZN => n4434);
   U2677 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n4548, B1 => 
                           REGISTERS_15_7_port, B2 => n4522, ZN => n4433);
   U2678 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n4549, B1 => 
                           REGISTERS_13_7_port, B2 => n4550, ZN => n4432);
   U2679 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n4634, B1 => 
                           REGISTERS_10_7_port, B2 => n4579, ZN => n4431);
   U2680 : NAND4_X1 port map( A1 => n4434, A2 => n4433, A3 => n4432, A4 => 
                           n4431, ZN => n4435);
   U2681 : AOI22_X1 port map( A1 => n4483, A2 => n4436, B1 => n4481, B2 => 
                           n4435, ZN => n4437);
   U2682 : OAI21_X1 port map( B1 => n4593, B2 => n4438, A => n4437, ZN => N392)
                           ;
   U2683 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n4572, B1 => 
                           REGISTERS_21_6_port, B2 => n4600, ZN => n4442);
   U2684 : AOI22_X1 port map( A1 => REGISTERS_18_6_port, A2 => n4597, B1 => 
                           REGISTERS_19_6_port, B2 => n4541, ZN => n4441);
   U2685 : AOI22_X1 port map( A1 => REGISTERS_17_6_port, A2 => n4608, B1 => 
                           REGISTERS_28_6_port, B2 => n4539, ZN => n4440);
   U2686 : AOI22_X1 port map( A1 => REGISTERS_22_6_port, A2 => n4510, B1 => 
                           REGISTERS_20_6_port, B2 => n4596, ZN => n4439);
   U2687 : NAND4_X1 port map( A1 => n4442, A2 => n4441, A3 => n4440, A4 => 
                           n4439, ZN => n4448);
   U2688 : AOI22_X1 port map( A1 => REGISTERS_26_6_port, A2 => n4601, B1 => 
                           REGISTERS_16_6_port, B2 => n4613, ZN => n4446);
   U2689 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n4606, B1 => 
                           REGISTERS_23_6_port, B2 => n4610, ZN => n4445);
   U2690 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n4612, B1 => 
                           REGISTERS_30_6_port, B2 => n4609, ZN => n4444);
   U2691 : AOI22_X1 port map( A1 => REGISTERS_31_6_port, A2 => n4611, B1 => 
                           REGISTERS_27_6_port, B2 => n4607, ZN => n4443);
   U2692 : NAND4_X1 port map( A1 => n4446, A2 => n4445, A3 => n4444, A4 => 
                           n4443, ZN => n4447);
   U2693 : NOR2_X1 port map( A1 => n4448, A2 => n4447, ZN => n4461);
   U2694 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n4620, B1 => 
                           REGISTERS_3_6_port, B2 => n4630, ZN => n4452);
   U2695 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n4557, B1 => 
                           REGISTERS_7_6_port, B2 => n4635, ZN => n4451);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_6_6_port, A2 => n4629, B1 => 
                           REGISTERS_1_6_port, B2 => n4621, ZN => n4450);
   U2697 : AOI22_X1 port map( A1 => REGISTERS_2_6_port, A2 => n4631, B1 => 
                           REGISTERS_4_6_port, B2 => n4636, ZN => n4449);
   U2698 : NAND4_X1 port map( A1 => n4452, A2 => n4451, A3 => n4450, A4 => 
                           n4449, ZN => n4458);
   U2699 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n4624, B1 => 
                           REGISTERS_12_6_port, B2 => n4549, ZN => n4456);
   U2700 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n4548, B1 => 
                           REGISTERS_14_6_port, B2 => n4629, ZN => n4455);
   U2701 : AOI22_X1 port map( A1 => REGISTERS_9_6_port, A2 => n4556, B1 => 
                           REGISTERS_10_6_port, B2 => n4631, ZN => n4454);
   U2702 : AOI22_X1 port map( A1 => REGISTERS_13_6_port, A2 => n4550, B1 => 
                           REGISTERS_8_6_port, B2 => n4620, ZN => n4453);
   U2703 : NAND4_X1 port map( A1 => n4456, A2 => n4455, A3 => n4454, A4 => 
                           n4453, ZN => n4457);
   U2704 : AOI22_X1 port map( A1 => n4459, A2 => n4458, B1 => n4481, B2 => 
                           n4457, ZN => n4460);
   U2705 : OAI21_X1 port map( B1 => n4647, B2 => n4461, A => n4460, ZN => N391)
                           ;
   U2706 : AOI22_X1 port map( A1 => REGISTERS_30_5_port, A2 => n4609, B1 => 
                           REGISTERS_22_5_port, B2 => n4594, ZN => n4465);
   U2707 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n4610, B1 => 
                           REGISTERS_26_5_port, B2 => n4601, ZN => n4464);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_21_5_port, A2 => n4570, B1 => 
                           REGISTERS_19_5_port, B2 => n4541, ZN => n4463);
   U2709 : AOI22_X1 port map( A1 => REGISTERS_18_5_port, A2 => n4597, B1 => 
                           REGISTERS_28_5_port, B2 => n4539, ZN => n4462);
   U2710 : NAND4_X1 port map( A1 => n4465, A2 => n4464, A3 => n4463, A4 => 
                           n4462, ZN => n4471);
   U2711 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n4596, B1 => 
                           REGISTERS_24_5_port, B2 => n4612, ZN => n4469);
   U2712 : AOI22_X1 port map( A1 => REGISTERS_25_5_port, A2 => n4606, B1 => 
                           REGISTERS_29_5_port, B2 => n4598, ZN => n4468);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_31_5_port, A2 => n4611, B1 => 
                           REGISTERS_16_5_port, B2 => n4613, ZN => n4467);
   U2714 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n4607, B1 => 
                           REGISTERS_17_5_port, B2 => n4608, ZN => n4466);
   U2715 : NAND4_X1 port map( A1 => n4469, A2 => n4468, A3 => n4467, A4 => 
                           n4466, ZN => n4470);
   U2716 : NOR2_X1 port map( A1 => n4471, A2 => n4470, ZN => n4485);
   U2717 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n4556, B1 => 
                           REGISTERS_4_5_port, B2 => n4636, ZN => n4475);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_3_5_port, A2 => n4548, B1 => 
                           REGISTERS_0_5_port, B2 => n4634, ZN => n4474);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n4624, B1 => 
                           REGISTERS_5_5_port, B2 => n4550, ZN => n4473);
   U2720 : AOI22_X1 port map( A1 => REGISTERS_2_5_port, A2 => n4631, B1 => 
                           REGISTERS_6_5_port, B2 => n4629, ZN => n4472);
   U2721 : NAND4_X1 port map( A1 => n4475, A2 => n4474, A3 => n4473, A4 => 
                           n4472, ZN => n4482);
   U2722 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n4636, B1 => 
                           REGISTERS_9_5_port, B2 => n4633, ZN => n4479);
   U2723 : AOI22_X1 port map( A1 => REGISTERS_13_5_port, A2 => n4550, B1 => 
                           REGISTERS_10_5_port, B2 => n4631, ZN => n4478);
   U2724 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n4580, B1 => 
                           REGISTERS_14_5_port, B2 => n4629, ZN => n4477);
   U2725 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n4624, B1 => 
                           REGISTERS_11_5_port, B2 => n4630, ZN => n4476);
   U2726 : NAND4_X1 port map( A1 => n4479, A2 => n4478, A3 => n4477, A4 => 
                           n4476, ZN => n4480);
   U2727 : AOI22_X1 port map( A1 => n4483, A2 => n4482, B1 => n4481, B2 => 
                           n4480, ZN => n4484);
   U2728 : OAI21_X1 port map( B1 => n4593, B2 => n4485, A => n4484, ZN => N390)
                           ;
   U2729 : AOI22_X1 port map( A1 => REGISTERS_31_4_port, A2 => n4611, B1 => 
                           REGISTERS_27_4_port, B2 => n4607, ZN => n4490);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_26_4_port, A2 => n4601, B1 => 
                           REGISTERS_18_4_port, B2 => n4540, ZN => n4489);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n4570, B1 => 
                           REGISTERS_29_4_port, B2 => n4598, ZN => n4488);
   U2732 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n4486, B1 => 
                           REGISTERS_25_4_port, B2 => n4606, ZN => n4487);
   U2733 : NAND4_X1 port map( A1 => n4490, A2 => n4489, A3 => n4488, A4 => 
                           n4487, ZN => n4496);
   U2734 : AOI22_X1 port map( A1 => REGISTERS_30_4_port, A2 => n4609, B1 => 
                           REGISTERS_24_4_port, B2 => n4612, ZN => n4494);
   U2735 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n4613, B1 => 
                           REGISTERS_23_4_port, B2 => n4610, ZN => n4493);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_22_4_port, A2 => n4510, B1 => 
                           REGISTERS_20_4_port, B2 => n4596, ZN => n4492);
   U2737 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n4595, B1 => 
                           REGISTERS_19_4_port, B2 => n4541, ZN => n4491);
   U2738 : NAND4_X1 port map( A1 => n4494, A2 => n4493, A3 => n4492, A4 => 
                           n4491, ZN => n4495);
   U2739 : NOR2_X1 port map( A1 => n4496, A2 => n4495, ZN => n4509);
   U2740 : AOI22_X1 port map( A1 => REGISTERS_2_4_port, A2 => n4631, B1 => 
                           REGISTERS_0_4_port, B2 => n4580, ZN => n4500);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n4624, B1 => 
                           REGISTERS_5_4_port, B2 => n4632, ZN => n4499);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n4555, B1 => 
                           REGISTERS_1_4_port, B2 => n4621, ZN => n4498);
   U2743 : AOI22_X1 port map( A1 => REGISTERS_6_4_port, A2 => n4629, B1 => 
                           REGISTERS_3_4_port, B2 => n4623, ZN => n4497);
   U2744 : NAND4_X1 port map( A1 => n4500, A2 => n4499, A3 => n4498, A4 => 
                           n4497, ZN => n4507);
   U2745 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n4556, B1 => 
                           REGISTERS_10_4_port, B2 => n4501, ZN => n4505);
   U2746 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n4624, B1 => 
                           REGISTERS_14_4_port, B2 => n4629, ZN => n4504);
   U2747 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n4555, B1 => 
                           REGISTERS_8_4_port, B2 => n4580, ZN => n4503);
   U2748 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n4548, B1 => 
                           REGISTERS_13_4_port, B2 => n4557, ZN => n4502);
   U2749 : NAND4_X1 port map( A1 => n4505, A2 => n4504, A3 => n4503, A4 => 
                           n4502, ZN => n4506);
   U2750 : AOI22_X1 port map( A1 => n4644, A2 => n4507, B1 => n4642, B2 => 
                           n4506, ZN => n4508);
   U2751 : OAI21_X1 port map( B1 => n4647, B2 => n4509, A => n4508, ZN => N389)
                           ;
   U2752 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n4612, B1 => 
                           REGISTERS_19_3_port, B2 => n4541, ZN => n4514);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_26_3_port, A2 => n4601, B1 => 
                           REGISTERS_17_3_port, B2 => n4608, ZN => n4513);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_22_3_port, A2 => n4510, B1 => 
                           REGISTERS_27_3_port, B2 => n4607, ZN => n4512);
   U2755 : AOI22_X1 port map( A1 => REGISTERS_23_3_port, A2 => n4610, B1 => 
                           REGISTERS_31_3_port, B2 => n4571, ZN => n4511);
   U2756 : NAND4_X1 port map( A1 => n4514, A2 => n4513, A3 => n4512, A4 => 
                           n4511, ZN => n4520);
   U2757 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n4595, B1 => 
                           REGISTERS_16_3_port, B2 => n4613, ZN => n4518);
   U2758 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n4572, B1 => 
                           REGISTERS_25_3_port, B2 => n4606, ZN => n4517);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_18_3_port, A2 => n4597, B1 => 
                           REGISTERS_30_3_port, B2 => n4609, ZN => n4516);
   U2760 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n4596, B1 => 
                           REGISTERS_21_3_port, B2 => n4600, ZN => n4515);
   U2761 : NAND4_X1 port map( A1 => n4518, A2 => n4517, A3 => n4516, A4 => 
                           n4515, ZN => n4519);
   U2762 : NOR2_X1 port map( A1 => n4520, A2 => n4519, ZN => n4534);
   U2763 : AOI22_X1 port map( A1 => REGISTERS_2_3_port, A2 => n4631, B1 => 
                           REGISTERS_6_3_port, B2 => n4521, ZN => n4526);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n4636, B1 => 
                           REGISTERS_1_3_port, B2 => n4621, ZN => n4525);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_3_3_port, A2 => n4548, B1 => 
                           REGISTERS_5_3_port, B2 => n4632, ZN => n4524);
   U2766 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n4580, B1 => 
                           REGISTERS_7_3_port, B2 => n4522, ZN => n4523);
   U2767 : NAND4_X1 port map( A1 => n4526, A2 => n4525, A3 => n4524, A4 => 
                           n4523, ZN => n4532);
   U2768 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n4632, B1 => 
                           REGISTERS_14_3_port, B2 => n4622, ZN => n4530);
   U2769 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n4548, B1 => 
                           REGISTERS_9_3_port, B2 => n4633, ZN => n4529);
   U2770 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n4580, B1 => 
                           REGISTERS_15_3_port, B2 => n4635, ZN => n4528);
   U2771 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n4555, B1 => 
                           REGISTERS_10_3_port, B2 => n4579, ZN => n4527);
   U2772 : NAND4_X1 port map( A1 => n4530, A2 => n4529, A3 => n4528, A4 => 
                           n4527, ZN => n4531);
   U2773 : AOI22_X1 port map( A1 => n4644, A2 => n4532, B1 => n4642, B2 => 
                           n4531, ZN => n4533);
   U2774 : OAI21_X1 port map( B1 => n4593, B2 => n4534, A => n4533, ZN => N388)
                           ;
   U2775 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n4610, B1 => 
                           REGISTERS_30_2_port, B2 => n4609, ZN => n4538);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n4607, B1 => 
                           REGISTERS_20_2_port, B2 => n4596, ZN => n4537);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n4570, B1 => 
                           REGISTERS_22_2_port, B2 => n4594, ZN => n4536);
   U2778 : AOI22_X1 port map( A1 => REGISTERS_26_2_port, A2 => n4601, B1 => 
                           REGISTERS_29_2_port, B2 => n4598, ZN => n4535);
   U2779 : NAND4_X1 port map( A1 => n4538, A2 => n4537, A3 => n4536, A4 => 
                           n4535, ZN => n4547);
   U2780 : AOI22_X1 port map( A1 => REGISTERS_31_2_port, A2 => n4611, B1 => 
                           REGISTERS_28_2_port, B2 => n4539, ZN => n4545);
   U2781 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n4613, B1 => 
                           REGISTERS_18_2_port, B2 => n4540, ZN => n4544);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_25_2_port, A2 => n4606, B1 => 
                           REGISTERS_24_2_port, B2 => n4612, ZN => n4543);
   U2783 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n4608, B1 => 
                           REGISTERS_19_2_port, B2 => n4541, ZN => n4542);
   U2784 : NAND4_X1 port map( A1 => n4545, A2 => n4544, A3 => n4543, A4 => 
                           n4542, ZN => n4546);
   U2785 : NOR2_X1 port map( A1 => n4547, A2 => n4546, ZN => n4565);
   U2786 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n4624, B1 => 
                           REGISTERS_0_2_port, B2 => n4580, ZN => n4554);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n4548, B1 => 
                           REGISTERS_6_2_port, B2 => n4622, ZN => n4553);
   U2788 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n4549, B1 => 
                           REGISTERS_1_2_port, B2 => n4621, ZN => n4552);
   U2789 : AOI22_X1 port map( A1 => REGISTERS_2_2_port, A2 => n4631, B1 => 
                           REGISTERS_5_2_port, B2 => n4550, ZN => n4551);
   U2790 : NAND4_X1 port map( A1 => n4554, A2 => n4553, A3 => n4552, A4 => 
                           n4551, ZN => n4563);
   U2791 : AOI22_X1 port map( A1 => REGISTERS_9_2_port, A2 => n4556, B1 => 
                           REGISTERS_12_2_port, B2 => n4555, ZN => n4561);
   U2792 : AOI22_X1 port map( A1 => REGISTERS_14_2_port, A2 => n4622, B1 => 
                           REGISTERS_11_2_port, B2 => n4623, ZN => n4560);
   U2793 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n4624, B1 => 
                           REGISTERS_8_2_port, B2 => n4620, ZN => n4559);
   U2794 : AOI22_X1 port map( A1 => REGISTERS_10_2_port, A2 => n4631, B1 => 
                           REGISTERS_13_2_port, B2 => n4557, ZN => n4558);
   U2795 : NAND4_X1 port map( A1 => n4561, A2 => n4560, A3 => n4559, A4 => 
                           n4558, ZN => n4562);
   U2796 : AOI22_X1 port map( A1 => n4644, A2 => n4563, B1 => n4642, B2 => 
                           n4562, ZN => n4564);
   U2797 : OAI21_X1 port map( B1 => n4647, B2 => n4565, A => n4564, ZN => N387)
                           ;
   U2798 : AOI22_X1 port map( A1 => REGISTERS_18_1_port, A2 => n4597, B1 => 
                           REGISTERS_17_1_port, B2 => n4608, ZN => n4569);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n4606, B1 => 
                           REGISTERS_20_1_port, B2 => n4596, ZN => n4568);
   U2800 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n4599, B1 => 
                           REGISTERS_27_1_port, B2 => n4607, ZN => n4567);
   U2801 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n4595, B1 => 
                           REGISTERS_16_1_port, B2 => n4613, ZN => n4566);
   U2802 : NAND4_X1 port map( A1 => n4569, A2 => n4568, A3 => n4567, A4 => 
                           n4566, ZN => n4578);
   U2803 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n4570, B1 => 
                           REGISTERS_24_1_port, B2 => n4612, ZN => n4576);
   U2804 : AOI22_X1 port map( A1 => REGISTERS_30_1_port, A2 => n4609, B1 => 
                           REGISTERS_22_1_port, B2 => n4594, ZN => n4575);
   U2805 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n4572, B1 => 
                           REGISTERS_31_1_port, B2 => n4571, ZN => n4574);
   U2806 : AOI22_X1 port map( A1 => REGISTERS_26_1_port, A2 => n4601, B1 => 
                           REGISTERS_23_1_port, B2 => n4610, ZN => n4573);
   U2807 : NAND4_X1 port map( A1 => n4576, A2 => n4575, A3 => n4574, A4 => 
                           n4573, ZN => n4577);
   U2808 : NOR2_X1 port map( A1 => n4578, A2 => n4577, ZN => n4592);
   U2809 : AOI22_X1 port map( A1 => REGISTERS_5_1_port, A2 => n4632, B1 => 
                           REGISTERS_2_1_port, B2 => n4579, ZN => n4584);
   U2810 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n4624, B1 => 
                           REGISTERS_4_1_port, B2 => n4636, ZN => n4583);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n4580, B1 => 
                           REGISTERS_3_1_port, B2 => n4623, ZN => n4582);
   U2812 : AOI22_X1 port map( A1 => REGISTERS_6_1_port, A2 => n4622, B1 => 
                           REGISTERS_1_1_port, B2 => n4621, ZN => n4581);
   U2813 : NAND4_X1 port map( A1 => n4584, A2 => n4583, A3 => n4582, A4 => 
                           n4581, ZN => n4590);
   U2814 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n4636, B1 => 
                           REGISTERS_8_1_port, B2 => n4620, ZN => n4588);
   U2815 : AOI22_X1 port map( A1 => REGISTERS_15_1_port, A2 => n4624, B1 => 
                           REGISTERS_14_1_port, B2 => n4629, ZN => n4587);
   U2816 : AOI22_X1 port map( A1 => REGISTERS_10_1_port, A2 => n4631, B1 => 
                           REGISTERS_11_1_port, B2 => n4623, ZN => n4586);
   U2817 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n4632, B1 => 
                           REGISTERS_9_1_port, B2 => n4621, ZN => n4585);
   U2818 : NAND4_X1 port map( A1 => n4588, A2 => n4587, A3 => n4586, A4 => 
                           n4585, ZN => n4589);
   U2819 : AOI22_X1 port map( A1 => n4644, A2 => n4590, B1 => n4642, B2 => 
                           n4589, ZN => n4591);
   U2820 : OAI21_X1 port map( B1 => n4593, B2 => n4592, A => n4591, ZN => N386)
                           ;
   U2821 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n4595, B1 => 
                           REGISTERS_22_0_port, B2 => n4594, ZN => n4605);
   U2822 : AOI22_X1 port map( A1 => REGISTERS_18_0_port, A2 => n4597, B1 => 
                           REGISTERS_20_0_port, B2 => n4596, ZN => n4604);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_19_0_port, A2 => n4599, B1 => 
                           REGISTERS_29_0_port, B2 => n4598, ZN => n4603);
   U2824 : AOI22_X1 port map( A1 => REGISTERS_26_0_port, A2 => n4601, B1 => 
                           REGISTERS_21_0_port, B2 => n4600, ZN => n4602);
   U2825 : NAND4_X1 port map( A1 => n4605, A2 => n4604, A3 => n4603, A4 => 
                           n4602, ZN => n4619);
   U2826 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n4607, B1 => 
                           REGISTERS_25_0_port, B2 => n4606, ZN => n4617);
   U2827 : AOI22_X1 port map( A1 => REGISTERS_30_0_port, A2 => n4609, B1 => 
                           REGISTERS_17_0_port, B2 => n4608, ZN => n4616);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_31_0_port, A2 => n4611, B1 => 
                           REGISTERS_23_0_port, B2 => n4610, ZN => n4615);
   U2829 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n4613, B1 => 
                           REGISTERS_24_0_port, B2 => n4612, ZN => n4614);
   U2830 : NAND4_X1 port map( A1 => n4617, A2 => n4616, A3 => n4615, A4 => 
                           n4614, ZN => n4618);
   U2831 : NOR2_X1 port map( A1 => n4619, A2 => n4618, ZN => n4646);
   U2832 : AOI22_X1 port map( A1 => REGISTERS_2_0_port, A2 => n4631, B1 => 
                           REGISTERS_0_0_port, B2 => n4620, ZN => n4628);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n4632, B1 => 
                           REGISTERS_4_0_port, B2 => n4636, ZN => n4627);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_6_0_port, A2 => n4622, B1 => 
                           REGISTERS_1_0_port, B2 => n4621, ZN => n4626);
   U2835 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n4624, B1 => 
                           REGISTERS_3_0_port, B2 => n4623, ZN => n4625);
   U2836 : NAND4_X1 port map( A1 => n4628, A2 => n4627, A3 => n4626, A4 => 
                           n4625, ZN => n4643);
   U2837 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n4630, B1 => 
                           REGISTERS_14_0_port, B2 => n4629, ZN => n4640);
   U2838 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n4632, B1 => 
                           REGISTERS_10_0_port, B2 => n4631, ZN => n4639);
   U2839 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n4634, B1 => 
                           REGISTERS_9_0_port, B2 => n4633, ZN => n4638);
   U2840 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n4636, B1 => 
                           REGISTERS_15_0_port, B2 => n4635, ZN => n4637);
   U2841 : NAND4_X1 port map( A1 => n4640, A2 => n4639, A3 => n4638, A4 => 
                           n4637, ZN => n4641);
   U2842 : AOI22_X1 port map( A1 => n4644, A2 => n4643, B1 => n4642, B2 => 
                           n4641, ZN => n4645);
   U2843 : OAI21_X1 port map( B1 => n4647, B2 => n4646, A => n4645, ZN => N385)
                           ;

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ENABLE_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, curr_instruction_to_cu_i_31_port, 
      curr_instruction_to_cu_i_30_port, curr_instruction_to_cu_i_29_port, 
      curr_instruction_to_cu_i_28_port, curr_instruction_to_cu_i_27_port, 
      curr_instruction_to_cu_i_26_port, curr_instruction_to_cu_i_20_port, 
      curr_instruction_to_cu_i_19_port, curr_instruction_to_cu_i_18_port, 
      curr_instruction_to_cu_i_17_port, curr_instruction_to_cu_i_16_port, 
      curr_instruction_to_cu_i_15_port, curr_instruction_to_cu_i_14_port, 
      curr_instruction_to_cu_i_13_port, curr_instruction_to_cu_i_12_port, 
      curr_instruction_to_cu_i_11_port, curr_instruction_to_cu_i_5_port, 
      curr_instruction_to_cu_i_4_port, curr_instruction_to_cu_i_3_port, 
      curr_instruction_to_cu_i_2_port, curr_instruction_to_cu_i_1_port, 
      curr_instruction_to_cu_i_0_port, enable_rf_i, read_rf_p2_i, alu_cin_i, 
      write_rf_i, cu_i_n134, cu_i_n132, cu_i_n131, cu_i_n127, cu_i_n126, 
      cu_i_n125, cu_i_n124, cu_i_n123, cu_i_n4, cu_i_n210, cu_i_n209, cu_i_n145
      , cu_i_n26, cu_i_n25, cu_i_n23, cu_i_cw1_i_4_port, cu_i_cw1_i_7_port, 
      cu_i_cw1_i_8_port, cu_i_cw3_6_port, cu_i_cw2_4_port, cu_i_cw2_5_port, 
      cu_i_cw2_6_port, cu_i_cw2_7_port, cu_i_cw2_8_port, cu_i_cw1_0_port, 
      cu_i_cw1_1_port, cu_i_cw1_2_port, cu_i_cw1_3_port, cu_i_cw1_4_port, 
      cu_i_cw1_5_port, cu_i_cw1_6_port, cu_i_cw1_7_port, cu_i_cw1_8_port, 
      cu_i_cw1_10_port, cu_i_cw1_11_port, cu_i_cw1_12_port, cu_i_cw1_13_port, 
      cu_i_N279, cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, 
      cu_i_N273, cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, 
      cu_i_cmd_alu_op_type_0_port, cu_i_cmd_alu_op_type_1_port, 
      cu_i_cmd_alu_op_type_2_port, cu_i_cmd_alu_op_type_3_port, 
      cu_i_cmd_word_1_port, cu_i_cmd_word_3_port, cu_i_cmd_word_4_port, 
      cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, cu_i_cmd_word_8_port, 
      cu_i_next_stall, cu_i_next_val_counter_mul_0_port, 
      cu_i_next_val_counter_mul_1_port, cu_i_next_val_counter_mul_2_port, 
      cu_i_next_val_counter_mul_3_port, datapath_i_data_from_alu_i_0_port, 
      datapath_i_data_from_alu_i_1_port, datapath_i_data_from_alu_i_2_port, 
      datapath_i_data_from_alu_i_3_port, datapath_i_data_from_alu_i_4_port, 
      datapath_i_data_from_alu_i_5_port, datapath_i_data_from_alu_i_6_port, 
      datapath_i_data_from_alu_i_7_port, datapath_i_data_from_alu_i_8_port, 
      datapath_i_data_from_alu_i_9_port, datapath_i_data_from_alu_i_10_port, 
      datapath_i_data_from_alu_i_11_port, datapath_i_data_from_alu_i_12_port, 
      datapath_i_data_from_alu_i_13_port, datapath_i_data_from_alu_i_14_port, 
      datapath_i_data_from_alu_i_15_port, datapath_i_data_from_alu_i_16_port, 
      datapath_i_data_from_alu_i_17_port, datapath_i_data_from_alu_i_18_port, 
      datapath_i_data_from_alu_i_19_port, datapath_i_data_from_alu_i_20_port, 
      datapath_i_data_from_alu_i_21_port, datapath_i_data_from_alu_i_22_port, 
      datapath_i_data_from_alu_i_23_port, datapath_i_data_from_alu_i_24_port, 
      datapath_i_data_from_alu_i_25_port, datapath_i_data_from_alu_i_26_port, 
      datapath_i_data_from_alu_i_27_port, datapath_i_data_from_alu_i_28_port, 
      datapath_i_data_from_alu_i_29_port, datapath_i_data_from_alu_i_30_port, 
      datapath_i_data_from_alu_i_31_port, datapath_i_data_from_memory_i_0_port,
      datapath_i_data_from_memory_i_1_port, 
      datapath_i_data_from_memory_i_2_port, 
      datapath_i_data_from_memory_i_3_port, 
      datapath_i_data_from_memory_i_4_port, 
      datapath_i_data_from_memory_i_5_port, 
      datapath_i_data_from_memory_i_6_port, 
      datapath_i_data_from_memory_i_7_port, 
      datapath_i_data_from_memory_i_8_port, 
      datapath_i_data_from_memory_i_9_port, 
      datapath_i_data_from_memory_i_10_port, 
      datapath_i_data_from_memory_i_11_port, 
      datapath_i_data_from_memory_i_12_port, 
      datapath_i_data_from_memory_i_13_port, 
      datapath_i_data_from_memory_i_14_port, 
      datapath_i_data_from_memory_i_15_port, 
      datapath_i_data_from_memory_i_16_port, 
      datapath_i_data_from_memory_i_17_port, 
      datapath_i_data_from_memory_i_18_port, 
      datapath_i_data_from_memory_i_19_port, 
      datapath_i_data_from_memory_i_20_port, 
      datapath_i_data_from_memory_i_21_port, 
      datapath_i_data_from_memory_i_22_port, 
      datapath_i_data_from_memory_i_23_port, 
      datapath_i_data_from_memory_i_24_port, 
      datapath_i_data_from_memory_i_25_port, 
      datapath_i_data_from_memory_i_26_port, 
      datapath_i_data_from_memory_i_27_port, 
      datapath_i_data_from_memory_i_28_port, 
      datapath_i_data_from_memory_i_29_port, 
      datapath_i_data_from_memory_i_30_port, 
      datapath_i_data_from_memory_i_31_port, datapath_i_value_to_mem_i_0_port, 
      datapath_i_value_to_mem_i_1_port, datapath_i_value_to_mem_i_2_port, 
      datapath_i_value_to_mem_i_3_port, datapath_i_value_to_mem_i_4_port, 
      datapath_i_value_to_mem_i_5_port, datapath_i_value_to_mem_i_6_port, 
      datapath_i_value_to_mem_i_7_port, datapath_i_value_to_mem_i_8_port, 
      datapath_i_value_to_mem_i_9_port, datapath_i_value_to_mem_i_10_port, 
      datapath_i_value_to_mem_i_11_port, datapath_i_value_to_mem_i_12_port, 
      datapath_i_value_to_mem_i_13_port, datapath_i_value_to_mem_i_14_port, 
      datapath_i_value_to_mem_i_15_port, datapath_i_value_to_mem_i_16_port, 
      datapath_i_value_to_mem_i_17_port, datapath_i_value_to_mem_i_18_port, 
      datapath_i_value_to_mem_i_19_port, datapath_i_value_to_mem_i_20_port, 
      datapath_i_value_to_mem_i_21_port, datapath_i_value_to_mem_i_22_port, 
      datapath_i_value_to_mem_i_23_port, datapath_i_value_to_mem_i_24_port, 
      datapath_i_value_to_mem_i_25_port, datapath_i_value_to_mem_i_26_port, 
      datapath_i_value_to_mem_i_27_port, datapath_i_value_to_mem_i_28_port, 
      datapath_i_value_to_mem_i_29_port, datapath_i_value_to_mem_i_30_port, 
      datapath_i_value_to_mem_i_31_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, datapath_i_val_immediate_i_0_port, 
      datapath_i_val_immediate_i_1_port, datapath_i_val_immediate_i_2_port, 
      datapath_i_val_immediate_i_3_port, datapath_i_val_immediate_i_4_port, 
      datapath_i_val_immediate_i_5_port, datapath_i_val_immediate_i_6_port, 
      datapath_i_val_immediate_i_7_port, datapath_i_val_immediate_i_8_port, 
      datapath_i_val_immediate_i_9_port, datapath_i_val_immediate_i_10_port, 
      datapath_i_val_immediate_i_11_port, datapath_i_val_immediate_i_12_port, 
      datapath_i_val_immediate_i_13_port, datapath_i_val_immediate_i_14_port, 
      datapath_i_val_immediate_i_15_port, datapath_i_val_immediate_i_16_port, 
      datapath_i_val_immediate_i_17_port, datapath_i_val_immediate_i_18_port, 
      datapath_i_val_immediate_i_19_port, datapath_i_val_immediate_i_20_port, 
      datapath_i_val_immediate_i_21_port, datapath_i_val_immediate_i_22_port, 
      datapath_i_val_immediate_i_23_port, datapath_i_val_immediate_i_24_port, 
      datapath_i_val_immediate_i_25_port, datapath_i_val_b_i_0_port, 
      datapath_i_val_b_i_1_port, datapath_i_val_b_i_2_port, 
      datapath_i_val_b_i_3_port, datapath_i_val_b_i_4_port, 
      datapath_i_val_b_i_5_port, datapath_i_val_b_i_6_port, 
      datapath_i_val_b_i_7_port, datapath_i_val_b_i_8_port, 
      datapath_i_val_b_i_9_port, datapath_i_val_b_i_10_port, 
      datapath_i_val_b_i_11_port, datapath_i_val_b_i_12_port, 
      datapath_i_val_b_i_13_port, datapath_i_val_b_i_14_port, 
      datapath_i_val_b_i_15_port, datapath_i_val_b_i_16_port, 
      datapath_i_val_b_i_17_port, datapath_i_val_b_i_18_port, 
      datapath_i_val_b_i_19_port, datapath_i_val_b_i_20_port, 
      datapath_i_val_b_i_21_port, datapath_i_val_b_i_22_port, 
      datapath_i_val_b_i_23_port, datapath_i_val_b_i_24_port, 
      datapath_i_val_b_i_25_port, datapath_i_val_b_i_26_port, 
      datapath_i_val_b_i_27_port, datapath_i_val_b_i_28_port, 
      datapath_i_val_b_i_29_port, datapath_i_val_b_i_30_port, 
      datapath_i_val_b_i_31_port, datapath_i_val_a_i_0_port, 
      datapath_i_val_a_i_1_port, datapath_i_val_a_i_2_port, 
      datapath_i_val_a_i_3_port, datapath_i_val_a_i_4_port, 
      datapath_i_val_a_i_5_port, datapath_i_val_a_i_6_port, 
      datapath_i_val_a_i_7_port, datapath_i_val_a_i_8_port, 
      datapath_i_val_a_i_9_port, datapath_i_val_a_i_10_port, 
      datapath_i_val_a_i_11_port, datapath_i_val_a_i_12_port, 
      datapath_i_val_a_i_13_port, datapath_i_val_a_i_14_port, 
      datapath_i_val_a_i_15_port, datapath_i_val_a_i_16_port, 
      datapath_i_val_a_i_17_port, datapath_i_val_a_i_18_port, 
      datapath_i_val_a_i_19_port, datapath_i_val_a_i_20_port, 
      datapath_i_val_a_i_21_port, datapath_i_val_a_i_22_port, 
      datapath_i_val_a_i_23_port, datapath_i_val_a_i_24_port, 
      datapath_i_val_a_i_25_port, datapath_i_val_a_i_26_port, 
      datapath_i_val_a_i_27_port, datapath_i_val_a_i_28_port, 
      datapath_i_val_a_i_29_port, datapath_i_val_a_i_30_port, 
      datapath_i_val_a_i_31_port, datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_branch_condition_i_0_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_5_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_7_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_9_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_11_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_13_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_15_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_17_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_19_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_21_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_23_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_25_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_27_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_29_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, 
      datapath_i_new_pc_value_mem_stage_i_31_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_n69, 
      datapath_i_fetch_stage_dp_n68, datapath_i_fetch_stage_dp_n67, 
      datapath_i_fetch_stage_dp_n66, datapath_i_fetch_stage_dp_n65, 
      datapath_i_fetch_stage_dp_n64, datapath_i_fetch_stage_dp_n63, 
      datapath_i_fetch_stage_dp_n62, datapath_i_fetch_stage_dp_n61, 
      datapath_i_fetch_stage_dp_n60, datapath_i_fetch_stage_dp_n59, 
      datapath_i_fetch_stage_dp_n58, datapath_i_fetch_stage_dp_n57, 
      datapath_i_fetch_stage_dp_n56, datapath_i_fetch_stage_dp_n55, 
      datapath_i_fetch_stage_dp_n54, datapath_i_fetch_stage_dp_n53, 
      datapath_i_fetch_stage_dp_n52, datapath_i_fetch_stage_dp_n51, 
      datapath_i_fetch_stage_dp_n50, datapath_i_fetch_stage_dp_n49, 
      datapath_i_fetch_stage_dp_n48, datapath_i_fetch_stage_dp_n47, 
      datapath_i_fetch_stage_dp_n46, datapath_i_fetch_stage_dp_n45, 
      datapath_i_fetch_stage_dp_n44, datapath_i_fetch_stage_dp_n43, 
      datapath_i_fetch_stage_dp_n42, datapath_i_fetch_stage_dp_n41, 
      datapath_i_fetch_stage_dp_n40, datapath_i_fetch_stage_dp_n39, 
      datapath_i_fetch_stage_dp_n38, datapath_i_fetch_stage_dp_n37, 
      datapath_i_fetch_stage_dp_n36, datapath_i_fetch_stage_dp_n35, 
      datapath_i_fetch_stage_dp_n34, datapath_i_fetch_stage_dp_n33, 
      datapath_i_fetch_stage_dp_n32, datapath_i_fetch_stage_dp_n31, 
      datapath_i_fetch_stage_dp_n30, datapath_i_fetch_stage_dp_n29, 
      datapath_i_fetch_stage_dp_n28, datapath_i_fetch_stage_dp_n27, 
      datapath_i_fetch_stage_dp_n26, datapath_i_fetch_stage_dp_n25, 
      datapath_i_fetch_stage_dp_n24, datapath_i_fetch_stage_dp_n23, 
      datapath_i_fetch_stage_dp_n22, datapath_i_fetch_stage_dp_n21, 
      datapath_i_fetch_stage_dp_n20, datapath_i_fetch_stage_dp_n19, 
      datapath_i_fetch_stage_dp_n18, datapath_i_fetch_stage_dp_n17, 
      datapath_i_fetch_stage_dp_n16, datapath_i_fetch_stage_dp_n15, 
      datapath_i_fetch_stage_dp_n14, datapath_i_fetch_stage_dp_n13, 
      datapath_i_fetch_stage_dp_n12, datapath_i_fetch_stage_dp_n11, 
      datapath_i_fetch_stage_dp_n10, datapath_i_fetch_stage_dp_n9, 
      datapath_i_fetch_stage_dp_n4, datapath_i_fetch_stage_dp_n3, 
      datapath_i_fetch_stage_dp_n2, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port, datapath_i_fetch_stage_dp_N6, 
      datapath_i_fetch_stage_dp_N5, datapath_i_decode_stage_dp_n80, 
      datapath_i_decode_stage_dp_n79, datapath_i_decode_stage_dp_n78, 
      datapath_i_decode_stage_dp_n77, datapath_i_decode_stage_dp_n76, 
      datapath_i_decode_stage_dp_n43, datapath_i_decode_stage_dp_n42, 
      datapath_i_decode_stage_dp_n41, datapath_i_decode_stage_dp_n40, 
      datapath_i_decode_stage_dp_n39, datapath_i_decode_stage_dp_n38, 
      datapath_i_decode_stage_dp_n37, datapath_i_decode_stage_dp_n36, 
      datapath_i_decode_stage_dp_n35, datapath_i_decode_stage_dp_n34, 
      datapath_i_decode_stage_dp_n33, datapath_i_decode_stage_dp_n32, 
      datapath_i_decode_stage_dp_n31, datapath_i_decode_stage_dp_n30, 
      datapath_i_decode_stage_dp_n29, datapath_i_decode_stage_dp_n28, 
      datapath_i_decode_stage_dp_n27, datapath_i_decode_stage_dp_n26, 
      datapath_i_decode_stage_dp_n25, datapath_i_decode_stage_dp_n24, 
      datapath_i_decode_stage_dp_n23, datapath_i_decode_stage_dp_n22, 
      datapath_i_decode_stage_dp_n21, datapath_i_decode_stage_dp_n20, 
      datapath_i_decode_stage_dp_n19, datapath_i_decode_stage_dp_n18, 
      datapath_i_decode_stage_dp_n17, datapath_i_decode_stage_dp_n16, 
      datapath_i_decode_stage_dp_n15, datapath_i_decode_stage_dp_n14, 
      datapath_i_decode_stage_dp_n13, datapath_i_decode_stage_dp_n12, 
      datapath_i_decode_stage_dp_pc_delay3_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_1_port, 
      datapath_i_decode_stage_dp_pc_delay2_2_port, 
      datapath_i_decode_stage_dp_pc_delay2_3_port, 
      datapath_i_decode_stage_dp_pc_delay2_4_port, 
      datapath_i_decode_stage_dp_pc_delay2_5_port, 
      datapath_i_decode_stage_dp_pc_delay2_6_port, 
      datapath_i_decode_stage_dp_pc_delay2_7_port, 
      datapath_i_decode_stage_dp_pc_delay2_8_port, 
      datapath_i_decode_stage_dp_pc_delay2_9_port, 
      datapath_i_decode_stage_dp_pc_delay2_10_port, 
      datapath_i_decode_stage_dp_pc_delay2_11_port, 
      datapath_i_decode_stage_dp_pc_delay2_12_port, 
      datapath_i_decode_stage_dp_pc_delay2_13_port, 
      datapath_i_decode_stage_dp_pc_delay2_14_port, 
      datapath_i_decode_stage_dp_pc_delay2_15_port, 
      datapath_i_decode_stage_dp_pc_delay2_16_port, 
      datapath_i_decode_stage_dp_pc_delay2_17_port, 
      datapath_i_decode_stage_dp_pc_delay2_18_port, 
      datapath_i_decode_stage_dp_pc_delay2_19_port, 
      datapath_i_decode_stage_dp_pc_delay2_20_port, 
      datapath_i_decode_stage_dp_pc_delay2_21_port, 
      datapath_i_decode_stage_dp_pc_delay2_22_port, 
      datapath_i_decode_stage_dp_pc_delay2_23_port, 
      datapath_i_decode_stage_dp_pc_delay2_24_port, 
      datapath_i_decode_stage_dp_pc_delay2_25_port, 
      datapath_i_decode_stage_dp_pc_delay2_26_port, 
      datapath_i_decode_stage_dp_pc_delay2_27_port, 
      datapath_i_decode_stage_dp_pc_delay2_28_port, 
      datapath_i_decode_stage_dp_pc_delay2_29_port, 
      datapath_i_decode_stage_dp_pc_delay2_30_port, 
      datapath_i_decode_stage_dp_pc_delay2_31_port, 
      datapath_i_decode_stage_dp_pc_delay2_32_port, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_0_port, 
      datapath_i_decode_stage_dp_address_rf_write_1_port, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_decode_stage_dp_address_rf_write_3_port, 
      datapath_i_decode_stage_dp_address_rf_write_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
      datapath_i_decode_stage_dp_enable_sign_extension_logic, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_out_0_port, 
      datapath_i_execute_stage_dp_alu_out_1_port, 
      datapath_i_execute_stage_dp_alu_out_2_port, 
      datapath_i_execute_stage_dp_alu_out_3_port, 
      datapath_i_execute_stage_dp_alu_out_4_port, 
      datapath_i_execute_stage_dp_alu_out_5_port, 
      datapath_i_execute_stage_dp_alu_out_6_port, 
      datapath_i_execute_stage_dp_alu_out_7_port, 
      datapath_i_execute_stage_dp_alu_out_8_port, 
      datapath_i_execute_stage_dp_alu_out_9_port, 
      datapath_i_execute_stage_dp_alu_out_10_port, 
      datapath_i_execute_stage_dp_alu_out_11_port, 
      datapath_i_execute_stage_dp_alu_out_12_port, 
      datapath_i_execute_stage_dp_alu_out_13_port, 
      datapath_i_execute_stage_dp_alu_out_14_port, 
      datapath_i_execute_stage_dp_alu_out_15_port, 
      datapath_i_execute_stage_dp_alu_out_16_port, 
      datapath_i_execute_stage_dp_alu_out_17_port, 
      datapath_i_execute_stage_dp_alu_out_18_port, 
      datapath_i_execute_stage_dp_alu_out_19_port, 
      datapath_i_execute_stage_dp_alu_out_20_port, 
      datapath_i_execute_stage_dp_alu_out_21_port, 
      datapath_i_execute_stage_dp_alu_out_22_port, 
      datapath_i_execute_stage_dp_alu_out_23_port, 
      datapath_i_execute_stage_dp_alu_out_24_port, 
      datapath_i_execute_stage_dp_alu_out_25_port, 
      datapath_i_execute_stage_dp_alu_out_26_port, 
      datapath_i_execute_stage_dp_alu_out_27_port, 
      datapath_i_execute_stage_dp_alu_out_28_port, 
      datapath_i_execute_stage_dp_alu_out_29_port, 
      datapath_i_execute_stage_dp_alu_out_30_port, 
      datapath_i_execute_stage_dp_alu_out_31_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_3_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, 
      datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
      datapath_i_memory_stage_dp_n2, datapath_i_memory_stage_dp_data_ir_0_port,
      datapath_i_memory_stage_dp_data_ir_1_port, 
      datapath_i_memory_stage_dp_data_ir_2_port, 
      datapath_i_memory_stage_dp_data_ir_3_port, 
      datapath_i_memory_stage_dp_data_ir_4_port, 
      datapath_i_memory_stage_dp_data_ir_5_port, 
      datapath_i_memory_stage_dp_data_ir_6_port, 
      datapath_i_memory_stage_dp_data_ir_7_port, 
      datapath_i_memory_stage_dp_data_ir_8_port, 
      datapath_i_memory_stage_dp_data_ir_9_port, 
      datapath_i_memory_stage_dp_data_ir_10_port, 
      datapath_i_memory_stage_dp_data_ir_11_port, 
      datapath_i_memory_stage_dp_data_ir_12_port, 
      datapath_i_memory_stage_dp_data_ir_13_port, 
      datapath_i_memory_stage_dp_data_ir_14_port, 
      datapath_i_memory_stage_dp_data_ir_15_port, 
      datapath_i_memory_stage_dp_data_ir_16_port, 
      datapath_i_memory_stage_dp_data_ir_17_port, 
      datapath_i_memory_stage_dp_data_ir_18_port, 
      datapath_i_memory_stage_dp_data_ir_19_port, 
      datapath_i_memory_stage_dp_data_ir_20_port, 
      datapath_i_memory_stage_dp_data_ir_21_port, 
      datapath_i_memory_stage_dp_data_ir_22_port, 
      datapath_i_memory_stage_dp_data_ir_23_port, 
      datapath_i_memory_stage_dp_data_ir_24_port, 
      datapath_i_memory_stage_dp_data_ir_25_port, 
      datapath_i_memory_stage_dp_data_ir_26_port, 
      datapath_i_memory_stage_dp_data_ir_27_port, 
      datapath_i_memory_stage_dp_data_ir_28_port, 
      datapath_i_memory_stage_dp_data_ir_29_port, 
      datapath_i_memory_stage_dp_data_ir_30_port, 
      datapath_i_memory_stage_dp_data_ir_31_port, n309, n310, n311, n313, n314,
      n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
      n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
      n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
      n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
      n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
      n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, 
      n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, 
      n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, 
      n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
      n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
      n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
      n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, DRAM_ENABLE_port, n768, 
      n769, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   DRAM_ENABLE <= DRAM_ENABLE_port;
   
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_counter_mul_reg_1_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_1_port, CK => CLK, RN => 
                           RST, Q => n735, QN => cu_i_n26);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_next_val_counter_mul_1_port);
   cu_i_counter_mul_reg_2_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_2_port, CK => CLK, RN => 
                           RST, Q => n754, QN => cu_i_n25);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_next_val_counter_mul_2_port);
   cu_i_counter_mul_reg_3_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_3_port, CK => CLK, RN => 
                           RST, Q => n738, QN => cu_i_n124);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_next_val_counter_mul_3_port);
   cu_i_counter_mul_reg_0_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_0_port, CK => CLK, RN => 
                           RST, Q => n694, QN => cu_i_n125);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_next_val_counter_mul_0_port);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => cu_i_n145, Q => 
                           cu_i_next_stall);
   cu_i_curr_state_reg_1_inst : DFFR_X1 port map( D => cu_i_n209, CK => CLK, RN
                           => RST, Q => n_1422, QN => cu_i_n123);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           ADD_WR(3) => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           ADD_WR(2) => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ADD_WR(1) => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ADD_WR(0) => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n12, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n43, OUT1(31) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
                           OUT1(30) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
                           OUT1(29) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
                           OUT1(28) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
                           OUT1(27) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
                           OUT1(26) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
                           OUT1(25) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
                           OUT1(24) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
                           OUT1(23) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
                           OUT1(22) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
                           OUT1(21) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
                           OUT1(20) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
                           OUT1(19) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
                           OUT1(18) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
                           OUT1(17) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
                           OUT1(16) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
                           OUT1(15) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
                           OUT1(14) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
                           OUT1(13) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
                           OUT1(12) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
                           OUT1(11) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
                           OUT1(10) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
                           OUT1(9) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
                           OUT1(8) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
                           OUT1(7) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
                           OUT1(6) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
                           OUT1(5) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
                           OUT1(4) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
                           OUT1(3) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
                           OUT1(2) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
                           OUT1(1) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
                           OUT1(0) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
                           OUT2(31) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
                           OUT2(30) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
                           OUT2(29) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
                           OUT2(28) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
                           OUT2(27) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
                           OUT2(26) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
                           OUT2(25) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
                           OUT2(24) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
                           OUT2(23) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
                           OUT2(22) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
                           OUT2(21) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
                           OUT2(20) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
                           OUT2(19) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
                           OUT2(18) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
                           OUT2(17) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
                           OUT2(16) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
                           OUT2(15) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
                           OUT2(14) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
                           OUT2(13) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
                           OUT2(12) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
                           OUT2(11) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
                           OUT2(10) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
                           OUT2(9) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
                           OUT2(8) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
                           OUT2(7) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
                           OUT2(6) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
                           OUT2(5) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
                           OUT2(4) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
                           OUT2(3) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
                           OUT2(2) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
                           OUT2(1) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
                           OUT2(0) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
                           RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_1423, mul_exeception => 
                           n_1424, FUNC(0) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_3_port, 
                           FUNC(1) => datapath_i_execute_stage_dp_n7, FUNC(2) 
                           => datapath_i_execute_stage_dp_alu_op_type_i_1_port,
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_1425, 
                           OUTALU(31) => 
                           datapath_i_execute_stage_dp_alu_out_31_port, 
                           OUTALU(30) => 
                           datapath_i_execute_stage_dp_alu_out_30_port, 
                           OUTALU(29) => 
                           datapath_i_execute_stage_dp_alu_out_29_port, 
                           OUTALU(28) => 
                           datapath_i_execute_stage_dp_alu_out_28_port, 
                           OUTALU(27) => 
                           datapath_i_execute_stage_dp_alu_out_27_port, 
                           OUTALU(26) => 
                           datapath_i_execute_stage_dp_alu_out_26_port, 
                           OUTALU(25) => 
                           datapath_i_execute_stage_dp_alu_out_25_port, 
                           OUTALU(24) => 
                           datapath_i_execute_stage_dp_alu_out_24_port, 
                           OUTALU(23) => 
                           datapath_i_execute_stage_dp_alu_out_23_port, 
                           OUTALU(22) => 
                           datapath_i_execute_stage_dp_alu_out_22_port, 
                           OUTALU(21) => 
                           datapath_i_execute_stage_dp_alu_out_21_port, 
                           OUTALU(20) => 
                           datapath_i_execute_stage_dp_alu_out_20_port, 
                           OUTALU(19) => 
                           datapath_i_execute_stage_dp_alu_out_19_port, 
                           OUTALU(18) => 
                           datapath_i_execute_stage_dp_alu_out_18_port, 
                           OUTALU(17) => 
                           datapath_i_execute_stage_dp_alu_out_17_port, 
                           OUTALU(16) => 
                           datapath_i_execute_stage_dp_alu_out_16_port, 
                           OUTALU(15) => 
                           datapath_i_execute_stage_dp_alu_out_15_port, 
                           OUTALU(14) => 
                           datapath_i_execute_stage_dp_alu_out_14_port, 
                           OUTALU(13) => 
                           datapath_i_execute_stage_dp_alu_out_13_port, 
                           OUTALU(12) => 
                           datapath_i_execute_stage_dp_alu_out_12_port, 
                           OUTALU(11) => 
                           datapath_i_execute_stage_dp_alu_out_11_port, 
                           OUTALU(10) => 
                           datapath_i_execute_stage_dp_alu_out_10_port, 
                           OUTALU(9) => 
                           datapath_i_execute_stage_dp_alu_out_9_port, 
                           OUTALU(8) => 
                           datapath_i_execute_stage_dp_alu_out_8_port, 
                           OUTALU(7) => 
                           datapath_i_execute_stage_dp_alu_out_7_port, 
                           OUTALU(6) => 
                           datapath_i_execute_stage_dp_alu_out_6_port, 
                           OUTALU(5) => 
                           datapath_i_execute_stage_dp_alu_out_5_port, 
                           OUTALU(4) => 
                           datapath_i_execute_stage_dp_alu_out_4_port, 
                           OUTALU(3) => 
                           datapath_i_execute_stage_dp_alu_out_3_port, 
                           OUTALU(2) => 
                           datapath_i_execute_stage_dp_alu_out_2_port, 
                           OUTALU(1) => 
                           datapath_i_execute_stage_dp_alu_out_1_port, 
                           OUTALU(0) => 
                           datapath_i_execute_stage_dp_alu_out_0_port, rst_BAR 
                           => RST);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n766, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n766, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n766, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n766, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n766, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n766, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n766, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n766, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n766, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n766, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n766, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n309, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n766, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n309, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n766, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n309, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n766, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n309, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n766, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n309, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n309, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n309, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n309, Z =>
                           DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n309, Z =>
                           DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n766, Z =>
                           DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n766, Z =>
                           DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n766, Z =>
                           DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n766, Z =>
                           DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n766, Z =>
                           DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n766, Z =>
                           DRAM_ADDRESS_2_port);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_9_port, EN => n768, Z => 
                           DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_31_port, EN => n768, Z => 
                           DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_30_port, EN => n768, Z => 
                           DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_29_port, EN => n768, Z => 
                           DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_28_port, EN => n768, Z => 
                           DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_27_port, EN => n768, Z => 
                           DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_26_port, EN => n768, Z => 
                           DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_25_port, EN => n768, Z => 
                           DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_24_port, EN => n768, Z => 
                           DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_23_port, EN => n768, Z => 
                           DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_22_port, EN => n768, Z => 
                           DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_21_port, EN => n768, Z => 
                           DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_20_port, EN => n768, Z => 
                           DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_19_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_18_port, EN => n768, Z => 
                           DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_17_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_16_port, EN => n768, Z => 
                           DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_15_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_14_port, EN => n768, Z => 
                           DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_13_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_12_port, EN => n768, Z => 
                           DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_11_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_10_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_8_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_7_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_6_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_5_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_4_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_3_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_2_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_1_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_0_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(0));
   cu_i_e_reg_D_I_0_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_0_port, QN => 
                           n_1426);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n765, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n765, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n765, D => datapath_i_n18, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n310, D => datapath_i_n17, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n765, D => datapath_i_n16, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n765, D => datapath_i_n15, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n310, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n769, D => datapath_i_n18, Q
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n17, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n769, D => datapath_i_n16, Q
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n15, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n769, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_16_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_17_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_18_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n769, D => 
                           curr_instruction_to_cu_i_19_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => curr_instruction_to_cu_i_20_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n769, D => datapath_i_n13, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n12, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n769, D => datapath_i_n11, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, D 
                           => datapath_i_n10, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n769, D => datapath_i_n9, Q =>
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   cu_i_wb_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n132, CK => CLK, RN =>
                           RST, Q => cu_i_cw3_6_port, QN => n_1427);
   cu_i_wb_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n131, CK => CLK, RN =>
                           RST, Q => n_1428, QN => n699);
   cu_i_m_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_8_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_8_port, QN => n_1429);
   cu_i_m_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_7_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_7_port, QN => n_1430);
   cu_i_m_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n127, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_6_port, QN => n_1431);
   cu_i_m_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n126, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_5_port, QN => n757);
   cu_i_m_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_4_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_4_port, QN => n756);
   cu_i_e_reg_D_I_13_Q_reg : DFFR_X1 port map( D => n310, CK => CLK, RN => RST,
                           Q => cu_i_cw1_13_port, QN => n_1432);
   cu_i_e_reg_D_I_12_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_12_port, QN => n_1433)
                           ;
   cu_i_e_reg_D_I_11_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_11_port, QN => n_1434)
                           ;
   cu_i_e_reg_D_I_10_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_10_port, QN => n_1435)
                           ;
   cu_i_e_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_8_port, QN => n_1436);
   cu_i_e_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_7_port, QN => n_1437);
   cu_i_e_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n311, CK => CLK, RN => RST, 
                           Q => cu_i_cw1_6_port, QN => n_1438);
   cu_i_e_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_1_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_5_port, QN => n_1439);
   cu_i_e_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_n134, CK => CLK, RN => 
                           RST, Q => cu_i_cw1_4_port, QN => n_1440);
   cu_i_e_reg_D_I_3_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_3_port, QN => 
                           n_1441);
   cu_i_e_reg_D_I_2_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_2_port, QN => 
                           n_1442);
   cu_i_e_reg_D_I_1_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_1_port, QN => 
                           n_1443);
   datapath_i_memory_stage_dp_delay_regg_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_31_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_31_port, QN 
                           => n_1444);
   datapath_i_memory_stage_dp_delay_regg_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_30_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_30_port, QN 
                           => n_1445);
   datapath_i_memory_stage_dp_delay_regg_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_29_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_29_port, QN 
                           => n_1446);
   datapath_i_memory_stage_dp_delay_regg_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_28_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_28_port, QN 
                           => n_1447);
   datapath_i_memory_stage_dp_delay_regg_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_27_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_27_port, QN 
                           => n_1448);
   datapath_i_memory_stage_dp_delay_regg_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_26_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_26_port, QN 
                           => n_1449);
   datapath_i_memory_stage_dp_delay_regg_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_25_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_25_port, QN 
                           => n_1450);
   datapath_i_memory_stage_dp_delay_regg_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_24_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_24_port, QN 
                           => n_1451);
   datapath_i_memory_stage_dp_delay_regg_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_23_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_23_port, QN 
                           => n_1452);
   datapath_i_memory_stage_dp_delay_regg_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_22_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_22_port, QN 
                           => n_1453);
   datapath_i_memory_stage_dp_delay_regg_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_21_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_21_port, QN 
                           => n_1454);
   datapath_i_memory_stage_dp_delay_regg_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_20_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_20_port, QN 
                           => n_1455);
   datapath_i_memory_stage_dp_delay_regg_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_19_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_19_port, QN 
                           => n_1456);
   datapath_i_memory_stage_dp_delay_regg_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_18_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_18_port, QN 
                           => n_1457);
   datapath_i_memory_stage_dp_delay_regg_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_17_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_17_port, QN 
                           => n_1458);
   datapath_i_memory_stage_dp_delay_regg_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_16_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_16_port, QN 
                           => n_1459);
   datapath_i_memory_stage_dp_delay_regg_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_15_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_15_port, QN 
                           => n_1460);
   datapath_i_memory_stage_dp_delay_regg_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_14_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_14_port, QN 
                           => n_1461);
   datapath_i_memory_stage_dp_delay_regg_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_13_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_13_port, QN 
                           => n_1462);
   datapath_i_memory_stage_dp_delay_regg_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_12_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_12_port, QN 
                           => n_1463);
   datapath_i_memory_stage_dp_delay_regg_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_11_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_11_port, QN 
                           => n_1464);
   datapath_i_memory_stage_dp_delay_regg_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_10_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_10_port, QN 
                           => n_1465);
   datapath_i_memory_stage_dp_delay_regg_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_9_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_9_port, QN => 
                           n_1466);
   datapath_i_memory_stage_dp_delay_regg_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_8_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_8_port, QN => 
                           n_1467);
   datapath_i_memory_stage_dp_delay_regg_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_7_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_7_port, QN => 
                           n_1468);
   datapath_i_memory_stage_dp_delay_regg_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_6_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_6_port, QN => 
                           n_1469);
   datapath_i_memory_stage_dp_delay_regg_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_5_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_5_port, QN => 
                           n_1470);
   datapath_i_memory_stage_dp_delay_regg_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_4_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_4_port, QN => 
                           n_1471);
   datapath_i_memory_stage_dp_delay_regg_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_3_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_3_port, QN => 
                           n_1472);
   datapath_i_memory_stage_dp_delay_regg_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_2_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_2_port, QN => 
                           n_1473);
   datapath_i_memory_stage_dp_delay_regg_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_1_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_1_port, QN => 
                           n_1474);
   datapath_i_memory_stage_dp_delay_regg_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_0_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_0_port, QN => 
                           n_1475);
   datapath_i_memory_stage_dp_lmd_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_31_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_31_port, QN => n_1476)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_30_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_30_port, QN => n_1477)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_29_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_29_port, QN => n_1478)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_28_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_28_port, QN => n_1479)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_27_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_27_port, QN => n_1480)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_26_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_26_port, QN => n_1481)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_25_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_25_port, QN => n_1482)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_24_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_24_port, QN => n_1483)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_23_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_23_port, QN => n_1484)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_22_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_22_port, QN => n_1485)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_21_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_21_port, QN => n_1486)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_20_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_20_port, QN => n_1487)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_19_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_19_port, QN => n_1488)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_18_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_18_port, QN => n_1489)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_17_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_17_port, QN => n_1490)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_16_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_16_port, QN => n_1491)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_15_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_15_port, QN => n_1492)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_14_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_14_port, QN => n_1493)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_13_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_13_port, QN => n_1494)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_12_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_12_port, QN => n_1495)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_11_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_11_port, QN => n_1496)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_10_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_10_port, QN => n_1497)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_9_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_9_port, QN => n_1498);
   datapath_i_memory_stage_dp_lmd_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_8_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_8_port, QN => n_1499);
   datapath_i_memory_stage_dp_lmd_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_7_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_7_port, QN => n_1500);
   datapath_i_memory_stage_dp_lmd_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_6_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_6_port, QN => n_1501);
   datapath_i_memory_stage_dp_lmd_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_5_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_5_port, QN => n_1502);
   datapath_i_memory_stage_dp_lmd_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_4_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_4_port, QN => n_1503);
   datapath_i_memory_stage_dp_lmd_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_3_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_3_port, QN => n_1504);
   datapath_i_memory_stage_dp_lmd_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_2_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_2_port, QN => n_1505);
   datapath_i_memory_stage_dp_lmd_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_1_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_1_port, QN => n_1506);
   datapath_i_memory_stage_dp_lmd_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_0_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_0_port, QN => n_1507);
   datapath_i_execute_stage_dp_reg_del_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_31_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_31_port, QN => n_1508);
   datapath_i_execute_stage_dp_reg_del_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_30_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_30_port, QN => n_1509);
   datapath_i_execute_stage_dp_reg_del_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_29_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_29_port, QN => n_1510);
   datapath_i_execute_stage_dp_reg_del_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_28_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_28_port, QN => n_1511);
   datapath_i_execute_stage_dp_reg_del_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_27_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_27_port, QN => n_1512);
   datapath_i_execute_stage_dp_reg_del_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_26_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_26_port, QN => n_1513);
   datapath_i_execute_stage_dp_reg_del_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_25_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_25_port, QN => n_1514);
   datapath_i_execute_stage_dp_reg_del_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_24_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_24_port, QN => n_1515);
   datapath_i_execute_stage_dp_reg_del_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_23_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_23_port, QN => n_1516);
   datapath_i_execute_stage_dp_reg_del_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_22_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_22_port, QN => n_1517);
   datapath_i_execute_stage_dp_reg_del_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_21_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_21_port, QN => n_1518);
   datapath_i_execute_stage_dp_reg_del_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_20_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_20_port, QN => n_1519);
   datapath_i_execute_stage_dp_reg_del_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_19_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_19_port, QN => n_1520);
   datapath_i_execute_stage_dp_reg_del_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_18_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_18_port, QN => n_1521);
   datapath_i_execute_stage_dp_reg_del_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_17_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_17_port, QN => n_1522);
   datapath_i_execute_stage_dp_reg_del_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_16_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_16_port, QN => n_1523);
   datapath_i_execute_stage_dp_reg_del_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_15_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_15_port, QN => n_1524);
   datapath_i_execute_stage_dp_reg_del_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_14_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_14_port, QN => n_1525);
   datapath_i_execute_stage_dp_reg_del_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_13_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_13_port, QN => n_1526);
   datapath_i_execute_stage_dp_reg_del_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_12_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_12_port, QN => n_1527);
   datapath_i_execute_stage_dp_reg_del_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_11_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_11_port, QN => n_1528);
   datapath_i_execute_stage_dp_reg_del_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_10_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_10_port, QN => n_1529);
   datapath_i_execute_stage_dp_reg_del_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_9_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_9_port, QN => n_1530);
   datapath_i_execute_stage_dp_reg_del_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_8_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_8_port, QN => n_1531);
   datapath_i_execute_stage_dp_reg_del_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_7_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_7_port, QN => n_1532);
   datapath_i_execute_stage_dp_reg_del_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_6_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_6_port, QN => n_1533);
   datapath_i_execute_stage_dp_reg_del_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_5_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_5_port, QN => n_1534);
   datapath_i_execute_stage_dp_reg_del_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_4_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_4_port, QN => n_1535);
   datapath_i_execute_stage_dp_reg_del_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_3_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_3_port, QN => n_1536);
   datapath_i_execute_stage_dp_reg_del_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_2_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_2_port, QN => n_1537);
   datapath_i_execute_stage_dp_reg_del_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_1_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_1_port, QN => n_1538);
   datapath_i_execute_stage_dp_reg_del_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_0_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_0_port, QN => n_1539);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_31_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_31_port, QN => n_1540);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_30_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_30_port, QN => n_1541);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_29_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_29_port, QN => n_1542);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_28_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_28_port, QN => n_1543);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_27_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_27_port, QN => n_1544);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_26_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_26_port, QN => n_1545);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_25_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_25_port, QN => n_1546);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_24_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_24_port, QN => n_1547);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_23_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_23_port, QN => n_1548);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_22_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_22_port, QN => n_1549);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_21_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_21_port, QN => n_1550);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_20_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_20_port, QN => n_1551);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_19_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_19_port, QN => n_1552);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_18_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_18_port, QN => n_1553);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_17_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_17_port, QN => n_1554);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_16_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_16_port, QN => n_1555);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_15_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_15_port, QN => n_1556);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_14_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_14_port, QN => n_1557);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_13_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_13_port, QN => n_1558);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_12_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_12_port, QN => n_1559);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_11_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_11_port, QN => n_1560);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_10_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_10_port, QN => n_1561);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_9_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_9_port, QN => n_1562);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_8_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_8_port, QN => n_1563);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_7_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_7_port, QN => n_1564);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_6_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_6_port, QN => n_1565);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_5_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_5_port, QN => n_1566);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_4_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_4_port, QN => n_1567);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_3_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_3_port, QN => n_1568);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_2_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_2_port, QN => n_1569);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_1_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_1_port, QN => n_1570);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_0_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_0_port, QN => n_1571);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_32_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_32_port, CK 
                           => CLK, RN => RST, Q => n_1572, QN => n703);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_31_port, CK 
                           => CLK, RN => RST, Q => n_1573, QN => n727);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_30_port, CK 
                           => CLK, RN => RST, Q => n_1574, QN => n726);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_29_port, CK 
                           => CLK, RN => RST, Q => n_1575, QN => n725);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_28_port, CK 
                           => CLK, RN => RST, Q => n_1576, QN => n724);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_27_port, CK 
                           => CLK, RN => RST, Q => n_1577, QN => n691);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_26_port, CK 
                           => CLK, RN => RST, Q => n_1578, QN => n723);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_25_port, CK 
                           => CLK, RN => RST, Q => n_1579, QN => n722);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_24_port, CK 
                           => CLK, RN => RST, Q => n_1580, QN => n721);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_23_port, CK 
                           => CLK, RN => RST, Q => n_1581, QN => n720);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_22_port, CK 
                           => CLK, RN => RST, Q => n_1582, QN => n719);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_21_port, CK 
                           => CLK, RN => RST, Q => n_1583, QN => n718);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_20_port, CK 
                           => CLK, RN => RST, Q => n_1584, QN => n717);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_19_port, CK 
                           => CLK, RN => RST, Q => n_1585, QN => n716);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_18_port, CK 
                           => CLK, RN => RST, Q => n_1586, QN => n715);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_17_port, CK 
                           => CLK, RN => RST, Q => n_1587, QN => n714);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_16_port, CK 
                           => CLK, RN => RST, Q => n_1588, QN => n713);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_15_port, CK 
                           => CLK, RN => RST, Q => n_1589, QN => n712);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_14_port, CK 
                           => CLK, RN => RST, Q => n_1590, QN => n711);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_13_port, CK 
                           => CLK, RN => RST, Q => n_1591, QN => n710);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_12_port, CK 
                           => CLK, RN => RST, Q => n_1592, QN => n709);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_11_port, CK 
                           => CLK, RN => RST, Q => n_1593, QN => n708);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_10_port, CK 
                           => CLK, RN => RST, Q => n_1594, QN => n707);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_9_port, CK 
                           => CLK, RN => RST, Q => n_1595, QN => n706);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_8_port, CK 
                           => CLK, RN => RST, Q => n_1596, QN => n705);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_7_port, CK 
                           => CLK, RN => RST, Q => n_1597, QN => n732);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_6_port, CK 
                           => CLK, RN => RST, Q => n_1598, QN => n731);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_5_port, CK 
                           => CLK, RN => RST, Q => n_1599, QN => n730);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_4_port, CK 
                           => CLK, RN => RST, Q => n_1600, QN => n729);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_3_port, CK 
                           => CLK, RN => RST, Q => n_1601, QN => n728);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_2_port, CK 
                           => CLK, RN => RST, Q => n_1602, QN => n734);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_1_port, CK 
                           => CLK, RN => RST, Q => n_1603, QN => n733);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_31_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_32_port, QN => 
                           n_1604);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_30_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_31_port, QN => 
                           n_1605);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_29_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_30_port, QN => 
                           n_1606);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_28_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_29_port, QN => 
                           n_1607);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_27_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_28_port, QN => 
                           n_1608);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_26_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_27_port, QN => 
                           n_1609);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_25_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_26_port, QN => 
                           n_1610);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_24_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_25_port, QN => 
                           n_1611);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_23_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_24_port, QN => 
                           n_1612);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_22_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_23_port, QN => 
                           n_1613);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_21_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_22_port, QN => 
                           n_1614);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_20_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_21_port, QN => 
                           n_1615);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_19_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_20_port, QN => 
                           n_1616);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_18_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_19_port, QN => 
                           n_1617);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_17_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_18_port, QN => 
                           n_1618);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_16_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_17_port, QN => 
                           n_1619);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_15_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_16_port, QN => 
                           n_1620);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_14_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_15_port, QN => 
                           n_1621);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_13_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_14_port, QN => 
                           n_1622);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_12_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_13_port, QN => 
                           n_1623);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_11_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_12_port, QN => 
                           n_1624);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_10_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_11_port, QN => 
                           n_1625);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_9_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_10_port, QN => 
                           n_1626);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_8_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_9_port, QN => 
                           n_1627);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_7_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_8_port, QN => 
                           n_1628);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_6_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_7_port, QN => 
                           n_1629);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_5_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_6_port, QN => 
                           n_1630);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_4_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_5_port, QN => 
                           n_1631);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_3_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_4_port, QN => 
                           n_1632);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_2_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_3_port, QN => 
                           n_1633);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_1_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_2_port, QN => 
                           n_1634);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_0_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_1_port, QN => 
                           n_1635);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_0_port, QN => 
                           n_1636);
   datapath_i_decode_stage_dp_reg_immediate_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_25_port, QN 
                           => n_1637);
   datapath_i_decode_stage_dp_reg_immediate_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_24_port, QN 
                           => n_1638);
   datapath_i_decode_stage_dp_reg_immediate_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_23_port, QN 
                           => n_1639);
   datapath_i_decode_stage_dp_reg_immediate_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_22_port, QN 
                           => n_1640);
   datapath_i_decode_stage_dp_reg_immediate_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_21_port, QN 
                           => n_1641);
   datapath_i_decode_stage_dp_reg_immediate_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_20_port, QN 
                           => n_1642);
   datapath_i_decode_stage_dp_reg_immediate_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_19_port, QN 
                           => n_1643);
   datapath_i_decode_stage_dp_reg_immediate_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_18_port, QN 
                           => n_1644);
   datapath_i_decode_stage_dp_reg_immediate_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_17_port, QN 
                           => n_1645);
   datapath_i_decode_stage_dp_reg_immediate_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_16_port, QN 
                           => n_1646);
   datapath_i_decode_stage_dp_reg_immediate_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_15_port, QN 
                           => n_1647);
   datapath_i_decode_stage_dp_reg_immediate_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_14_port, QN 
                           => n_1648);
   datapath_i_decode_stage_dp_reg_immediate_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_13_port, QN 
                           => n_1649);
   datapath_i_decode_stage_dp_reg_immediate_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_12_port, QN 
                           => n_1650);
   datapath_i_decode_stage_dp_reg_immediate_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_11_port, QN 
                           => n_1651);
   datapath_i_decode_stage_dp_reg_immediate_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_10_port, QN 
                           => n_1652);
   datapath_i_decode_stage_dp_reg_immediate_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_9_port, QN 
                           => n_1653);
   datapath_i_decode_stage_dp_reg_immediate_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_8_port, QN 
                           => n_1654);
   datapath_i_decode_stage_dp_reg_immediate_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_7_port, QN 
                           => n_1655);
   datapath_i_decode_stage_dp_reg_immediate_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_6_port, QN 
                           => n_1656);
   datapath_i_decode_stage_dp_reg_immediate_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_5_port, QN 
                           => n_1657);
   datapath_i_decode_stage_dp_reg_immediate_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_4_port, QN 
                           => n_1658);
   datapath_i_decode_stage_dp_reg_immediate_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_3_port, QN 
                           => n_1659);
   datapath_i_decode_stage_dp_reg_immediate_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_2_port, QN 
                           => n_1660);
   datapath_i_decode_stage_dp_reg_immediate_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_1_port, QN 
                           => n_1661);
   datapath_i_decode_stage_dp_reg_immediate_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_0_port, QN 
                           => n_1662);
   datapath_i_decode_stage_dp_reg_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_31_port, 
                           QN => n764);
   datapath_i_decode_stage_dp_reg_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_30_port, 
                           QN => n763);
   datapath_i_decode_stage_dp_reg_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_29_port, 
                           QN => n762);
   datapath_i_decode_stage_dp_reg_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_28_port, 
                           QN => n761);
   datapath_i_decode_stage_dp_reg_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_27_port, 
                           QN => n760);
   datapath_i_decode_stage_dp_reg_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_26_port, 
                           QN => n759);
   datapath_i_decode_stage_dp_reg_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_25_port, 
                           QN => n758);
   datapath_i_decode_stage_dp_reg_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_24_port, 
                           QN => n_1663);
   datapath_i_decode_stage_dp_reg_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_23_port, 
                           QN => n_1664);
   datapath_i_decode_stage_dp_reg_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_22_port, 
                           QN => n_1665);
   datapath_i_decode_stage_dp_reg_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_21_port, 
                           QN => n_1666);
   datapath_i_decode_stage_dp_reg_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_20_port, 
                           QN => n_1667);
   datapath_i_decode_stage_dp_reg_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_19_port, 
                           QN => n_1668);
   datapath_i_decode_stage_dp_reg_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_18_port, 
                           QN => n_1669);
   datapath_i_decode_stage_dp_reg_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_17_port, 
                           QN => n_1670);
   datapath_i_decode_stage_dp_reg_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_16_port, 
                           QN => n_1671);
   datapath_i_decode_stage_dp_reg_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_15_port, 
                           QN => n_1672);
   datapath_i_decode_stage_dp_reg_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_14_port, 
                           QN => n_1673);
   datapath_i_decode_stage_dp_reg_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_13_port, 
                           QN => n_1674);
   datapath_i_decode_stage_dp_reg_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_12_port, 
                           QN => n_1675);
   datapath_i_decode_stage_dp_reg_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_11_port, 
                           QN => n_1676);
   datapath_i_decode_stage_dp_reg_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_10_port, 
                           QN => n_1677);
   datapath_i_decode_stage_dp_reg_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_9_port, QN 
                           => n_1678);
   datapath_i_decode_stage_dp_reg_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_8_port, QN 
                           => n_1679);
   datapath_i_decode_stage_dp_reg_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_7_port, QN 
                           => n_1680);
   datapath_i_decode_stage_dp_reg_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_6_port, QN 
                           => n_1681);
   datapath_i_decode_stage_dp_reg_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_5_port, QN 
                           => n_1682);
   datapath_i_decode_stage_dp_reg_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_4_port, QN 
                           => n_1683);
   datapath_i_decode_stage_dp_reg_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_3_port, QN 
                           => n_1684);
   datapath_i_decode_stage_dp_reg_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_2_port, QN 
                           => n_1685);
   datapath_i_decode_stage_dp_reg_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_1_port, QN 
                           => n_1686);
   datapath_i_decode_stage_dp_reg_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_0_port, QN 
                           => n_1687);
   datapath_i_decode_stage_dp_reg_a_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_31_port, 
                           QN => n_1688);
   datapath_i_decode_stage_dp_reg_a_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_30_port, 
                           QN => n_1689);
   datapath_i_decode_stage_dp_reg_a_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_29_port, 
                           QN => n_1690);
   datapath_i_decode_stage_dp_reg_a_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_28_port, 
                           QN => n_1691);
   datapath_i_decode_stage_dp_reg_a_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_27_port, 
                           QN => n_1692);
   datapath_i_decode_stage_dp_reg_a_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_26_port, 
                           QN => n_1693);
   datapath_i_decode_stage_dp_reg_a_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_25_port, 
                           QN => n_1694);
   datapath_i_decode_stage_dp_reg_a_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_24_port, 
                           QN => n_1695);
   datapath_i_decode_stage_dp_reg_a_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_23_port, 
                           QN => n_1696);
   datapath_i_decode_stage_dp_reg_a_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_22_port, 
                           QN => n_1697);
   datapath_i_decode_stage_dp_reg_a_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_21_port, 
                           QN => n_1698);
   datapath_i_decode_stage_dp_reg_a_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_20_port, 
                           QN => n_1699);
   datapath_i_decode_stage_dp_reg_a_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_19_port, 
                           QN => n_1700);
   datapath_i_decode_stage_dp_reg_a_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_18_port, 
                           QN => n_1701);
   datapath_i_decode_stage_dp_reg_a_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_17_port, 
                           QN => n_1702);
   datapath_i_decode_stage_dp_reg_a_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_16_port, 
                           QN => n_1703);
   datapath_i_decode_stage_dp_reg_a_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_15_port, 
                           QN => n_1704);
   datapath_i_decode_stage_dp_reg_a_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_14_port, 
                           QN => n_1705);
   datapath_i_decode_stage_dp_reg_a_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_13_port, 
                           QN => n_1706);
   datapath_i_decode_stage_dp_reg_a_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_12_port, 
                           QN => n_1707);
   datapath_i_decode_stage_dp_reg_a_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_11_port, 
                           QN => n_1708);
   datapath_i_decode_stage_dp_reg_a_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_10_port, 
                           QN => n_1709);
   datapath_i_decode_stage_dp_reg_a_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_9_port, QN 
                           => n_1710);
   datapath_i_decode_stage_dp_reg_a_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_8_port, QN 
                           => n_1711);
   datapath_i_decode_stage_dp_reg_a_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_7_port, QN 
                           => n_1712);
   datapath_i_decode_stage_dp_reg_a_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_6_port, QN 
                           => n_1713);
   datapath_i_decode_stage_dp_reg_a_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_5_port, QN 
                           => n_1714);
   datapath_i_decode_stage_dp_reg_a_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_4_port, QN 
                           => n_1715);
   datapath_i_decode_stage_dp_reg_a_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_3_port, QN 
                           => n_1716);
   datapath_i_decode_stage_dp_reg_a_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_2_port, QN 
                           => n_1717);
   datapath_i_decode_stage_dp_reg_a_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_1_port, QN 
                           => n_1718);
   datapath_i_decode_stage_dp_reg_a_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_0_port, QN 
                           => n_1719);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           QN => n_1720);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           QN => n_1721);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           QN => n_1722);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           QN => n_1723);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           QN => n_1724);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_4_port, QN 
                           => n_1725);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_3_port, QN 
                           => n_1726);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_2_port, QN 
                           => n_1727);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_1_port, QN 
                           => n_1728);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_0_port, QN 
                           => n_1729);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n80, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_4_port, QN 
                           => n_1730);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n79, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_3_port, QN 
                           => n_1731);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n78, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_2_port, QN 
                           => n_1732);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n77, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_1_port, QN 
                           => n_1733);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n76, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_0_port, QN 
                           => n_1734);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n69, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_31_port, QN => 
                           n702);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n68, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_30_port, QN => 
                           n_1735);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n67, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_29_port, QN => 
                           n737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n66, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_28_port, QN => 
                           n695);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n65, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_27_port, QN => 
                           n700);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n64, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_26_port, QN => 
                           n693);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n63, CK => CLK, RN => 
                           RST, Q => datapath_i_n9, QN => n_1736);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n62, CK => CLK, RN => 
                           RST, Q => datapath_i_n10, QN => n_1737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n61, CK => CLK, RN => 
                           RST, Q => datapath_i_n11, QN => n_1738);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n60, CK => CLK, RN => 
                           RST, Q => datapath_i_n12, QN => n_1739);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n59, CK => CLK, RN => 
                           RST, Q => datapath_i_n13, QN => n_1740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n58, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_20_port, QN => 
                           n_1741);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n57, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_19_port, QN => 
                           n_1742);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n56, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_18_port, QN => 
                           n697);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n55, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_17_port, QN => 
                           n_1743);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n54, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_16_port, QN => 
                           n_1744);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n53, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_15_port, QN => 
                           n_1745);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n52, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_14_port, QN => 
                           n_1746);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n51, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_13_port, QN => 
                           n740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n50, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_12_port, QN => 
                           n_1747);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n49, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_11_port, QN => 
                           n_1748);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n48, CK => CLK, RN => 
                           RST, Q => datapath_i_n14, QN => n_1749);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n47, CK => CLK, RN => 
                           RST, Q => datapath_i_n15, QN => n_1750);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n46, CK => CLK, RN => 
                           RST, Q => datapath_i_n16, QN => n_1751);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n45, CK => CLK, RN => 
                           RST, Q => datapath_i_n17, QN => n_1752);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n44, CK => CLK, RN => 
                           RST, Q => datapath_i_n18, QN => n_1753);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n43, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_5_port, QN => 
                           n696);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n42, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_4_port, QN => 
                           n698);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n41, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_3_port, QN => 
                           n739);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n40, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_2_port, QN => 
                           n701);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n39, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_1_port, QN => 
                           n690);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n38, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_0_port, QN => 
                           n692);
   datapath_i_fetch_stage_dp_new_program_counter_D_I_31_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n2, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_31_port, QN => n_1754
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_30_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n3, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_30_port, QN => n_1755
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_29_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n4, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_29_port, QN => n_1756
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_28_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n9, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_28_port, QN => n_1757
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_27_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n10, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_27_port, QN => n_1758
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_26_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n11, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_26_port, QN => n_1759
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_25_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n12, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_25_port, QN => n_1760
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_24_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n13, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_24_port, QN => n_1761
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_23_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n14, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_23_port, QN => n_1762
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_22_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n15, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_22_port, QN => n_1763
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_21_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n16, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_21_port, QN => n_1764
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_20_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n17, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_20_port, QN => n_1765
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_19_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n18, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_19_port, QN => n_1766
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_18_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n19, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_18_port, QN => n_1767
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_17_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n20, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_17_port, QN => n_1768
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_16_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n21, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_16_port, QN => n_1769
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_15_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n22, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_15_port, QN => n_1770
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_14_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n23, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_14_port, QN => n_1771
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_13_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n24, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_13_port, QN => n_1772
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_12_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n25, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_12_port, QN => n_1773
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_11_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n26, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_11_port, QN => n_1774
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_10_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n27, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_10_port, QN => n_1775
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_9_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n28, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_9_port, QN => n_1776)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_8_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n29, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_8_port, QN => n_1777)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_7_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n30, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_7_port, QN => n_1778)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_6_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n31, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_6_port, QN => n_1779)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_5_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n32, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_5_port, QN => n_1780)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_4_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n33, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_4_port, QN => n_1781)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_3_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n34, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_3_port, QN => n_1782)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_2_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n35, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_2_port, QN => n_1783)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_1_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n36, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_1_port, QN => n_1784)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n37, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_0_port, QN => n_1785)
                           ;
   datapath_i_fetch_stage_dp_program_counter_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_31_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_31_port, QN => 
                           n_1786);
   datapath_i_fetch_stage_dp_program_counter_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_30_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_30_port, QN => 
                           n_1787);
   datapath_i_fetch_stage_dp_program_counter_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_29_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_29_port, QN => 
                           n753);
   datapath_i_fetch_stage_dp_program_counter_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_28_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_28_port, QN => 
                           n_1788);
   datapath_i_fetch_stage_dp_program_counter_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_27_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_27_port, QN => 
                           n751);
   datapath_i_fetch_stage_dp_program_counter_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_26_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_26_port, QN => 
                           n_1789);
   datapath_i_fetch_stage_dp_program_counter_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_25_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_25_port, QN => 
                           n750);
   datapath_i_fetch_stage_dp_program_counter_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_24_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_24_port, QN => 
                           n_1790);
   datapath_i_fetch_stage_dp_program_counter_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_23_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_23_port, QN => 
                           n749);
   datapath_i_fetch_stage_dp_program_counter_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_22_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_22_port, QN => 
                           n_1791);
   datapath_i_fetch_stage_dp_program_counter_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_21_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_21_port, QN => 
                           n748);
   datapath_i_fetch_stage_dp_program_counter_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_20_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_20_port, QN => 
                           n_1792);
   datapath_i_fetch_stage_dp_program_counter_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_19_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_19_port, QN => 
                           n747);
   datapath_i_fetch_stage_dp_program_counter_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_18_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_18_port, QN => 
                           n_1793);
   datapath_i_fetch_stage_dp_program_counter_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_17_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_17_port, QN => 
                           n746);
   datapath_i_fetch_stage_dp_program_counter_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_16_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_16_port, QN => 
                           n_1794);
   datapath_i_fetch_stage_dp_program_counter_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_15_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_15_port, QN => 
                           n745);
   datapath_i_fetch_stage_dp_program_counter_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_14_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_14_port, QN => 
                           n_1795);
   datapath_i_fetch_stage_dp_program_counter_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_13_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_13_port, QN => 
                           n752);
   datapath_i_fetch_stage_dp_program_counter_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_12_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_12_port, QN => 
                           n_1796);
   datapath_i_fetch_stage_dp_program_counter_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_11_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_11_port, QN => 
                           n744);
   datapath_i_fetch_stage_dp_program_counter_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_10_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_10_port, QN => 
                           n_1797);
   datapath_i_fetch_stage_dp_program_counter_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_9_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_9_port, QN => n743
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_8_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_8_port, QN => 
                           n_1798);
   datapath_i_fetch_stage_dp_program_counter_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_7_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_7_port, QN => n742
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_6_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_6_port, QN => 
                           n_1799);
   datapath_i_fetch_stage_dp_program_counter_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_5_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_5_port, QN => n741
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_4_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_1800);
   datapath_i_fetch_stage_dp_program_counter_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_3_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_1801);
   datapath_i_fetch_stage_dp_program_counter_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_2_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_2_port, QN => 
                           n_1802);
   datapath_i_fetch_stage_dp_program_counter_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N6, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N40_port, QN => 
                           n_1803);
   datapath_i_fetch_stage_dp_program_counter_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N5, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N39_port, QN => 
                           n_1804);
   U305 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(9), ZN => 
                           datapath_i_memory_stage_dp_data_ir_9_port);
   U306 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(8), ZN => 
                           datapath_i_memory_stage_dp_data_ir_8_port);
   U307 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(7), ZN => 
                           datapath_i_memory_stage_dp_data_ir_7_port);
   U308 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(6), ZN => 
                           datapath_i_memory_stage_dp_data_ir_6_port);
   U309 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(5), ZN => 
                           datapath_i_memory_stage_dp_data_ir_5_port);
   U310 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(4), ZN => 
                           datapath_i_memory_stage_dp_data_ir_4_port);
   U311 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(3), ZN => 
                           datapath_i_memory_stage_dp_data_ir_3_port);
   U312 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(31), ZN => 
                           datapath_i_memory_stage_dp_data_ir_31_port);
   U313 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(30), ZN => 
                           datapath_i_memory_stage_dp_data_ir_30_port);
   U314 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(2), ZN => 
                           datapath_i_memory_stage_dp_data_ir_2_port);
   U315 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(29), ZN => 
                           datapath_i_memory_stage_dp_data_ir_29_port);
   U316 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(28), ZN => 
                           datapath_i_memory_stage_dp_data_ir_28_port);
   U317 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(27), ZN => 
                           datapath_i_memory_stage_dp_data_ir_27_port);
   U318 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(26), ZN => 
                           datapath_i_memory_stage_dp_data_ir_26_port);
   U319 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(25), ZN => 
                           datapath_i_memory_stage_dp_data_ir_25_port);
   U320 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(24), ZN => 
                           datapath_i_memory_stage_dp_data_ir_24_port);
   U321 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(23), ZN => 
                           datapath_i_memory_stage_dp_data_ir_23_port);
   U322 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(22), ZN => 
                           datapath_i_memory_stage_dp_data_ir_22_port);
   U323 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(21), ZN => 
                           datapath_i_memory_stage_dp_data_ir_21_port);
   U324 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(20), ZN => 
                           datapath_i_memory_stage_dp_data_ir_20_port);
   U325 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(1), ZN => 
                           datapath_i_memory_stage_dp_data_ir_1_port);
   U326 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(19), ZN => 
                           datapath_i_memory_stage_dp_data_ir_19_port);
   U327 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(18), ZN => 
                           datapath_i_memory_stage_dp_data_ir_18_port);
   U328 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(17), ZN => 
                           datapath_i_memory_stage_dp_data_ir_17_port);
   U329 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(16), ZN => 
                           datapath_i_memory_stage_dp_data_ir_16_port);
   U330 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(15), ZN => 
                           datapath_i_memory_stage_dp_data_ir_15_port);
   U331 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(14), ZN => 
                           datapath_i_memory_stage_dp_data_ir_14_port);
   U332 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(13), ZN => 
                           datapath_i_memory_stage_dp_data_ir_13_port);
   U333 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(12), ZN => 
                           datapath_i_memory_stage_dp_data_ir_12_port);
   U334 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(11), ZN => 
                           datapath_i_memory_stage_dp_data_ir_11_port);
   U335 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(10), ZN => 
                           datapath_i_memory_stage_dp_data_ir_10_port);
   U336 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(0), ZN => 
                           datapath_i_memory_stage_dp_data_ir_0_port);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   cu_i_curr_state_reg_0_inst : DFFS_X1 port map( D => cu_i_n210, CK => CLK, SN
                           => RST, Q => n736, QN => cu_i_n23);
   datapath_i_execute_stage_dp_condition_delay_reg_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_branch_condition_i_0_port, QN => n755);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_0_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, QN => 
                           n_1805);
   cu_i_stall_reg : DFFR_X2 port map( D => cu_i_next_stall, CK => CLK, RN => 
                           RST, Q => n704, QN => cu_i_n4);
   U596 : NOR2_X1 port map( A1 => cu_i_n123, A2 => n736, ZN => n320);
   U597 : NAND2_X1 port map( A1 => n738, A2 => n321, ZN => n447);
   U598 : NAND2_X1 port map( A1 => cu_i_n25, A2 => cu_i_n26, ZN => n321);
   U599 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => 
                           curr_instruction_to_cu_i_29_port, ZN => n318);
   U600 : AND4_X1 port map( A1 => n394, A2 => curr_instruction_to_cu_i_4_port, 
                           A3 => n444, A4 => curr_instruction_to_cu_i_2_port, 
                           ZN => n432);
   U601 : NOR4_X1 port map( A1 => n465, A2 => n702, A3 => n313, A4 => n693, ZN 
                           => cu_i_cmd_word_4_port);
   U602 : OAI21_X2 port map( B1 => n691, B2 => n689, A => n671, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U603 : AOI21_X1 port map( B1 => n573, B2 => n572, A => cu_i_cw3_6_port, ZN 
                           => n574);
   U604 : OAI21_X1 port map( B1 => n448, B2 => n447, A => n699, ZN => 
                           write_rf_i);
   U605 : AOI22_X1 port map( A1 => cu_i_n4, A2 => cu_i_cw1_0_port, B1 => 
                           cu_i_cmd_alu_op_type_0_port, B2 => n704, ZN => n614)
                           ;
   U606 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U607 : NOR2_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, ZN => 
                           n468);
   U608 : NOR2_X1 port map( A1 => n614, A2 => n397, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U609 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           curr_instruction_to_cu_i_28_port, ZN => n319);
   U610 : CLKBUF_X1 port map( A => n685, Z => n689);
   U611 : CLKBUF_X1 port map( A => n415, Z => n470);
   U612 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n755, ZN => n415);
   U613 : AOI21_X1 port map( B1 => n337, B2 => n432, A => n392, ZN => n570);
   U614 : INV_X1 port map( A => n704, ZN => n617);
   U615 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => n695,
                           A3 => n314, A4 => n429, ZN => cu_i_cmd_word_7_port);
   U616 : INV_X1 port map( A => n320, ZN => n465);
   U617 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => n319
                           , ZN => n313);
   U618 : NAND2_X1 port map( A1 => n320, A2 => n318, ZN => n314);
   U619 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => n700
                           , ZN => n429);
   U620 : NOR2_X1 port map( A1 => n314, A2 => n313, ZN => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic);
   U621 : NAND2_X1 port map( A1 => n700, A2 => n693, ZN => n435);
   U622 : INV_X1 port map( A => n435, ZN => n317);
   U623 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n317
                           , ZN => n421);
   U624 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           curr_instruction_to_cu_i_29_port, A3 => n702, ZN => 
                           n428);
   U625 : AOI21_X1 port map( B1 => n421, B2 => n429, A => n428, ZN => n396);
   U626 : NOR4_X1 port map( A1 => n695, A2 => n737, A3 => 
                           curr_instruction_to_cu_i_30_port, A4 => 
                           curr_instruction_to_cu_i_31_port, ZN => n439);
   U627 : INV_X1 port map( A => n439, ZN => n434);
   U628 : NOR2_X1 port map( A1 => n429, A2 => n434, ZN => n438);
   U629 : AND4_X1 port map( A1 => n693, A2 => curr_instruction_to_cu_i_28_port,
                           A3 => curr_instruction_to_cu_i_30_port, A4 => n318, 
                           ZN => n422);
   U630 : NAND3_X1 port map( A1 => n319, A2 => curr_instruction_to_cu_i_29_port
                           , A3 => n702, ZN => n416);
   U631 : AOI21_X1 port map( B1 => n416, B2 => n434, A => 
                           curr_instruction_to_cu_i_26_port, ZN => n315);
   U632 : NOR4_X1 port map( A1 => n396, A2 => n438, A3 => n422, A4 => n315, ZN 
                           => n456);
   U633 : INV_X1 port map( A => n318, ZN => n316);
   U634 : OR3_X1 port map( A1 => n316, A2 => n421, A3 => 
                           curr_instruction_to_cu_i_30_port, ZN => n336);
   U635 : NAND2_X1 port map( A1 => n456, A2 => n336, ZN => n454);
   U636 : AOI211_X1 port map( C1 => n320, C2 => n454, A => cu_i_cmd_word_4_port
                           , B => cu_i_cmd_word_7_port, ZN => n405);
   U637 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           ZN => n568);
   U638 : NAND2_X1 port map( A1 => n405, A2 => n568, ZN => n310);
   U639 : NAND3_X1 port map( A1 => n319, A2 => n318, A3 => n317, ZN => n461);
   U640 : INV_X1 port map( A => n461, ZN => n459);
   U641 : NAND2_X1 port map( A1 => n320, A2 => n459, ZN => n392);
   U642 : INV_X1 port map( A => n392, ZN => n450);
   U643 : OR2_X1 port map( A1 => n310, A2 => n450, ZN => cu_i_N278);
   U644 : OAI22_X1 port map( A1 => n704, A2 => cu_i_cw2_8_port, B1 => 
                           cu_i_cmd_word_4_port, B2 => cu_i_n4, ZN => n309);
   U645 : INV_X1 port map( A => n309, ZN => DRAM_ENABLE_port);
   U646 : INV_X1 port map( A => DRAM_ENABLE_port, ZN => n766);
   U647 : INV_X1 port map( A => cu_i_cmd_word_4_port, ZN => n567);
   U648 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_29_port, A2 => n567,
                           ZN => cu_i_cmd_word_3_port);
   U649 : OAI22_X1 port map( A1 => n704, A2 => cu_i_cw2_7_port, B1 => 
                           cu_i_cmd_word_3_port, B2 => n617, ZN => n406);
   U650 : NAND2_X1 port map( A1 => DRAM_ENABLE_port, A2 => n406, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U651 : CLKBUF_X1 port map( A => datapath_i_memory_stage_dp_n2, Z => n768);
   U652 : NAND4_X1 port map( A1 => cu_i_n25, A2 => cu_i_n26, A3 => n738, A4 => 
                           n694, ZN => cu_i_n145);
   U653 : NAND2_X1 port map( A1 => n447, A2 => cu_i_n145, ZN => n337);
   U654 : NOR2_X1 port map( A1 => n696, A2 => n739, ZN => n394);
   U655 : NOR2_X1 port map( A1 => n692, A2 => n690, ZN => n444);
   U656 : INV_X1 port map( A => n570, ZN => n569);
   U657 : AOI221_X1 port map( B1 => n569, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n570, C2 => 
                           curr_instruction_to_cu_i_11_port, A => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           ZN => n322);
   U658 : INV_X1 port map( A => n322, ZN => datapath_i_decode_stage_dp_n76);
   U659 : AOI221_X1 port map( B1 => n569, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n570, C2 => 
                           curr_instruction_to_cu_i_12_port, A => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           ZN => n323);
   U660 : INV_X1 port map( A => n323, ZN => datapath_i_decode_stage_dp_n77);
   U661 : AOI221_X1 port map( B1 => n569, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n570, C2 => 
                           curr_instruction_to_cu_i_14_port, A => 
                           datapath_i_decode_stage_dp_enable_sign_extension_logic, 
                           ZN => n324);
   U662 : INV_X1 port map( A => n324, ZN => datapath_i_decode_stage_dp_n79);
   U663 : INV_X1 port map( A => n568, ZN => n769);
   U664 : AOI221_X1 port map( B1 => n569, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n570, C2 => 
                           curr_instruction_to_cu_i_15_port, A => n769, ZN => 
                           n325);
   U665 : INV_X1 port map( A => n325, ZN => datapath_i_decode_stage_dp_n80);
   U666 : CLKBUF_X1 port map( A => n468, Z => n412);
   U667 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_11_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_11_port, ZN => 
                           n326);
   U668 : OAI21_X1 port map( B1 => n470, B2 => n709, A => n326, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_11_port);
   U669 : CLKBUF_X1 port map( A => datapath_i_branch_condition_i_0_port, Z => 
                           n413);
   U670 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_9_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_9_port, ZN => n327
                           );
   U671 : OAI21_X1 port map( B1 => n470, B2 => n707, A => n327, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_9_port);
   U672 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_7_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_7_port, ZN => n328
                           );
   U673 : OAI21_X1 port map( B1 => n470, B2 => n705, A => n328, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_7_port);
   U674 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_5_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_5_port, ZN => n329
                           );
   U675 : OAI21_X1 port map( B1 => n470, B2 => n731, A => n329, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_5_port);
   U676 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_4_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_4_port, ZN => n330
                           );
   U677 : OAI21_X1 port map( B1 => n470, B2 => n730, A => n330, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U678 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_3_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_3_port, ZN => n331
                           );
   U679 : OAI21_X1 port map( B1 => n415, B2 => n729, A => n331, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U680 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_2_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_2_port, ZN => n332
                           );
   U681 : OAI21_X1 port map( B1 => n415, B2 => n728, A => n332, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U682 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_6_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_6_port, ZN => n333
                           );
   U683 : OAI21_X1 port map( B1 => n470, B2 => n732, A => n333, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U684 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_8_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_8_port, ZN => n334
                           );
   U685 : OAI21_X1 port map( B1 => n470, B2 => n706, A => n334, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U686 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_10_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_10_port, ZN => 
                           n335);
   U687 : OAI21_X1 port map( B1 => n470, B2 => n708, A => n335, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U688 : OAI21_X1 port map( B1 => n465, B2 => n336, A => n568, ZN => 
                           cu_i_cmd_word_6_port);
   U689 : NOR2_X1 port map( A1 => cu_i_cmd_word_7_port, A2 => 
                           cu_i_cmd_word_6_port, ZN => n464);
   U690 : INV_X1 port map( A => n464, ZN => cu_i_n134);
   U691 : NOR2_X1 port map( A1 => n461, A2 => n337, ZN => n338);
   U692 : AOI21_X1 port map( B1 => n338, B2 => n432, A => n465, ZN => n339);
   U693 : INV_X1 port map( A => n339, ZN => n340);
   U694 : NAND2_X1 port map( A1 => cu_i_n123, A2 => n736, ZN => n463);
   U695 : AOI21_X1 port map( B1 => n340, B2 => n463, A => n704, ZN => 
                           IRAM_ENABLE_port);
   U696 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_11_port, ZN
                           => n341);
   U697 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_9_port, ZN 
                           => n389);
   U698 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_7_port, ZN 
                           => n402);
   U699 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_5_port, ZN 
                           => n399);
   U700 : NAND3_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, A3
                           => datapath_i_new_pc_value_mem_stage_i_2_port, ZN =>
                           n476);
   U701 : NOR2_X1 port map( A1 => n399, A2 => n476, ZN => n483);
   U702 : NAND2_X1 port map( A1 => n483, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, ZN => 
                           n482);
   U703 : NOR2_X1 port map( A1 => n402, A2 => n482, ZN => n489);
   U704 : NAND2_X1 port map( A1 => n489, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, ZN => 
                           n488);
   U705 : NOR2_X1 port map( A1 => n389, A2 => n488, ZN => n495);
   U706 : NAND2_X1 port map( A1 => n495, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, ZN => 
                           n494);
   U707 : AOI221_X1 port map( B1 => cu_i_cw2_4_port, B2 => cu_i_n4, C1 => 
                           cu_i_n134, C2 => n704, A => 
                           datapath_i_branch_condition_i_0_port, ZN => n566);
   U708 : INV_X1 port map( A => n566, ZN => n537);
   U709 : CLKBUF_X1 port map( A => n537, Z => n563);
   U710 : INV_X1 port map( A => n563, ZN => n540);
   U711 : NOR2_X1 port map( A1 => n341, A2 => n494, ZN => n501);
   U712 : AOI211_X1 port map( C1 => n341, C2 => n494, A => n540, B => n501, ZN 
                           => n343);
   U713 : NAND2_X1 port map( A1 => IRAM_ENABLE_port, A2 => IRAM_ADDRESS_2_port,
                           ZN => n471);
   U714 : INV_X1 port map( A => n471, ZN => n473);
   U715 : AND2_X1 port map( A1 => n473, A2 => IRAM_ADDRESS_3_port, ZN => n479);
   U716 : NAND2_X1 port map( A1 => n479, A2 => IRAM_ADDRESS_4_port, ZN => n478)
                           ;
   U717 : NOR2_X1 port map( A1 => n478, A2 => n741, ZN => n485);
   U718 : NAND2_X1 port map( A1 => n485, A2 => IRAM_ADDRESS_6_port, ZN => n484)
                           ;
   U719 : NOR2_X1 port map( A1 => n484, A2 => n742, ZN => n491);
   U720 : NAND2_X1 port map( A1 => n491, A2 => IRAM_ADDRESS_8_port, ZN => n490)
                           ;
   U721 : NOR2_X1 port map( A1 => n490, A2 => n743, ZN => n497);
   U722 : NAND2_X1 port map( A1 => n497, A2 => IRAM_ADDRESS_10_port, ZN => n496
                           );
   U723 : NOR2_X1 port map( A1 => n496, A2 => n744, ZN => n503);
   U724 : AOI211_X1 port map( C1 => n496, C2 => n744, A => n503, B => n563, ZN 
                           => n342);
   U725 : OR2_X1 port map( A1 => n343, A2 => n342, ZN => 
                           datapath_i_fetch_stage_dp_n26);
   U726 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_13_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_13_port, ZN => 
                           n344);
   U727 : OAI21_X1 port map( B1 => n470, B2 => n711, A => n344, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_13_port);
   U728 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_12_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_12_port, ZN => 
                           n345);
   U729 : OAI21_X1 port map( B1 => n470, B2 => n710, A => n345, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U730 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_13_port, ZN
                           => n346);
   U731 : NAND2_X1 port map( A1 => n501, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, ZN => 
                           n500);
   U732 : INV_X1 port map( A => n537, ZN => n557);
   U733 : NOR2_X1 port map( A1 => n346, A2 => n500, ZN => n507);
   U734 : AOI211_X1 port map( C1 => n346, C2 => n500, A => n557, B => n507, ZN 
                           => n348);
   U735 : NAND2_X1 port map( A1 => n503, A2 => IRAM_ADDRESS_12_port, ZN => n502
                           );
   U736 : NOR2_X1 port map( A1 => n502, A2 => n752, ZN => n509);
   U737 : AOI211_X1 port map( C1 => n502, C2 => n752, A => n509, B => n537, ZN 
                           => n347);
   U738 : OR2_X1 port map( A1 => n348, A2 => n347, ZN => 
                           datapath_i_fetch_stage_dp_n24);
   U739 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_15_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_15_port, ZN => 
                           n349);
   U740 : OAI21_X1 port map( B1 => n415, B2 => n713, A => n349, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_15_port);
   U741 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_14_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_14_port, ZN => 
                           n350);
   U742 : OAI21_X1 port map( B1 => n470, B2 => n712, A => n350, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U743 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_15_port, ZN
                           => n351);
   U744 : NAND2_X1 port map( A1 => n507, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, ZN => 
                           n506);
   U745 : NOR2_X1 port map( A1 => n351, A2 => n506, ZN => n513);
   U746 : AOI211_X1 port map( C1 => n351, C2 => n506, A => n540, B => n513, ZN 
                           => n353);
   U747 : NAND2_X1 port map( A1 => n509, A2 => IRAM_ADDRESS_14_port, ZN => n508
                           );
   U748 : NOR2_X1 port map( A1 => n508, A2 => n745, ZN => n515);
   U749 : AOI211_X1 port map( C1 => n508, C2 => n745, A => n515, B => n537, ZN 
                           => n352);
   U750 : OR2_X1 port map( A1 => n353, A2 => n352, ZN => 
                           datapath_i_fetch_stage_dp_n22);
   U751 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_17_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_17_port, ZN => 
                           n354);
   U752 : OAI21_X1 port map( B1 => n415, B2 => n715, A => n354, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_17_port);
   U753 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_16_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_16_port, ZN => 
                           n355);
   U754 : OAI21_X1 port map( B1 => n470, B2 => n714, A => n355, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U755 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_17_port, ZN
                           => n356);
   U756 : NAND2_X1 port map( A1 => n513, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, ZN => 
                           n512);
   U757 : NOR2_X1 port map( A1 => n356, A2 => n512, ZN => n519);
   U758 : AOI211_X1 port map( C1 => n356, C2 => n512, A => n557, B => n519, ZN 
                           => n358);
   U759 : NAND2_X1 port map( A1 => n515, A2 => IRAM_ADDRESS_16_port, ZN => n514
                           );
   U760 : NOR2_X1 port map( A1 => n514, A2 => n746, ZN => n521);
   U761 : AOI211_X1 port map( C1 => n514, C2 => n746, A => n521, B => n537, ZN 
                           => n357);
   U762 : OR2_X1 port map( A1 => n358, A2 => n357, ZN => 
                           datapath_i_fetch_stage_dp_n20);
   U763 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_19_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_19_port, ZN => 
                           n359);
   U764 : OAI21_X1 port map( B1 => n415, B2 => n717, A => n359, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_19_port);
   U765 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_18_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_18_port, ZN => 
                           n360);
   U766 : OAI21_X1 port map( B1 => n470, B2 => n716, A => n360, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U767 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_19_port, ZN
                           => n361);
   U768 : NAND2_X1 port map( A1 => n519, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, ZN => 
                           n518);
   U769 : NOR2_X1 port map( A1 => n361, A2 => n518, ZN => n525);
   U770 : AOI211_X1 port map( C1 => n361, C2 => n518, A => n557, B => n525, ZN 
                           => n363);
   U771 : NAND2_X1 port map( A1 => n521, A2 => IRAM_ADDRESS_18_port, ZN => n520
                           );
   U772 : NOR2_X1 port map( A1 => n520, A2 => n747, ZN => n527);
   U773 : AOI211_X1 port map( C1 => n520, C2 => n747, A => n527, B => n563, ZN 
                           => n362);
   U774 : OR2_X1 port map( A1 => n363, A2 => n362, ZN => 
                           datapath_i_fetch_stage_dp_n18);
   U775 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_21_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_21_port, ZN => 
                           n364);
   U776 : OAI21_X1 port map( B1 => n415, B2 => n719, A => n364, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_21_port);
   U777 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_20_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_20_port, ZN => 
                           n365);
   U778 : OAI21_X1 port map( B1 => n470, B2 => n718, A => n365, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U779 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_21_port, ZN
                           => n366);
   U780 : NAND2_X1 port map( A1 => n525, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, ZN => 
                           n524);
   U781 : NOR2_X1 port map( A1 => n366, A2 => n524, ZN => n531);
   U782 : AOI211_X1 port map( C1 => n366, C2 => n524, A => n557, B => n531, ZN 
                           => n368);
   U783 : NAND2_X1 port map( A1 => n527, A2 => IRAM_ADDRESS_20_port, ZN => n526
                           );
   U784 : NOR2_X1 port map( A1 => n526, A2 => n748, ZN => n533);
   U785 : AOI211_X1 port map( C1 => n526, C2 => n748, A => n533, B => n537, ZN 
                           => n367);
   U786 : OR2_X1 port map( A1 => n368, A2 => n367, ZN => 
                           datapath_i_fetch_stage_dp_n16);
   U787 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_23_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_23_port, ZN => 
                           n369);
   U788 : OAI21_X1 port map( B1 => n415, B2 => n721, A => n369, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_23_port);
   U789 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_22_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_22_port, ZN => 
                           n370);
   U790 : OAI21_X1 port map( B1 => n470, B2 => n720, A => n370, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U791 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_23_port, ZN
                           => n371);
   U792 : NAND2_X1 port map( A1 => n531, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, ZN => 
                           n530);
   U793 : NOR2_X1 port map( A1 => n371, A2 => n530, ZN => n538);
   U794 : AOI211_X1 port map( C1 => n371, C2 => n530, A => n557, B => n538, ZN 
                           => n373);
   U795 : NAND2_X1 port map( A1 => n533, A2 => IRAM_ADDRESS_22_port, ZN => n532
                           );
   U796 : NOR2_X1 port map( A1 => n532, A2 => n749, ZN => n541);
   U797 : AOI211_X1 port map( C1 => n532, C2 => n749, A => n541, B => n537, ZN 
                           => n372);
   U798 : OR2_X1 port map( A1 => n373, A2 => n372, ZN => 
                           datapath_i_fetch_stage_dp_n14);
   U799 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_25_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_25_port, ZN => 
                           n374);
   U800 : OAI21_X1 port map( B1 => n415, B2 => n723, A => n374, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_25_port);
   U801 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_24_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_24_port, ZN => 
                           n375);
   U802 : OAI21_X1 port map( B1 => n415, B2 => n722, A => n375, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U803 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_25_port, ZN
                           => n376);
   U804 : NAND2_X1 port map( A1 => n538, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, ZN => 
                           n536);
   U805 : NOR2_X1 port map( A1 => n376, A2 => n536, ZN => n545);
   U806 : AOI211_X1 port map( C1 => n376, C2 => n536, A => n557, B => n545, ZN 
                           => n378);
   U807 : NAND2_X1 port map( A1 => n541, A2 => IRAM_ADDRESS_24_port, ZN => n539
                           );
   U808 : NOR2_X1 port map( A1 => n539, A2 => n750, ZN => n547);
   U809 : AOI211_X1 port map( C1 => n539, C2 => n750, A => n547, B => n537, ZN 
                           => n377);
   U810 : OR2_X1 port map( A1 => n378, A2 => n377, ZN => 
                           datapath_i_fetch_stage_dp_n12);
   U811 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_27_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_27_port, ZN => 
                           n379);
   U812 : OAI21_X1 port map( B1 => n415, B2 => n724, A => n379, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_27_port);
   U813 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_26_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_26_port, ZN => 
                           n380);
   U814 : OAI21_X1 port map( B1 => n415, B2 => n691, A => n380, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U815 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_27_port, ZN
                           => n381);
   U816 : NAND2_X1 port map( A1 => n545, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, ZN => 
                           n544);
   U817 : NOR2_X1 port map( A1 => n381, A2 => n544, ZN => n551);
   U818 : AOI211_X1 port map( C1 => n381, C2 => n544, A => n557, B => n551, ZN 
                           => n383);
   U819 : NAND2_X1 port map( A1 => n547, A2 => IRAM_ADDRESS_26_port, ZN => n546
                           );
   U820 : NOR2_X1 port map( A1 => n546, A2 => n751, ZN => n553);
   U821 : AOI211_X1 port map( C1 => n546, C2 => n751, A => n553, B => n563, ZN 
                           => n382);
   U822 : OR2_X1 port map( A1 => n383, A2 => n382, ZN => 
                           datapath_i_fetch_stage_dp_n10);
   U823 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_29_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_29_port, ZN => 
                           n384);
   U824 : OAI21_X1 port map( B1 => n415, B2 => n726, A => n384, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_29_port);
   U825 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_28_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_28_port, ZN => 
                           n385);
   U826 : OAI21_X1 port map( B1 => n415, B2 => n725, A => n385, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U827 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_29_port, ZN
                           => n386);
   U828 : NAND2_X1 port map( A1 => n551, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, ZN => 
                           n550);
   U829 : NOR2_X1 port map( A1 => n386, A2 => n550, ZN => n556);
   U830 : AOI211_X1 port map( C1 => n386, C2 => n550, A => n540, B => n556, ZN 
                           => n388);
   U831 : NAND2_X1 port map( A1 => n553, A2 => IRAM_ADDRESS_28_port, ZN => n552
                           );
   U832 : NOR2_X1 port map( A1 => n552, A2 => n753, ZN => n558);
   U833 : AOI211_X1 port map( C1 => n552, C2 => n753, A => n558, B => n537, ZN 
                           => n387);
   U834 : OR2_X1 port map( A1 => n388, A2 => n387, ZN => 
                           datapath_i_fetch_stage_dp_n4);
   U835 : AOI211_X1 port map( C1 => n389, C2 => n488, A => n540, B => n495, ZN 
                           => n391);
   U836 : AOI211_X1 port map( C1 => n490, C2 => n743, A => n497, B => n563, ZN 
                           => n390);
   U837 : OR2_X1 port map( A1 => n391, A2 => n390, ZN => 
                           datapath_i_fetch_stage_dp_n28);
   U838 : OAI222_X1 port map( A1 => n693, A2 => n568, B1 => n392, B2 => n432, 
                           C1 => n465, C2 => n456, ZN => n311);
   U839 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n311, ZN => 
                           cu_i_cmd_word_1_port);
   U840 : OAI22_X1 port map( A1 => n704, A2 => cu_i_cw2_6_port, B1 => 
                           cu_i_cw3_6_port, B2 => n617, ZN => n393);
   U841 : INV_X1 port map( A => n393, ZN => cu_i_n132);
   U842 : NAND3_X1 port map( A1 => n394, A2 => n698, A3 => n690, ZN => n425);
   U843 : AOI211_X1 port map( C1 => n692, C2 => n701, A => n461, B => n425, ZN 
                           => n395);
   U844 : OR2_X1 port map( A1 => n396, A2 => n395, ZN => cu_i_N267);
   U845 : CLKBUF_X1 port map( A => n310, Z => n765);
   U846 : AOI22_X1 port map( A1 => cu_i_n4, A2 => cu_i_cw1_1_port, B1 => 
                           cu_i_cmd_alu_op_type_1_port, B2 => n704, ZN => n616)
                           ;
   U847 : AOI22_X1 port map( A1 => n617, A2 => cu_i_cw1_2_port, B1 => 
                           cu_i_cmd_alu_op_type_2_port, B2 => n704, ZN => n633)
                           ;
   U848 : AOI22_X1 port map( A1 => cu_i_n4, A2 => cu_i_cw1_3_port, B1 => 
                           cu_i_cmd_alu_op_type_3_port, B2 => n704, ZN => n613)
                           ;
   U849 : AOI21_X1 port map( B1 => n616, B2 => n633, A => n613, ZN => n397);
   U850 : INV_X1 port map( A => n613, ZN => n632);
   U851 : OAI211_X1 port map( C1 => n614, C2 => n616, A => n632, B => n633, ZN 
                           => n398);
   U852 : INV_X1 port map( A => n398, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_3_port);
   U853 : AOI211_X1 port map( C1 => n399, C2 => n476, A => n540, B => n483, ZN 
                           => n401);
   U854 : AOI211_X1 port map( C1 => n478, C2 => n741, A => n485, B => n537, ZN 
                           => n400);
   U855 : OR2_X1 port map( A1 => n401, A2 => n400, ZN => 
                           datapath_i_fetch_stage_dp_n32);
   U856 : AOI211_X1 port map( C1 => n402, C2 => n482, A => n540, B => n489, ZN 
                           => n404);
   U857 : AOI211_X1 port map( C1 => n484, C2 => n742, A => n491, B => n537, ZN 
                           => n403);
   U858 : OR2_X1 port map( A1 => n404, A2 => n403, ZN => 
                           datapath_i_fetch_stage_dp_n30);
   U859 : NAND2_X1 port map( A1 => n405, A2 => n569, ZN => enable_rf_i);
   U860 : NAND2_X1 port map( A1 => n450, A2 => n432, ZN => n448);
   U861 : AND2_X1 port map( A1 => n310, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U862 : INV_X1 port map( A => n406, ZN => DRAM_READNOTWRITE);
   U863 : AOI22_X1 port map( A1 => n617, A2 => cu_i_cw1_13_port, B1 => n310, B2
                           => n704, ZN => n407);
   U864 : INV_X1 port map( A => n407, ZN => n647);
   U865 : CLKBUF_X1 port map( A => n647, Z => n648);
   U866 : MUX2_X1 port map( A => datapath_i_val_b_i_0_port, B => 
                           datapath_i_val_immediate_i_0_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U867 : MUX2_X1 port map( A => datapath_i_val_b_i_2_port, B => 
                           datapath_i_val_immediate_i_2_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U868 : NOR2_X1 port map( A1 => n694, A2 => n448, ZN => cu_i_N273);
   U869 : INV_X1 port map( A => n448, ZN => n573);
   U870 : AOI221_X1 port map( B1 => cu_i_n25, B2 => n573, C1 => cu_i_n26, C2 =>
                           n573, A => cu_i_N273, ZN => n408);
   U871 : INV_X1 port map( A => n408, ZN => n410);
   U872 : NAND3_X1 port map( A1 => n573, A2 => n735, A3 => n694, ZN => n446);
   U873 : NOR2_X1 port map( A1 => cu_i_n25, A2 => n446, ZN => n409);
   U874 : MUX2_X1 port map( A => n410, B => n409, S => cu_i_n124, Z => 
                           cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U876 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_31_port, B1 => 
                           datapath_i_new_pc_value_decode_31_port, B2 => n468, 
                           ZN => n411);
   U877 : OAI21_X1 port map( B1 => n703, B2 => n415, A => n411, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_31_port);
   U878 : AOI22_X1 port map( A1 => n413, A2 => 
                           datapath_i_alu_output_val_i_30_port, B1 => n412, B2 
                           => datapath_i_new_pc_value_decode_30_port, ZN => 
                           n414);
   U879 : OAI21_X1 port map( B1 => n415, B2 => n727, A => n414, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   U880 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => n700,
                           A3 => n416, ZN => n449);
   U881 : AOI21_X1 port map( B1 => n439, B2 => n693, A => n449, ZN => n420);
   U882 : OAI221_X1 port map( B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           curr_instruction_to_cu_i_5_port, C1 => n690, C2 => 
                           n739, A => n698, ZN => n417);
   U883 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_4_port, A3 => n696, ZN => 
                           n437);
   U884 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_1_port, A2 => n437,
                           ZN => n452);
   U885 : AOI221_X1 port map( B1 => n417, B2 => n452, C1 => n701, C2 => n452, A
                           => curr_instruction_to_cu_i_0_port, ZN => n418);
   U886 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => n422
                           , B1 => n459, B2 => n418, ZN => n419);
   U887 : OAI211_X1 port map( C1 => n421, C2 => n428, A => n420, B => n419, ZN 
                           => cu_i_N264);
   U888 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_4_port, ZN => n424);
   U889 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => 
                           curr_instruction_to_cu_i_5_port, A3 => n461, A4 => 
                           n701, ZN => n423);
   U890 : AOI21_X1 port map( B1 => n424, B2 => n423, A => n422, ZN => n442);
   U891 : NOR2_X1 port map( A1 => n692, A2 => n425, ZN => n427);
   U892 : AND3_X1 port map( A1 => n437, A2 => n692, A3 => n690, ZN => n426);
   U893 : MUX2_X1 port map( A => n427, B => n426, S => 
                           curr_instruction_to_cu_i_2_port, Z => n431);
   U894 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n429,
                           A3 => n428, ZN => n430);
   U895 : AOI221_X1 port map( B1 => n432, B2 => n459, C1 => n431, C2 => n459, A
                           => n430, ZN => n433);
   U896 : OAI211_X1 port map( C1 => n435, C2 => n434, A => n442, B => n433, ZN 
                           => cu_i_N265);
   U897 : NAND2_X1 port map( A1 => n692, A2 => n690, ZN => n436);
   U898 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => n459,
                           A3 => n437, A4 => n436, ZN => n443);
   U899 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => n700,
                           ZN => n440);
   U900 : AOI21_X1 port map( B1 => n440, B2 => n439, A => n438, ZN => n441);
   U901 : OAI211_X1 port map( C1 => n444, C2 => n443, A => n442, B => n441, ZN 
                           => cu_i_N266);
   U902 : NAND2_X1 port map( A1 => n704, A2 => n448, ZN => cu_i_N274);
   U903 : AOI221_X1 port map( B1 => cu_i_n125, B2 => cu_i_n26, C1 => n694, C2 
                           => n735, A => n448, ZN => cu_i_N275);
   U904 : OAI21_X1 port map( B1 => cu_i_n26, B2 => cu_i_n125, A => n573, ZN => 
                           n445);
   U905 : AOI22_X1 port map( A1 => cu_i_n25, A2 => n446, B1 => n445, B2 => n754
                           , ZN => cu_i_N276);
   U906 : INV_X1 port map( A => n447, ZN => n572);
   U907 : AOI211_X1 port map( C1 => n704, C2 => cu_i_n145, A => n572, B => n448
                           , ZN => cu_i_N279);
   U908 : INV_X1 port map( A => n449, ZN => n453);
   U909 : NAND3_X1 port map( A1 => n450, A2 => n692, A3 => n701, ZN => n451);
   U910 : OAI22_X1 port map( A1 => n465, A2 => n453, B1 => n452, B2 => n451, ZN
                           => cu_i_cmd_word_8_port);
   U911 : MUX2_X1 port map( A => cu_i_cmd_word_8_port, B => cu_i_cw1_12_port, S
                           => cu_i_n4, Z => alu_cin_i);
   U912 : NOR2_X1 port map( A1 => cu_i_cw1_4_port, A2 => n704, ZN => n649);
   U913 : AOI21_X1 port map( B1 => n704, B2 => n756, A => n649, ZN => 
                           cu_i_cw1_i_4_port);
   U914 : MUX2_X1 port map( A => cu_i_cw2_7_port, B => cu_i_cw1_7_port, S => 
                           cu_i_n4, Z => cu_i_cw1_i_7_port);
   U915 : MUX2_X1 port map( A => cu_i_cw2_8_port, B => cu_i_cw1_8_port, S => 
                           n617, Z => cu_i_cw1_i_8_port);
   U916 : INV_X1 port map( A => n454, ZN => n462);
   U917 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_14_port, A2 => 
                           curr_instruction_to_cu_i_15_port, A3 => 
                           curr_instruction_to_cu_i_11_port, A4 => 
                           curr_instruction_to_cu_i_12_port, ZN => n455);
   U918 : NAND2_X1 port map( A1 => n455, A2 => n740, ZN => n460);
   U919 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_19_port, A2 => 
                           curr_instruction_to_cu_i_20_port, A3 => 
                           curr_instruction_to_cu_i_16_port, A4 => 
                           curr_instruction_to_cu_i_17_port, ZN => n457);
   U920 : AOI21_X1 port map( B1 => n457, B2 => n697, A => n456, ZN => n458);
   U921 : AOI221_X1 port map( B1 => n462, B2 => n461, C1 => n460, C2 => n459, A
                           => n458, ZN => n466);
   U922 : OAI211_X1 port map( C1 => n466, C2 => n465, A => n464, B => n463, ZN 
                           => cu_i_n209);
   U923 : NOR2_X1 port map( A1 => cu_i_n123, A2 => cu_i_n23, ZN => cu_i_n210);
   U924 : AOI22_X1 port map( A1 => cu_i_n4, A2 => n757, B1 => n699, B2 => n704,
                           ZN => cu_i_n131);
   U925 : MUX2_X1 port map( A => cu_i_cw2_6_port, B => cu_i_cw1_6_port, S => 
                           n617, Z => cu_i_n127);
   U926 : MUX2_X1 port map( A => cu_i_cw2_5_port, B => cu_i_cw1_5_port, S => 
                           n617, Z => cu_i_n126);
   U927 : MUX2_X1 port map( A => curr_instruction_to_cu_i_31_port, B => 
                           IRAM_DATA(31), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n69);
   U928 : MUX2_X1 port map( A => curr_instruction_to_cu_i_30_port, B => 
                           IRAM_DATA(30), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n68);
   U929 : MUX2_X1 port map( A => curr_instruction_to_cu_i_29_port, B => 
                           IRAM_DATA(29), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n67);
   U930 : MUX2_X1 port map( A => curr_instruction_to_cu_i_28_port, B => 
                           IRAM_DATA(28), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n66);
   U931 : MUX2_X1 port map( A => curr_instruction_to_cu_i_27_port, B => 
                           IRAM_DATA(27), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n65);
   U932 : MUX2_X1 port map( A => curr_instruction_to_cu_i_26_port, B => 
                           IRAM_DATA(26), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n64);
   U933 : MUX2_X1 port map( A => datapath_i_n9, B => IRAM_DATA(25), S => 
                           cu_i_n4, Z => datapath_i_fetch_stage_dp_n63);
   U934 : MUX2_X1 port map( A => datapath_i_n10, B => IRAM_DATA(24), S => n617,
                           Z => datapath_i_fetch_stage_dp_n62);
   U935 : MUX2_X1 port map( A => datapath_i_n11, B => IRAM_DATA(23), S => 
                           cu_i_n4, Z => datapath_i_fetch_stage_dp_n61);
   U936 : MUX2_X1 port map( A => datapath_i_n12, B => IRAM_DATA(22), S => 
                           cu_i_n4, Z => datapath_i_fetch_stage_dp_n60);
   U937 : MUX2_X1 port map( A => datapath_i_n13, B => IRAM_DATA(21), S => 
                           cu_i_n4, Z => datapath_i_fetch_stage_dp_n59);
   U938 : MUX2_X1 port map( A => curr_instruction_to_cu_i_20_port, B => 
                           IRAM_DATA(20), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n58);
   U939 : MUX2_X1 port map( A => curr_instruction_to_cu_i_19_port, B => 
                           IRAM_DATA(19), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n57);
   U940 : MUX2_X1 port map( A => curr_instruction_to_cu_i_18_port, B => 
                           IRAM_DATA(18), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n56);
   U941 : MUX2_X1 port map( A => curr_instruction_to_cu_i_17_port, B => 
                           IRAM_DATA(17), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n55);
   U942 : MUX2_X1 port map( A => curr_instruction_to_cu_i_16_port, B => 
                           IRAM_DATA(16), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n54);
   U943 : MUX2_X1 port map( A => curr_instruction_to_cu_i_15_port, B => 
                           IRAM_DATA(15), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n53);
   U944 : MUX2_X1 port map( A => curr_instruction_to_cu_i_14_port, B => 
                           IRAM_DATA(14), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n52);
   U945 : MUX2_X1 port map( A => curr_instruction_to_cu_i_13_port, B => 
                           IRAM_DATA(13), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n51);
   U946 : MUX2_X1 port map( A => curr_instruction_to_cu_i_12_port, B => 
                           IRAM_DATA(12), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n50);
   U947 : MUX2_X1 port map( A => curr_instruction_to_cu_i_11_port, B => 
                           IRAM_DATA(11), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n49);
   U948 : MUX2_X1 port map( A => datapath_i_n14, B => IRAM_DATA(10), S => n617,
                           Z => datapath_i_fetch_stage_dp_n48);
   U949 : MUX2_X1 port map( A => datapath_i_n15, B => IRAM_DATA(9), S => 
                           cu_i_n4, Z => datapath_i_fetch_stage_dp_n47);
   U950 : MUX2_X1 port map( A => datapath_i_n16, B => IRAM_DATA(8), S => n617, 
                           Z => datapath_i_fetch_stage_dp_n46);
   U951 : MUX2_X1 port map( A => datapath_i_n17, B => IRAM_DATA(7), S => 
                           cu_i_n4, Z => datapath_i_fetch_stage_dp_n45);
   U952 : MUX2_X1 port map( A => datapath_i_n18, B => IRAM_DATA(6), S => n617, 
                           Z => datapath_i_fetch_stage_dp_n44);
   U953 : MUX2_X1 port map( A => curr_instruction_to_cu_i_5_port, B => 
                           IRAM_DATA(5), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n43);
   U954 : MUX2_X1 port map( A => curr_instruction_to_cu_i_4_port, B => 
                           IRAM_DATA(4), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n42);
   U955 : MUX2_X1 port map( A => curr_instruction_to_cu_i_3_port, B => 
                           IRAM_DATA(3), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n41);
   U956 : MUX2_X1 port map( A => curr_instruction_to_cu_i_2_port, B => 
                           IRAM_DATA(2), S => n617, Z => 
                           datapath_i_fetch_stage_dp_n40);
   U957 : MUX2_X1 port map( A => curr_instruction_to_cu_i_1_port, B => 
                           IRAM_DATA(1), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n39);
   U958 : MUX2_X1 port map( A => curr_instruction_to_cu_i_0_port, B => 
                           IRAM_DATA(0), S => cu_i_n4, Z => 
                           datapath_i_fetch_stage_dp_n38);
   U959 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_0_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_0_port, ZN => n467
                           );
   U960 : OAI21_X1 port map( B1 => n470, B2 => n733, A => n467, ZN => 
                           datapath_i_fetch_stage_dp_N5);
   U961 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N5, B => 
                           datapath_i_fetch_stage_dp_N39_port, S => n566, Z => 
                           datapath_i_fetch_stage_dp_n37);
   U962 : AOI22_X1 port map( A1 => datapath_i_branch_condition_i_0_port, A2 => 
                           datapath_i_alu_output_val_i_1_port, B1 => n468, B2 
                           => datapath_i_new_pc_value_decode_1_port, ZN => n469
                           );
   U963 : OAI21_X1 port map( B1 => n470, B2 => n734, A => n469, ZN => 
                           datapath_i_fetch_stage_dp_N6);
   U964 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N6, B => 
                           datapath_i_fetch_stage_dp_N40_port, S => n566, Z => 
                           datapath_i_fetch_stage_dp_n36);
   U965 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port,
                           A => n471, ZN => n472);
   U966 : AOI22_X1 port map( A1 => n566, A2 => n472, B1 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B2 => 
                           n537, ZN => datapath_i_fetch_stage_dp_n35);
   U967 : OAI21_X1 port map( B1 => n473, B2 => IRAM_ADDRESS_3_port, A => n566, 
                           ZN => n475);
   U968 : AND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_3_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_2_port, ZN
                           => n477);
   U969 : OAI21_X1 port map( B1 => datapath_i_new_pc_value_mem_stage_i_3_port, 
                           B2 => datapath_i_new_pc_value_mem_stage_i_2_port, A 
                           => n537, ZN => n474);
   U970 : OAI22_X1 port map( A1 => n479, A2 => n475, B1 => n477, B2 => n474, ZN
                           => datapath_i_fetch_stage_dp_n34);
   U971 : OAI211_X1 port map( C1 => n477, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n563, B => n476, ZN => n481);
   U972 : OAI211_X1 port map( C1 => n479, C2 => IRAM_ADDRESS_4_port, A => n557,
                           B => n478, ZN => n480);
   U973 : NAND2_X1 port map( A1 => n481, A2 => n480, ZN => 
                           datapath_i_fetch_stage_dp_n33);
   U974 : OAI211_X1 port map( C1 => n483, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, A => 
                           n537, B => n482, ZN => n487);
   U975 : OAI211_X1 port map( C1 => n485, C2 => IRAM_ADDRESS_6_port, A => n557,
                           B => n484, ZN => n486);
   U976 : NAND2_X1 port map( A1 => n487, A2 => n486, ZN => 
                           datapath_i_fetch_stage_dp_n31);
   U977 : OAI211_X1 port map( C1 => n489, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, A => 
                           n563, B => n488, ZN => n493);
   U978 : OAI211_X1 port map( C1 => n491, C2 => IRAM_ADDRESS_8_port, A => n540,
                           B => n490, ZN => n492);
   U979 : NAND2_X1 port map( A1 => n493, A2 => n492, ZN => 
                           datapath_i_fetch_stage_dp_n29);
   U980 : OAI211_X1 port map( C1 => n495, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, A => 
                           n537, B => n494, ZN => n499);
   U981 : OAI211_X1 port map( C1 => n497, C2 => IRAM_ADDRESS_10_port, A => n540
                           , B => n496, ZN => n498);
   U982 : NAND2_X1 port map( A1 => n499, A2 => n498, ZN => 
                           datapath_i_fetch_stage_dp_n27);
   U983 : OAI211_X1 port map( C1 => n501, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, A => 
                           n563, B => n500, ZN => n505);
   U984 : OAI211_X1 port map( C1 => n503, C2 => IRAM_ADDRESS_12_port, A => n540
                           , B => n502, ZN => n504);
   U985 : NAND2_X1 port map( A1 => n505, A2 => n504, ZN => 
                           datapath_i_fetch_stage_dp_n25);
   U986 : OAI211_X1 port map( C1 => n507, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, A => 
                           n563, B => n506, ZN => n511);
   U987 : OAI211_X1 port map( C1 => n509, C2 => IRAM_ADDRESS_14_port, A => n540
                           , B => n508, ZN => n510);
   U988 : NAND2_X1 port map( A1 => n511, A2 => n510, ZN => 
                           datapath_i_fetch_stage_dp_n23);
   U989 : OAI211_X1 port map( C1 => n513, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, A => 
                           n563, B => n512, ZN => n517);
   U990 : OAI211_X1 port map( C1 => n515, C2 => IRAM_ADDRESS_16_port, A => n540
                           , B => n514, ZN => n516);
   U991 : NAND2_X1 port map( A1 => n517, A2 => n516, ZN => 
                           datapath_i_fetch_stage_dp_n21);
   U992 : OAI211_X1 port map( C1 => n519, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, A => 
                           n563, B => n518, ZN => n523);
   U993 : OAI211_X1 port map( C1 => n521, C2 => IRAM_ADDRESS_18_port, A => n540
                           , B => n520, ZN => n522);
   U994 : NAND2_X1 port map( A1 => n523, A2 => n522, ZN => 
                           datapath_i_fetch_stage_dp_n19);
   U995 : OAI211_X1 port map( C1 => n525, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, A => 
                           n563, B => n524, ZN => n529);
   U996 : OAI211_X1 port map( C1 => n527, C2 => IRAM_ADDRESS_20_port, A => n540
                           , B => n526, ZN => n528);
   U997 : NAND2_X1 port map( A1 => n529, A2 => n528, ZN => 
                           datapath_i_fetch_stage_dp_n17);
   U998 : OAI211_X1 port map( C1 => n531, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, A => 
                           n563, B => n530, ZN => n535);
   U999 : OAI211_X1 port map( C1 => n533, C2 => IRAM_ADDRESS_22_port, A => n557
                           , B => n532, ZN => n534);
   U1000 : NAND2_X1 port map( A1 => n535, A2 => n534, ZN => 
                           datapath_i_fetch_stage_dp_n15);
   U1001 : OAI211_X1 port map( C1 => n538, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, A => 
                           n537, B => n536, ZN => n543);
   U1002 : OAI211_X1 port map( C1 => n541, C2 => IRAM_ADDRESS_24_port, A => 
                           n540, B => n539, ZN => n542);
   U1003 : NAND2_X1 port map( A1 => n543, A2 => n542, ZN => 
                           datapath_i_fetch_stage_dp_n13);
   U1004 : OAI211_X1 port map( C1 => n545, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, A => 
                           n563, B => n544, ZN => n549);
   U1005 : OAI211_X1 port map( C1 => n547, C2 => IRAM_ADDRESS_26_port, A => 
                           n557, B => n546, ZN => n548);
   U1006 : NAND2_X1 port map( A1 => n549, A2 => n548, ZN => 
                           datapath_i_fetch_stage_dp_n11);
   U1007 : OAI211_X1 port map( C1 => n551, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, A => 
                           n563, B => n550, ZN => n555);
   U1008 : OAI211_X1 port map( C1 => n553, C2 => IRAM_ADDRESS_28_port, A => 
                           n557, B => n552, ZN => n554);
   U1009 : NAND2_X1 port map( A1 => n555, A2 => n554, ZN => 
                           datapath_i_fetch_stage_dp_n9);
   U1010 : NAND2_X1 port map( A1 => n556, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, ZN => 
                           n562);
   U1011 : OAI211_X1 port map( C1 => n556, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, A => 
                           n563, B => n562, ZN => n560);
   U1012 : NAND2_X1 port map( A1 => n558, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n561);
   U1013 : OAI211_X1 port map( C1 => n558, C2 => IRAM_ADDRESS_30_port, A => 
                           n557, B => n561, ZN => n559);
   U1014 : NAND2_X1 port map( A1 => n560, A2 => n559, ZN => 
                           datapath_i_fetch_stage_dp_n3);
   U1015 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n561, Z => n565);
   U1016 : XOR2_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_31_port, 
                           B => n562, Z => n564);
   U1017 : AOI22_X1 port map( A1 => n566, A2 => n565, B1 => n564, B2 => n563, 
                           ZN => datapath_i_fetch_stage_dp_n2);
   U1018 : OAI21_X1 port map( B1 => n567, B2 => n737, A => n569, ZN => 
                           read_rf_p2_i);
   U1019 : OAI221_X1 port map( B1 => n570, B2 => n697, C1 => n569, C2 => n740, 
                           A => n568, ZN => datapath_i_decode_stage_dp_n78);
   U1020 : AND4_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           A2 => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           A3 => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           A4 => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ZN => n571);
   U1021 : AND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           A2 => n571, ZN => n587);
   U1022 : INV_X1 port map( A => n587, ZN => n596);
   U1023 : AND2_X2 port map( A1 => n596, A2 => n574, ZN => n610);
   U1024 : NOR2_X1 port map( A1 => n587, A2 => n574, ZN => n609);
   U1025 : CLKBUF_X1 port map( A => n609, Z => n600);
   U1026 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_0_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_0_port, ZN => n575);
   U1027 : OAI21_X1 port map( B1 => n733, B2 => n596, A => n575, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U1028 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_1_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_1_port, ZN => n576);
   U1029 : OAI21_X1 port map( B1 => n734, B2 => n596, A => n576, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U1030 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_2_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_2_port, ZN => n577);
   U1031 : OAI21_X1 port map( B1 => n728, B2 => n596, A => n577, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U1032 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_3_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_3_port, ZN => n578);
   U1033 : OAI21_X1 port map( B1 => n729, B2 => n596, A => n578, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U1034 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_4_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_4_port, ZN => n579);
   U1035 : OAI21_X1 port map( B1 => n730, B2 => n596, A => n579, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U1036 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_5_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_5_port, ZN => n580);
   U1037 : OAI21_X1 port map( B1 => n731, B2 => n596, A => n580, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U1038 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_6_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_6_port, ZN => n581);
   U1039 : OAI21_X1 port map( B1 => n732, B2 => n596, A => n581, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U1040 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_7_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_7_port, ZN => n582);
   U1041 : OAI21_X1 port map( B1 => n705, B2 => n596, A => n582, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U1042 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_8_port, B1 => n600, B2
                           => datapath_i_data_from_alu_i_8_port, ZN => n583);
   U1043 : OAI21_X1 port map( B1 => n706, B2 => n596, A => n583, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U1044 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_9_port, B1 => n609, B2
                           => datapath_i_data_from_alu_i_9_port, ZN => n584);
   U1045 : OAI21_X1 port map( B1 => n707, B2 => n596, A => n584, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U1046 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_10_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_10_port, ZN => n585
                           );
   U1047 : OAI21_X1 port map( B1 => n708, B2 => n596, A => n585, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U1048 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_11_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_11_port, ZN => n586
                           );
   U1049 : OAI21_X1 port map( B1 => n709, B2 => n596, A => n586, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U1050 : INV_X1 port map( A => n587, ZN => n612);
   U1051 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_12_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_12_port, ZN => n588
                           );
   U1052 : OAI21_X1 port map( B1 => n710, B2 => n612, A => n588, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U1053 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_13_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_13_port, ZN => n589
                           );
   U1054 : OAI21_X1 port map( B1 => n711, B2 => n596, A => n589, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U1055 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_14_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_14_port, ZN => n590
                           );
   U1056 : OAI21_X1 port map( B1 => n712, B2 => n612, A => n590, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U1057 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_15_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_15_port, ZN => n591
                           );
   U1058 : OAI21_X1 port map( B1 => n713, B2 => n596, A => n591, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U1059 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_16_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_16_port, ZN => n592
                           );
   U1060 : OAI21_X1 port map( B1 => n714, B2 => n612, A => n592, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U1061 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_17_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_17_port, ZN => n593
                           );
   U1062 : OAI21_X1 port map( B1 => n715, B2 => n596, A => n593, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U1063 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_18_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_18_port, ZN => n594
                           );
   U1064 : OAI21_X1 port map( B1 => n716, B2 => n612, A => n594, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U1065 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_19_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_19_port, ZN => n595
                           );
   U1066 : OAI21_X1 port map( B1 => n717, B2 => n596, A => n595, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U1067 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_20_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_20_port, ZN => n597
                           );
   U1068 : OAI21_X1 port map( B1 => n718, B2 => n612, A => n597, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U1069 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_21_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_21_port, ZN => n598
                           );
   U1070 : OAI21_X1 port map( B1 => n719, B2 => n612, A => n598, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U1071 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_22_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_22_port, ZN => n599
                           );
   U1072 : OAI21_X1 port map( B1 => n720, B2 => n612, A => n599, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U1073 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_23_port, B1 => n600, 
                           B2 => datapath_i_data_from_alu_i_23_port, ZN => n601
                           );
   U1074 : OAI21_X1 port map( B1 => n721, B2 => n612, A => n601, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U1075 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_24_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_24_port, ZN => n602
                           );
   U1076 : OAI21_X1 port map( B1 => n722, B2 => n612, A => n602, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U1077 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_25_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_25_port, ZN => n603
                           );
   U1078 : OAI21_X1 port map( B1 => n723, B2 => n612, A => n603, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U1079 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_26_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_26_port, ZN => n604
                           );
   U1080 : OAI21_X1 port map( B1 => n691, B2 => n612, A => n604, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U1081 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_27_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_27_port, ZN => n605
                           );
   U1082 : OAI21_X1 port map( B1 => n724, B2 => n612, A => n605, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U1083 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_28_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_28_port, ZN => n606
                           );
   U1084 : OAI21_X1 port map( B1 => n725, B2 => n612, A => n606, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U1085 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_29_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_29_port, ZN => n607
                           );
   U1086 : OAI21_X1 port map( B1 => n726, B2 => n612, A => n607, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U1087 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_30_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_30_port, ZN => n608
                           );
   U1088 : OAI21_X1 port map( B1 => n727, B2 => n612, A => n608, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U1089 : AOI22_X1 port map( A1 => n610, A2 => 
                           datapath_i_data_from_memory_i_31_port, B1 => n609, 
                           B2 => datapath_i_data_from_alu_i_31_port, ZN => n611
                           );
   U1090 : OAI21_X1 port map( B1 => n703, B2 => n612, A => n611, ZN => 
                           datapath_i_decode_stage_dp_n12);
   U1091 : AOI21_X1 port map( B1 => n633, B2 => n614, A => n613, ZN => n615);
   U1092 : NOR2_X1 port map( A1 => n616, A2 => n615, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U1093 : AOI22_X1 port map( A1 => n617, A2 => cu_i_cw1_10_port, B1 => 
                           cu_i_cmd_word_6_port, B2 => n704, ZN => n631);
   U1094 : NOR4_X1 port map( A1 => datapath_i_val_a_i_15_port, A2 => 
                           datapath_i_val_a_i_16_port, A3 => 
                           datapath_i_val_a_i_17_port, A4 => 
                           datapath_i_val_a_i_18_port, ZN => n621);
   U1095 : NOR4_X1 port map( A1 => datapath_i_val_a_i_19_port, A2 => 
                           datapath_i_val_a_i_20_port, A3 => 
                           datapath_i_val_a_i_21_port, A4 => 
                           datapath_i_val_a_i_22_port, ZN => n620);
   U1096 : NOR4_X1 port map( A1 => datapath_i_val_a_i_7_port, A2 => 
                           datapath_i_val_a_i_8_port, A3 => 
                           datapath_i_val_a_i_9_port, A4 => 
                           datapath_i_val_a_i_10_port, ZN => n619);
   U1097 : NOR4_X1 port map( A1 => datapath_i_val_a_i_11_port, A2 => 
                           datapath_i_val_a_i_12_port, A3 => 
                           datapath_i_val_a_i_13_port, A4 => 
                           datapath_i_val_a_i_14_port, ZN => n618);
   U1098 : NAND4_X1 port map( A1 => n621, A2 => n620, A3 => n619, A4 => n618, 
                           ZN => n627);
   U1099 : NOR4_X1 port map( A1 => datapath_i_val_a_i_30_port, A2 => 
                           datapath_i_val_a_i_31_port, A3 => 
                           datapath_i_val_a_i_1_port, A4 => 
                           datapath_i_val_a_i_2_port, ZN => n625);
   U1100 : NOR4_X1 port map( A1 => datapath_i_val_a_i_3_port, A2 => 
                           datapath_i_val_a_i_4_port, A3 => 
                           datapath_i_val_a_i_5_port, A4 => 
                           datapath_i_val_a_i_6_port, ZN => n624);
   U1101 : NOR4_X1 port map( A1 => datapath_i_val_a_i_23_port, A2 => 
                           datapath_i_val_a_i_24_port, A3 => 
                           datapath_i_val_a_i_25_port, A4 => 
                           datapath_i_val_a_i_26_port, ZN => n623);
   U1102 : NOR4_X1 port map( A1 => datapath_i_val_a_i_0_port, A2 => 
                           datapath_i_val_a_i_27_port, A3 => 
                           datapath_i_val_a_i_28_port, A4 => 
                           datapath_i_val_a_i_29_port, ZN => n622);
   U1103 : NAND4_X1 port map( A1 => n625, A2 => n624, A3 => n623, A4 => n622, 
                           ZN => n626);
   U1104 : NOR2_X1 port map( A1 => n627, A2 => n626, ZN => n629);
   U1105 : AOI22_X1 port map( A1 => cu_i_n4, A2 => cu_i_cw1_11_port, B1 => 
                           cu_i_cmd_word_7_port, B2 => n704, ZN => n628);
   U1106 : NAND2_X1 port map( A1 => n629, A2 => n628, ZN => n630);
   U1107 : OAI22_X1 port map( A1 => n631, A2 => n630, B1 => n629, B2 => n628, 
                           ZN => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port);
   U1108 : NOR2_X1 port map( A1 => n633, A2 => n632, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U1109 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port)
                           ;
   U1110 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port)
                           ;
   U1111 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port)
                           ;
   U1112 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           );
   U1113 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           );
   U1114 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           );
   U1115 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           );
   U1116 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           );
   U1117 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
                           ZN => n634);
   U1118 : NAND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
                           A2 => n310, ZN => n644);
   U1119 : OAI21_X1 port map( B1 => n310, B2 => n634, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           );
   U1120 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
                           ZN => n635);
   U1121 : OAI21_X1 port map( B1 => n310, B2 => n635, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           );
   U1122 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
                           ZN => n636);
   U1123 : OAI21_X1 port map( B1 => n310, B2 => n636, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           );
   U1124 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
                           ZN => n637);
   U1125 : OAI21_X1 port map( B1 => n765, B2 => n637, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           );
   U1126 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
                           ZN => n638);
   U1127 : OAI21_X1 port map( B1 => n765, B2 => n638, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           );
   U1128 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
                           ZN => n639);
   U1129 : OAI21_X1 port map( B1 => n310, B2 => n639, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           );
   U1130 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
                           ZN => n640);
   U1131 : OAI21_X1 port map( B1 => n765, B2 => n640, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           );
   U1132 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
                           ZN => n641);
   U1133 : OAI21_X1 port map( B1 => n310, B2 => n641, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           );
   U1134 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
                           ZN => n642);
   U1135 : OAI21_X1 port map( B1 => n765, B2 => n642, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           );
   U1136 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
                           ZN => n643);
   U1137 : OAI21_X1 port map( B1 => n310, B2 => n643, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           );
   U1138 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, S 
                           => n310, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port)
                           ;
   U1139 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
                           ZN => n645);
   U1140 : OAI21_X1 port map( B1 => n310, B2 => n645, A => n644, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           );
   U1141 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, S 
                           => n310, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port)
                           ;
   U1142 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port)
                           ;
   U1143 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port)
                           ;
   U1144 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port)
                           ;
   U1145 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port)
                           ;
   U1146 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, S 
                           => n765, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port)
                           ;
   U1147 : MUX2_X1 port map( A => datapath_i_val_b_i_7_port, B => 
                           datapath_i_val_immediate_i_7_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U1148 : MUX2_X1 port map( A => datapath_i_val_b_i_8_port, B => 
                           datapath_i_val_immediate_i_8_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U1149 : MUX2_X1 port map( A => datapath_i_val_b_i_9_port, B => 
                           datapath_i_val_immediate_i_9_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U1150 : MUX2_X1 port map( A => datapath_i_val_b_i_10_port, B => 
                           datapath_i_val_immediate_i_10_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_10_port);
   U1151 : MUX2_X1 port map( A => datapath_i_val_b_i_11_port, B => 
                           datapath_i_val_immediate_i_11_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_11_port);
   U1152 : MUX2_X1 port map( A => datapath_i_val_b_i_12_port, B => 
                           datapath_i_val_immediate_i_12_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_12_port);
   U1153 : MUX2_X1 port map( A => datapath_i_val_b_i_13_port, B => 
                           datapath_i_val_immediate_i_13_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_13_port);
   U1154 : MUX2_X1 port map( A => datapath_i_val_b_i_14_port, B => 
                           datapath_i_val_immediate_i_14_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_14_port);
   U1155 : MUX2_X1 port map( A => datapath_i_val_b_i_15_port, B => 
                           datapath_i_val_immediate_i_15_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_15_port);
   U1156 : MUX2_X1 port map( A => datapath_i_val_b_i_16_port, B => 
                           datapath_i_val_immediate_i_16_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_16_port);
   U1157 : MUX2_X1 port map( A => datapath_i_val_b_i_17_port, B => 
                           datapath_i_val_immediate_i_17_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_17_port);
   U1158 : MUX2_X1 port map( A => datapath_i_val_b_i_18_port, B => 
                           datapath_i_val_immediate_i_18_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_18_port);
   U1159 : MUX2_X1 port map( A => datapath_i_val_b_i_19_port, B => 
                           datapath_i_val_immediate_i_19_port, S => n647, Z => 
                           datapath_i_execute_stage_dp_opb_19_port);
   U1160 : MUX2_X1 port map( A => datapath_i_val_b_i_20_port, B => 
                           datapath_i_val_immediate_i_20_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_20_port);
   U1161 : MUX2_X1 port map( A => datapath_i_val_b_i_21_port, B => 
                           datapath_i_val_immediate_i_21_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_21_port);
   U1162 : MUX2_X1 port map( A => datapath_i_val_b_i_22_port, B => 
                           datapath_i_val_immediate_i_22_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_22_port);
   U1163 : MUX2_X1 port map( A => datapath_i_val_b_i_23_port, B => 
                           datapath_i_val_immediate_i_23_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_23_port);
   U1164 : MUX2_X1 port map( A => datapath_i_val_b_i_24_port, B => 
                           datapath_i_val_immediate_i_24_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_24_port);
   U1165 : NAND2_X1 port map( A1 => datapath_i_val_immediate_i_25_port, A2 => 
                           n647, ZN => n646);
   U1166 : OAI21_X1 port map( B1 => n647, B2 => n758, A => n646, ZN => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U1167 : OAI21_X1 port map( B1 => n647, B2 => n759, A => n646, ZN => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U1168 : OAI21_X1 port map( B1 => n647, B2 => n760, A => n646, ZN => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U1169 : OAI21_X1 port map( B1 => n647, B2 => n761, A => n646, ZN => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U1170 : OAI21_X1 port map( B1 => n647, B2 => n762, A => n646, ZN => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U1171 : OAI21_X1 port map( B1 => n647, B2 => n763, A => n646, ZN => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U1172 : OAI21_X1 port map( B1 => n647, B2 => n764, A => n646, ZN => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U1173 : MUX2_X1 port map( A => datapath_i_val_b_i_1_port, B => 
                           datapath_i_val_immediate_i_1_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U1174 : MUX2_X1 port map( A => datapath_i_val_b_i_3_port, B => 
                           datapath_i_val_immediate_i_3_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U1175 : MUX2_X1 port map( A => datapath_i_val_b_i_4_port, B => 
                           datapath_i_val_immediate_i_4_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U1176 : MUX2_X1 port map( A => datapath_i_val_b_i_5_port, B => 
                           datapath_i_val_immediate_i_5_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U1177 : MUX2_X1 port map( A => datapath_i_val_b_i_6_port, B => 
                           datapath_i_val_immediate_i_6_port, S => n648, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U1178 : NOR2_X1 port map( A1 => cu_i_n4, A2 => cu_i_n134, ZN => n650);
   U1179 : NOR2_X1 port map( A1 => n650, A2 => n649, ZN => n651);
   U1180 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n651, ZN => n685);
   U1181 : INV_X1 port map( A => n651, ZN => n674);
   U1182 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n674, ZN => n687);
   U1183 : CLKBUF_X1 port map( A => n687, Z => n676);
   U1184 : CLKBUF_X1 port map( A => n674, Z => n686);
   U1185 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n676, B1 => datapath_i_val_a_i_7_port, B2 => n686
                           , ZN => n652);
   U1186 : OAI21_X1 port map( B1 => n705, B2 => n689, A => n652, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U1187 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n676, B1 => datapath_i_val_a_i_8_port, B2 => n674
                           , ZN => n653);
   U1188 : OAI21_X1 port map( B1 => n706, B2 => n685, A => n653, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U1189 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n676, B1 => datapath_i_val_a_i_9_port, B2 => n686
                           , ZN => n654);
   U1190 : OAI21_X1 port map( B1 => n707, B2 => n685, A => n654, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U1191 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n676, B1 => datapath_i_val_a_i_10_port, B2 => 
                           n674, ZN => n655);
   U1192 : OAI21_X1 port map( B1 => n708, B2 => n685, A => n655, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U1193 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n676, B1 => datapath_i_val_a_i_11_port, B2 => 
                           n686, ZN => n656);
   U1194 : OAI21_X1 port map( B1 => n709, B2 => n685, A => n656, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U1195 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n676, B1 => datapath_i_val_a_i_12_port, B2 => 
                           n674, ZN => n657);
   U1196 : OAI21_X1 port map( B1 => n710, B2 => n685, A => n657, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U1197 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n676, B1 => datapath_i_val_a_i_13_port, B2 => 
                           n686, ZN => n658);
   U1198 : OAI21_X1 port map( B1 => n711, B2 => n685, A => n658, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U1199 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n676, B1 => datapath_i_val_a_i_14_port, B2 => 
                           n674, ZN => n659);
   U1200 : OAI21_X1 port map( B1 => n712, B2 => n685, A => n659, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U1201 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n676, B1 => datapath_i_val_a_i_15_port, B2 => 
                           n686, ZN => n660);
   U1202 : OAI21_X1 port map( B1 => n713, B2 => n685, A => n660, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U1203 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n687, B1 => datapath_i_val_a_i_16_port, B2 => 
                           n674, ZN => n661);
   U1204 : OAI21_X1 port map( B1 => n714, B2 => n689, A => n661, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U1205 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n687, B1 => datapath_i_val_a_i_17_port, B2 => 
                           n674, ZN => n662);
   U1206 : OAI21_X1 port map( B1 => n715, B2 => n689, A => n662, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U1207 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n687, B1 => datapath_i_val_a_i_18_port, B2 => 
                           n686, ZN => n663);
   U1208 : OAI21_X1 port map( B1 => n716, B2 => n689, A => n663, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U1209 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n676, B1 => datapath_i_val_a_i_19_port, B2 => 
                           n674, ZN => n664);
   U1210 : OAI21_X1 port map( B1 => n717, B2 => n689, A => n664, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U1211 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n676, B1 => datapath_i_val_a_i_20_port, B2 => 
                           n686, ZN => n665);
   U1212 : OAI21_X1 port map( B1 => n718, B2 => n689, A => n665, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U1213 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n676, B1 => datapath_i_val_a_i_21_port, B2 => 
                           n674, ZN => n666);
   U1214 : OAI21_X1 port map( B1 => n719, B2 => n689, A => n666, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U1215 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n676, B1 => datapath_i_val_a_i_22_port, B2 => 
                           n686, ZN => n667);
   U1216 : OAI21_X1 port map( B1 => n720, B2 => n689, A => n667, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U1217 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n676, B1 => datapath_i_val_a_i_23_port, B2 => 
                           n674, ZN => n668);
   U1218 : OAI21_X1 port map( B1 => n721, B2 => n689, A => n668, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U1219 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n676, B1 => datapath_i_val_a_i_24_port, B2 => 
                           n674, ZN => n669);
   U1220 : OAI21_X1 port map( B1 => n722, B2 => n689, A => n669, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U1221 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n676, B1 => datapath_i_val_a_i_25_port, B2 => 
                           n674, ZN => n670);
   U1222 : OAI21_X1 port map( B1 => n723, B2 => n689, A => n670, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U1223 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n676, B1 => datapath_i_val_a_i_26_port, B2 => 
                           n674, ZN => n671);
   U1224 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n676, B1 => datapath_i_val_a_i_0_port, B2 => n674
                           , ZN => n672);
   U1225 : OAI21_X1 port map( B1 => n685, B2 => n733, A => n672, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U1226 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n676, B1 => datapath_i_val_a_i_27_port, B2 => 
                           n674, ZN => n673);
   U1227 : OAI21_X1 port map( B1 => n724, B2 => n689, A => n673, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U1228 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n676, B1 => datapath_i_val_a_i_28_port, B2 => 
                           n674, ZN => n675);
   U1229 : OAI21_X1 port map( B1 => n725, B2 => n685, A => n675, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U1230 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n676, B1 => datapath_i_val_a_i_29_port, B2 => 
                           n686, ZN => n677);
   U1231 : OAI21_X1 port map( B1 => n726, B2 => n689, A => n677, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U1232 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n687, B1 => datapath_i_val_a_i_30_port, B2 => 
                           n686, ZN => n678);
   U1233 : OAI21_X1 port map( B1 => n727, B2 => n685, A => n678, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U1234 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n687, B1 => datapath_i_val_a_i_31_port, B2 => 
                           n686, ZN => n679);
   U1235 : OAI21_X1 port map( B1 => n703, B2 => n689, A => n679, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U1236 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n687, B1 => datapath_i_val_a_i_1_port, B2 => n686
                           , ZN => n680);
   U1237 : OAI21_X1 port map( B1 => n685, B2 => n734, A => n680, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U1238 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n687, B1 => datapath_i_val_a_i_2_port, B2 => n686
                           , ZN => n681);
   U1239 : OAI21_X1 port map( B1 => n728, B2 => n689, A => n681, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U1240 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n687, B1 => datapath_i_val_a_i_3_port, B2 => n686
                           , ZN => n682);
   U1241 : OAI21_X1 port map( B1 => n729, B2 => n685, A => n682, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U1242 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n687, B1 => datapath_i_val_a_i_4_port, B2 => n686
                           , ZN => n683);
   U1243 : OAI21_X1 port map( B1 => n730, B2 => n685, A => n683, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U1244 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n687, B1 => datapath_i_val_a_i_5_port, B2 => n686
                           , ZN => n684);
   U1245 : OAI21_X1 port map( B1 => n731, B2 => n685, A => n684, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U1246 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n687, B1 => datapath_i_val_a_i_6_port, B2 => n686
                           , ZN => n688);
   U1247 : OAI21_X1 port map( B1 => n732, B2 => n689, A => n688, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);

end SYN_dlx_rtl;
