
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_0_port, data2_mul_2_port, data2_mul_1_port, 
      dataout_mul_31_port, dataout_mul_30_port, dataout_mul_29_port, 
      dataout_mul_28_port, dataout_mul_27_port, dataout_mul_26_port, 
      dataout_mul_25_port, dataout_mul_24_port, dataout_mul_23_port, 
      dataout_mul_22_port, dataout_mul_21_port, dataout_mul_20_port, 
      dataout_mul_19_port, dataout_mul_18_port, dataout_mul_17_port, 
      dataout_mul_16_port, dataout_mul_15_port, dataout_mul_13_port, 
      dataout_mul_12_port, dataout_mul_11_port, dataout_mul_10_port, 
      dataout_mul_9_port, dataout_mul_8_port, dataout_mul_7_port, 
      dataout_mul_6_port, dataout_mul_5_port, dataout_mul_4_port, 
      dataout_mul_3_port, dataout_mul_2_port, dataout_mul_1_port, 
      dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521, N2522, N2523, 
      N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, 
      N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2543, 
      N2544, N2545, N2546, N2547, N2548, n554, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_34_port, 
      boothmul_pipelined_i_muxes_in_4_33_port, 
      boothmul_pipelined_i_muxes_in_4_32_port, 
      boothmul_pipelined_i_muxes_in_4_31_port, 
      boothmul_pipelined_i_muxes_in_4_30_port, 
      boothmul_pipelined_i_muxes_in_4_29_port, 
      boothmul_pipelined_i_muxes_in_4_28_port, 
      boothmul_pipelined_i_muxes_in_4_27_port, 
      boothmul_pipelined_i_sum_B_in_7_14_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_12_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_10_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_8_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_6_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_4_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_3_port, 
      boothmul_pipelined_i_sum_B_in_1_4_port, 
      boothmul_pipelined_i_sum_B_in_1_5_port, 
      boothmul_pipelined_i_sum_B_in_1_6_port, 
      boothmul_pipelined_i_sum_B_in_1_7_port, 
      boothmul_pipelined_i_sum_B_in_1_8_port, 
      boothmul_pipelined_i_sum_B_in_1_9_port, 
      boothmul_pipelined_i_sum_B_in_1_10_port, 
      boothmul_pipelined_i_sum_B_in_1_11_port, 
      boothmul_pipelined_i_sum_B_in_1_12_port, 
      boothmul_pipelined_i_sum_B_in_1_13_port, 
      boothmul_pipelined_i_sum_B_in_1_14_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_6_28_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_5_26_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_4_24_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_3_22_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_7_15_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n1068, 
      n1084, n1094, n1095, n1102, n1104, n1105, n1109, n1110, n1120, n1129, 
      n1142, n1157, n1167, n1178, n1194, n1203, n1219, n1235, n1236, n1247, 
      n1249, n1254, n1256, n1277, n1278, n1286, n1301, n1302, n1319, n1321, 
      n1322, n1324, n1328, n1334, n1349, n1353, n1354, n1366, n1389, n1392, 
      n1393, n1394, n1403, n1425, n1428, n1429, n1430, n1441, n1467, n1469, 
      n1470, n1531, n1534, n1535, n1537, n1542, n1546, n1550, n1556, n1559, 
      n1560, n1580, n1581, n1584, n1593, n1594, n1595, n1615, n1633, n1655, 
      n1677, n1680, n1682, n1708, n1720, n1722, n1724, n1728, n1803, n1974, 
      n1976, n1978, n1979, n1986, n2008, n2011, n2026, n2028, n2031, n2052, 
      n2058, n2070, n2075, n2078, n2082, n2084, n2085, n2094, n2097, n2116, 
      n2127, n2131, n2134, n2143, n2144, n2150, n2157, n2161, n2163, n2165, 
      n2204, n2209, n2210, n2212, n2219, n2220, n2226, n2240, n2244, n2245, 
      n2250, n2261, n2262, n2264, n2267, n2271, n2275, n2294, n2300, n2313, 
      n2319, n2321, n2322, n2323, n2332, n2333, n2337, n2338, n2340, n2355, 
      n2361, n2378, n2379, n2381, n2399, n2401, n2403, n2407, n2425, n2433, 
      n2435, n2441, n2445, n2513, n2519_port, n2520_port, n2521_port, 
      n2527_port, n2529_port, n2539_port, n2541_port, n2542_port, n2594, n2595,
      n2596, n2622, n2635, n2669, n2670, n2671, n2672, n2690, n2693, n2694, 
      n2773, n2802, n2806, n2808, n3020, n3026, n3027, n3028, n3029, n3030, 
      n3036, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3802, n3804, 
      n3805, n3807, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, 
      n3817, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3875, n3876, n3877, n3878, 
      n3879, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, 
      n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, 
      n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3910, 
      n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, 
      n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, 
      n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, 
      n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, 
      n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, 
      n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3970, n3971, 
      n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, 
      n3982, n3983, n3984, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4003, 
      n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, 
      n4014, n4015, n4016, n4017, n4018, n4020, n4021, n4022, n4023, n4024, 
      n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, 
      n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, 
      n4045, n4046, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, 
      n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, 
      n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, 
      n4076, n4077, n4078, n4079, n4081, n4082, n4083, n4084, n4085, n4086, 
      n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, 
      n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, 
      n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, 
      n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, 
      n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, 
      n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, 
      n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, 
      n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4298, n4299, 
      n4300, n4302, n4303, n4304, n4305, n4306, n4308, n4309, n4310, n4311, 
      n4312, n4313, n4314, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, 
      n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4542, n4545, n4546, 
      n4548, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
      n6015, n6016, n6017, n6018, n6019, n6021, n6022, n6023, n1840, n1841, 
      n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, 
      n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, 
      n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, 
      n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, 
      n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, 
      n1892, n1893, n1894, n1895, n1896, n1898, n1900, n1901, n1902, n1903, 
      n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, 
      n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
      n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, 
      n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, 
      n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
      n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, 
      n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
      n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, 
      n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
      n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, 
      n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, 
      n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, 
      n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
      n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, 
      n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, 
      n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, 
      n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
      n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, 
      n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
      n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
      n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
      n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
      n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
      n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
      n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
      n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, 
      n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
      n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
      n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
      n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
      n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
      n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
      n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
      n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, 
      n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, 
      n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
      n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, 
      n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, 
      n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
      n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, 
      n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, 
      n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, 
      n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, 
      n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
      n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
      n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, 
      n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
      n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, 
      n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, 
      n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, 
      n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, 
      n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, 
      n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, 
      n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
      n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, 
      n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, 
      n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, 
      n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, 
      n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, 
      n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, 
      n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, 
      n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, 
      n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, 
      n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, 
      n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
      n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
      n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, 
      n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, 
      n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, 
      n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, 
      n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, 
      n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
      n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, 
      n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, 
      n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, 
      n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, 
      n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, 
      n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, 
      n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, 
      n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, 
      n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, 
      n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, 
      n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, 
      n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, 
      n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, 
      n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, 
      n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, 
      n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, 
      n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, 
      n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, 
      n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, 
      n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, 
      n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, 
      n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, 
      n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, 
      n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, 
      n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, 
      n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, 
      n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, 
      n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, 
      n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, 
      n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, 
      n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, 
      n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, 
      n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, 
      n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, 
      n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, 
      n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, 
      n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, 
      n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, 
      n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, 
      n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, 
      n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, 
      n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, 
      n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, 
      n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, 
      n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, 
      n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, 
      n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, 
      n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, 
      n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, 
      n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, 
      n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, 
      n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, 
      n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, 
      n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, 
      n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, 
      n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, 
      n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, 
      n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, 
      n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, 
      n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, 
      n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, 
      n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, 
      n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, 
      n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, 
      n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, 
      n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, 
      n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, 
      n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, 
      n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, 
      n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, 
      n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, 
      n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, 
      n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, 
      n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, 
      n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, 
      n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, 
      n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, 
      n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, 
      n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, 
      n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, 
      n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n_1004, n_1005, 
      n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, 
      n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, 
      n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, 
      n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, 
      n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, 
      n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, 
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, 
      n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, 
      n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, 
      n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, 
      n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, 
      n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, 
      n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, 
      n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, 
      n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, 
      n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, 
      n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, 
      n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, 
      n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, 
      n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, 
      n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, 
      n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, 
      n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, 
      n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, 
      n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, 
      n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, 
      n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, 
      n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, 
      n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, 
      n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, 
      n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, 
      n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, 
      n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, 
      n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, 
      n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, 
      n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, 
      n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, 
      n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, 
      n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, 
      n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, 
      n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, 
      n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, 
      n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, 
      n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, 
      n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, 
      n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, 
      n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, 
      n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, 
      n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, 
      n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, 
      n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, 
      n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, 
      n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, 
      n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, 
      n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, 
      n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, 
      n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, 
      n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, 
      n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671 : 
      std_logic;

begin
   
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n554, Q => 
                           DATA2_I_29_port);
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n554, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n554, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n554, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n554, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n554, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n554, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n554, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n554, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n554, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n7829, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n7829, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n554, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n7829, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n7829, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n7829, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n7829, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n7829, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n554, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n554, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n554, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n554, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n554, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n554, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n554, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n7829, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n554, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n554, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n554, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n554, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n7822, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => DATA1(14), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_27_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_28_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => DATA1(12), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_29_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_30_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => DATA1(10), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_31_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_32_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_33_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_34_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => DATA1(3), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n7822, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n7822, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n7822, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n7822, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n7829, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1893, B => n1894, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1891, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1889, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1887, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1885, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1883, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1881, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1879, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1877, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1875, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1873, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1871, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1869, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1867, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1865, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_3_port, CI => n3036,
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => dataout_mul_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_4_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_5_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_6_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_7_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_8_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_9_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_10_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_11_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_12_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_13_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_14_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_2_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1004, S => 
                           boothmul_pipelined_i_sum_B_in_2_20_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => n4046, 
                           CI => n3026, CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => dataout_mul_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => n4045, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => n4044, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => n4043, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => n4042, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => n4041, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => n4040, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => n4039, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => n4038, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => n4037, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => n4036, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => n4035, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => n4034, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => n4033, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => n4033, 
                           CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_3_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n3800, B => n4032, CI => n4026, CO => n_1005, S => 
                           boothmul_pipelined_i_sum_B_in_3_22_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3030,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => dataout_mul_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           n4190, B => n4025, CI => n4009, CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           n4189, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           n4188, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_4_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n4187, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1006, S => 
                           boothmul_pipelined_i_sum_B_in_4_24_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => n4018, 
                           CI => n3029, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => dataout_mul_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => n4017, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => n4016, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => n4015, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => n4014, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => n4013, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => n4012, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => n4011, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => n4010, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => n4008, 
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n4186, B => n4007, CI => n3991, CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           n4185, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_B_in_5_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n4184, B => n4007, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1007, S => 
                           boothmul_pipelined_i_sum_B_in_5_26_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => n4001, 
                           CI => n3028, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => dataout_mul_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => n4000, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => n3999, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => n3998, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => n3997, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => n3996, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => n3995, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => n3994, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => n3993, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => n3992, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => n3990, 
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n4183, B => n3989, CI => n3974, CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           n4182, B => n3989, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_B_in_6_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n4181, B => n3989, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1008, S => 
                           boothmul_pipelined_i_sum_B_in_6_28_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => n3984, 
                           CI => n3027, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => dataout_mul_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => n3983, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => n3982, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => n3981, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => n3980, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => n3979, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => n3978, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => n3977, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => n3976, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => n3975, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => n3973, 
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n4180, B => n3972, CI => n3958, CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           n4179, B => n3972, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_B_in_7_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n4178, B => n3972, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1009, S => 
                           boothmul_pipelined_i_sum_B_in_7_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => n3968, 
                           CI => n3020, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => n3967, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => n3966, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => n3965, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => n3964, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => n3963, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => n3962, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => n3961, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => n3960, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => n3959, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => n3957, 
                           CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n4177, B => n3956, CI => n3940, CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           n4176, B => n3956, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           n4175, B => n3956, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           n4175, B => n3956, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1010, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n7822, Q => 
                           data2_mul_1_port);
   clk_r_REG3467_S7 : DFFR_X1 port map( D => n1903, CK => clk, RN => n6055, Q 
                           => n_1011, QN => n4548);
   clk_r_REG3456_S7 : DFFR_X1 port map( D => n1904, CK => clk, RN => rst_BAR, Q
                           => n_1012, QN => n4546);
   clk_r_REG3465_S7 : DFFS_X1 port map( D => n1905, CK => clk, SN => rst_BAR, Q
                           => n_1013, QN => n4545);
   clk_r_REG117_S52 : DFFS_X1 port map( D => DATA1(31), CK => clk, SN => 
                           rst_BAR, Q => n7726, QN => n5995);
   clk_r_REG113_S51 : DFFR_X1 port map( D => DATA1(30), CK => clk, RN => 
                           rst_BAR, Q => n7742, QN => n6022);
   clk_r_REG112_S51 : DFFS_X1 port map( D => DATA1(30), CK => clk, SN => 
                           rst_BAR, Q => n4542, QN => n_1014);
   clk_r_REG107_S49 : DFFR_X1 port map( D => DATA1(29), CK => clk, RN => 
                           rst_BAR, Q => n7762, QN => n6016);
   clk_r_REG106_S49 : DFFS_X1 port map( D => DATA1(29), CK => clk, SN => 
                           rst_BAR, Q => n4540, QN => n_1015);
   clk_r_REG101_S48 : DFFR_X1 port map( D => n1906, CK => clk, RN => n6056, Q 
                           => n_1016, QN => n4539);
   clk_r_REG92_S46 : DFFR_X1 port map( D => n1907, CK => clk, RN => rst_BAR, Q 
                           => n_1017, QN => n4538);
   clk_r_REG86_S45 : DFFS_X1 port map( D => n1910, CK => clk, SN => rst_BAR, Q 
                           => n_1018, QN => n4537);
   clk_r_REG80_S43 : DFFS_X1 port map( D => n1911, CK => clk, SN => rst_BAR, Q 
                           => n_1019, QN => n4536);
   clk_r_REG62_S38 : DFFR_X1 port map( D => n1922, CK => clk, RN => n6054, Q =>
                           n_1020, QN => n4535);
   clk_r_REG51_S35 : DFFR_X1 port map( D => n1925, CK => clk, RN => rst_BAR, Q 
                           => n_1021, QN => n4534);
   clk_r_REG43_S32 : DFFR_X1 port map( D => n1929, CK => clk, RN => rst_BAR, Q 
                           => n_1022, QN => n4533);
   clk_r_REG334_S7 : DFFR_X1 port map( D => n1933, CK => clk, RN => rst_BAR, Q 
                           => n_1023, QN => n4532);
   clk_r_REG20_S14 : DFFR_X1 port map( D => n1939, CK => clk, RN => rst_BAR, Q 
                           => n_1024, QN => n4531);
   clk_r_REG126_S3 : DFFR_X1 port map( D => n1941, CK => clk, RN => rst_BAR, Q 
                           => n_1025, QN => n4530);
   clk_r_REG2176_S3 : DFFS_X1 port map( D => n1942, CK => clk, SN => rst_BAR, Q
                           => n_1026, QN => n4529);
   clk_r_REG2253_S3 : DFFR_X1 port map( D => n1943, CK => clk, RN => rst_BAR, Q
                           => n_1027, QN => n4528);
   clk_r_REG2327_S3 : DFFR_X1 port map( D => n1944, CK => clk, RN => rst_BAR, Q
                           => n_1028, QN => n4527);
   clk_r_REG2642_S3 : DFFS_X1 port map( D => n1945, CK => clk, SN => rst_BAR, Q
                           => n_1029, QN => n4526);
   clk_r_REG390_S3 : DFFR_X1 port map( D => n1946, CK => clk, RN => rst_BAR, Q 
                           => n_1030, QN => n4525);
   clk_r_REG1491_S3 : DFFR_X1 port map( D => n1970, CK => clk, RN => n6055, Q 
                           => n_1031, QN => n4524);
   clk_r_REG3249_S2 : DFFR_X1 port map( D => cin, CK => clk, RN => n6054, Q => 
                           n4523, QN => n_1032);
   clk_r_REG660_S3 : DFFS_X1 port map( D => n7827, CK => clk, SN => rst_BAR, Q 
                           => n4522, QN => n_1033);
   clk_r_REG591_S3 : DFFR_X1 port map( D => n1950, CK => clk, RN => rst_BAR, Q 
                           => n4520, QN => n7790);
   clk_r_REG605_S3 : DFFR_X1 port map( D => n1068, CK => clk, RN => rst_BAR, Q 
                           => n4517, QN => n7741);
   clk_r_REG604_S3 : DFFS_X1 port map( D => n1068, CK => clk, SN => rst_BAR, Q 
                           => n4516, QN => n_1034);
   clk_r_REG664_S3 : DFFR_X1 port map( D => n7709, CK => clk, RN => rst_BAR, Q 
                           => n4515, QN => n_1035);
   clk_r_REG3457_S7 : DFFS_X1 port map( D => n1904, CK => clk, SN => rst_BAR, Q
                           => n4514, QN => n_1036);
   clk_r_REG3466_S7 : DFFR_X1 port map( D => n1905, CK => clk, RN => n6054, Q 
                           => n4513, QN => n7816);
   clk_r_REG566_S3 : DFFS_X1 port map( D => n1959, CK => clk, SN => rst_BAR, Q 
                           => n4512, QN => n7731);
   clk_r_REG651_S3 : DFFR_X1 port map( D => n7709, CK => clk, RN => rst_BAR, Q 
                           => n_1037, QN => n4511);
   clk_r_REG514_S10 : DFFR_X1 port map( D => n7823, CK => clk, RN => rst_BAR, Q
                           => n4510, QN => n_1038);
   clk_r_REG3463_S7 : DFFR_X1 port map( D => n7821, CK => clk, RN => n6054, Q 
                           => n4509, QN => n_1039);
   clk_r_REG538_S3 : DFFR_X1 port map( D => n6023, CK => clk, RN => n6055, Q =>
                           n4508, QN => n7748);
   clk_r_REG565_S3 : DFFS_X1 port map( D => n1962, CK => clk, SN => rst_BAR, Q 
                           => n4507, QN => n7804);
   clk_r_REG549_S3 : DFFR_X1 port map( D => n1964, CK => clk, RN => rst_BAR, Q 
                           => n4506, QN => n7757);
   clk_r_REG584_S3 : DFFR_X1 port map( D => n1949, CK => clk, RN => rst_BAR, Q 
                           => n4505, QN => n7770);
   clk_r_REG613_S3 : DFFR_X1 port map( D => n1952, CK => clk, RN => rst_BAR, Q 
                           => n4504, QN => n_1040);
   clk_r_REG612_S3 : DFFS_X1 port map( D => n1952, CK => clk, SN => rst_BAR, Q 
                           => n4503, QN => n_1041);
   clk_r_REG623_S3 : DFFR_X1 port map( D => n7826, CK => clk, RN => rst_BAR, Q 
                           => n4502, QN => n_1042);
   clk_r_REG622_S3 : DFFS_X1 port map( D => n7825, CK => clk, SN => rst_BAR, Q 
                           => n4501, QN => n_1043);
   clk_r_REG670_S3 : DFFR_X1 port map( D => n7824, CK => clk, RN => rst_BAR, Q 
                           => n4500, QN => n_1044);
   clk_r_REG669_S3 : DFFS_X1 port map( D => n7824, CK => clk, SN => rst_BAR, Q 
                           => n4499, QN => n_1045);
   clk_r_REG594_S3 : DFFS_X1 port map( D => n1958, CK => clk, SN => rst_BAR, Q 
                           => n_1046, QN => n4498);
   clk_r_REG593_S3 : DFFR_X1 port map( D => n1958, CK => clk, RN => rst_BAR, Q 
                           => n_1047, QN => n4497);
   clk_r_REG602_S3 : DFFR_X1 port map( D => n1958, CK => clk, RN => rst_BAR, Q 
                           => n4496, QN => n_1048);
   clk_r_REG601_S3 : DFFS_X1 port map( D => n1958, CK => clk, SN => rst_BAR, Q 
                           => n4495, QN => n_1049);
   clk_r_REG1794_S42 : DFFS_X1 port map( D => n1914, CK => clk, SN => rst_BAR, 
                           Q => n4494, QN => n_1050);
   clk_r_REG2715_S39 : DFFS_X1 port map( D => n1921, CK => clk, SN => rst_BAR, 
                           Q => n4493, QN => n_1051);
   clk_r_REG668_S3 : DFFR_X1 port map( D => n7824, CK => clk, RN => rst_BAR, Q 
                           => n4492, QN => n_1052);
   clk_r_REG2711_S42 : DFFS_X1 port map( D => n1912, CK => clk, SN => rst_BAR, 
                           Q => n4491, QN => n_1053);
   clk_r_REG2555_S45 : DFFS_X1 port map( D => n1910, CK => clk, SN => rst_BAR, 
                           Q => n4490, QN => n_1054);
   clk_r_REG587_S3 : DFFS_X1 port map( D => n1950, CK => clk, SN => rst_BAR, Q 
                           => n7725, QN => n4489);
   clk_r_REG655_S3 : DFFR_X1 port map( D => n7828, CK => clk, RN => rst_BAR, Q 
                           => n4488, QN => n7818);
   clk_r_REG618_S3 : DFFS_X1 port map( D => n1917, CK => clk, SN => n6054, Q =>
                           n4487, QN => n7785);
   clk_r_REG609_S3 : DFFS_X1 port map( D => n1952, CK => clk, SN => rst_BAR, Q 
                           => n_1055, QN => n4486);
   clk_r_REG608_S3 : DFFR_X1 port map( D => n1952, CK => clk, RN => rst_BAR, Q 
                           => n_1056, QN => n4485);
   clk_r_REG611_S3 : DFFR_X1 port map( D => n1952, CK => clk, RN => rst_BAR, Q 
                           => n4484, QN => n_1057);
   clk_r_REG610_S3 : DFFS_X1 port map( D => n1952, CK => clk, SN => n6055, Q =>
                           n4483, QN => n_1058);
   clk_r_REG597_S3 : DFFS_X1 port map( D => n1958, CK => clk, SN => rst_BAR, Q 
                           => n4482, QN => n_1059);
   clk_r_REG617_S3 : DFFS_X1 port map( D => n1913, CK => clk, SN => rst_BAR, Q 
                           => n4481, QN => n7784);
   clk_r_REG545_S3 : DFFS_X1 port map( D => n1965, CK => clk, SN => rst_BAR, Q 
                           => n7763, QN => n4480);
   clk_r_REG547_S3 : DFFR_X1 port map( D => n1965, CK => clk, RN => rst_BAR, Q 
                           => n4479, QN => n_1060);
   clk_r_REG571_S3 : DFFR_X1 port map( D => n1947, CK => clk, RN => rst_BAR, Q 
                           => n4476, QN => n7761);
   clk_r_REG578_S3 : DFFR_X1 port map( D => n5994, CK => clk, RN => rst_BAR, Q 
                           => n4475, QN => n7768);
   clk_r_REG582_S3 : DFFS_X1 port map( D => n5992, CK => clk, SN => rst_BAR, Q 
                           => n4474, QN => n7767);
   clk_r_REG567_S3 : DFFS_X1 port map( D => n1102, CK => clk, SN => n6054, Q =>
                           n4473, QN => n7734);
   clk_r_REG569_S3 : DFFR_X1 port map( D => n2332, CK => clk, RN => rst_BAR, Q 
                           => n7727, QN => n4472);
   clk_r_REG570_S3 : DFFR_X1 port map( D => n2332, CK => clk, RN => rst_BAR, Q 
                           => n4471, QN => n7766);
   clk_r_REG637_S32 : DFFR_X1 port map( D => n1927, CK => clk, RN => n6057, Q 
                           => n4470, QN => n_1061);
   clk_r_REG583_S3 : DFFS_X1 port map( D => n5992, CK => clk, SN => rst_BAR, Q 
                           => n4469, QN => n_1062);
   clk_r_REG573_S3 : DFFR_X1 port map( D => n5997, CK => clk, RN => n6056, Q =>
                           n4468, QN => n7719);
   clk_r_REG633_S7 : DFFR_X1 port map( D => n1930, CK => clk, RN => rst_BAR, Q 
                           => n4467, QN => n_1063);
   clk_r_REG577_S3 : DFFR_X1 port map( D => n5994, CK => clk, RN => rst_BAR, Q 
                           => n4466, QN => n7722);
   clk_r_REG630_S7 : DFFR_X1 port map( D => n1932, CK => clk, RN => rst_BAR, Q 
                           => n4465, QN => n_1064);
   clk_r_REG674_S3 : DFFR_X1 port map( D => n1960, CK => clk, RN => n6057, Q =>
                           n4464, QN => n7736);
   clk_r_REG543_S3 : DFFS_X1 port map( D => n6003, CK => clk, SN => rst_BAR, Q 
                           => n4463, QN => n7723);
   clk_r_REG561_S3 : DFFS_X1 port map( D => n1963, CK => clk, SN => rst_BAR, Q 
                           => n4462, QN => n7794);
   clk_r_REG557_S3 : DFFR_X1 port map( D => n1961, CK => clk, RN => n6055, Q =>
                           n4461, QN => n7808);
   clk_r_REG559_S3 : DFFR_X1 port map( D => n6000, CK => clk, RN => n6057, Q =>
                           n4460, QN => n_1065);
   clk_r_REG585_S3 : DFFS_X1 port map( D => n1949, CK => clk, SN => rst_BAR, Q 
                           => n4459, QN => n7772);
   clk_r_REG2397_S48 : DFFR_X1 port map( D => n1906, CK => clk, RN => rst_BAR, 
                           Q => n4458, QN => n_1066);
   clk_r_REG2396_S48 : DFFS_X1 port map( D => n1906, CK => clk, SN => rst_BAR, 
                           Q => n4457, QN => n_1067);
   clk_r_REG551_S3 : DFFR_X1 port map( D => n5987, CK => clk, RN => rst_BAR, Q 
                           => n4456, QN => n7730);
   clk_r_REG548_S3 : DFFR_X1 port map( D => n1219, CK => clk, RN => rst_BAR, Q 
                           => n4455, QN => n7720);
   clk_r_REG541_S3 : DFFR_X1 port map( D => n5996, CK => clk, RN => rst_BAR, Q 
                           => n4454, QN => n7801);
   clk_r_REG563_S3 : DFFR_X1 port map( D => n5991, CK => clk, RN => rst_BAR, Q 
                           => n4453, QN => n7749);
   clk_r_REG510_S7 : DFFS_X1 port map( D => n5990, CK => clk, SN => rst_BAR, Q 
                           => n4452, QN => n_1068);
   clk_r_REG505_S10 : DFFS_X1 port map( D => n1859, CK => clk, SN => rst_BAR, Q
                           => n4451, QN => n_1069);
   clk_r_REG3462_S7 : DFFR_X1 port map( D => n1900, CK => clk, RN => rst_BAR, Q
                           => n4450, QN => n_1070);
   clk_r_REG3459_S7 : DFFR_X1 port map( D => n1901, CK => clk, RN => n6057, Q 
                           => n4449, QN => n7817);
   clk_r_REG491_S7 : DFFS_X1 port map( D => n1937, CK => clk, SN => rst_BAR, Q 
                           => n4448, QN => n_1071);
   clk_r_REG534_S3 : DFFR_X1 port map( D => n1902, CK => clk, RN => rst_BAR, Q 
                           => n4447, QN => n7803);
   clk_r_REG832_S7 : DFFS_X1 port map( D => n1858, CK => clk, SN => rst_BAR, Q 
                           => n4446, QN => n_1072);
   clk_r_REG931_S3 : DFFS_X1 port map( D => n1967, CK => clk, SN => rst_BAR, Q 
                           => n4445, QN => n7797);
   clk_r_REG933_S3 : DFFS_X1 port map( D => n1966, CK => clk, SN => rst_BAR, Q 
                           => n4444, QN => n_1073);
   clk_r_REG930_S3 : DFFR_X1 port map( D => n5986, CK => clk, RN => rst_BAR, Q 
                           => n4443, QN => n7747);
   clk_r_REG917_S10 : DFFR_X1 port map( D => n1861, CK => clk, RN => rst_BAR, Q
                           => n4442, QN => n_1074);
   clk_r_REG922_S3 : DFFS_X1 port map( D => n1969, CK => clk, SN => rst_BAR, Q 
                           => n4441, QN => n_1075);
   clk_r_REG921_S3 : DFFR_X1 port map( D => n5999, CK => clk, RN => rst_BAR, Q 
                           => n4440, QN => n_1076);
   clk_r_REG556_S3 : DFFS_X1 port map( D => n6002, CK => clk, SN => rst_BAR, Q 
                           => n4439, QN => n7805);
   clk_r_REG456_S10 : DFFS_X1 port map( D => n1936, CK => clk, SN => rst_BAR, Q
                           => n4438, QN => n_1077);
   clk_r_REG511_S10 : DFFS_X1 port map( D => n7823, CK => clk, SN => rst_BAR, Q
                           => n4437, QN => n_1078);
   clk_r_REG554_S3 : DFFS_X1 port map( D => n6001, CK => clk, SN => rst_BAR, Q 
                           => n4436, QN => n_1079);
   clk_r_REG644_S35 : DFFR_X1 port map( D => n1926, CK => clk, RN => rst_BAR, Q
                           => n4435, QN => n_1080);
   clk_r_REG355_S35 : DFFR_X1 port map( D => n1928, CK => clk, RN => rst_BAR, Q
                           => n4434, QN => n_1081);
   clk_r_REG615_S32 : DFFR_X1 port map( D => n1931, CK => clk, RN => n6055, Q 
                           => n4433, QN => n7788);
   clk_r_REG171_S42 : DFFR_X1 port map( D => n1915, CK => clk, RN => rst_BAR, Q
                           => n4432, QN => n_1082);
   clk_r_REG648_S39 : DFFR_X1 port map( D => n1918, CK => clk, RN => rst_BAR, Q
                           => n4431, QN => n_1083);
   clk_r_REG596_S3 : DFFR_X1 port map( D => n1919, CK => clk, RN => rst_BAR, Q 
                           => n4430, QN => n_1084);
   clk_r_REG173_S42 : DFFR_X1 port map( D => n1916, CK => clk, RN => n6055, Q 
                           => n4429, QN => n_1085);
   clk_r_REG315_S32 : DFFR_X1 port map( D => n1924, CK => clk, RN => rst_BAR, Q
                           => n4428, QN => n_1086);
   clk_r_REG636_S46 : DFFS_X1 port map( D => n1908, CK => clk, SN => rst_BAR, Q
                           => n4427, QN => n_1087);
   clk_r_REG467_S6 : DFFR_X1 port map( D => n1934, CK => clk, RN => n6054, Q =>
                           n4426, QN => n_1088);
   clk_r_REG422_S24 : DFFR_X1 port map( D => n1935, CK => clk, RN => rst_BAR, Q
                           => n4425, QN => n_1089);
   clk_r_REG926_S3 : DFFS_X1 port map( D => n5998, CK => clk, SN => rst_BAR, Q 
                           => n4424, QN => n7753);
   clk_r_REG742_S6 : DFFS_X1 port map( D => n1857, CK => clk, SN => rst_BAR, Q 
                           => n4423, QN => n_1090);
   clk_r_REG1875_S4 : DFFS_X1 port map( D => n1847, CK => clk, SN => rst_BAR, Q
                           => n4422, QN => n_1091);
   clk_r_REG2410_S46 : DFFS_X1 port map( D => n1840, CK => clk, SN => rst_BAR, 
                           Q => n4421, QN => n_1092);
   clk_r_REG2569_S43 : DFFS_X1 port map( D => n1843, CK => clk, SN => rst_BAR, 
                           Q => n4420, QN => n_1093);
   clk_r_REG2567_S42 : DFFS_X1 port map( D => n6017, CK => clk, SN => n6057, Q 
                           => n4419, QN => n_1094);
   clk_r_REG168_S42 : DFFS_X1 port map( D => n1846, CK => clk, SN => rst_BAR, Q
                           => n4418, QN => n7752);
   clk_r_REG170_S42 : DFFR_X1 port map( D => n6018, CK => clk, RN => rst_BAR, Q
                           => n4417, QN => n7754);
   clk_r_REG924_S3 : DFFR_X1 port map( D => n5988, CK => clk, RN => rst_BAR, Q 
                           => n4416, QN => n7814);
   clk_r_REG2179_S3 : DFFS_X1 port map( D => n1942, CK => clk, SN => rst_BAR, Q
                           => n4415, QN => n7815);
   clk_r_REG2255_S3 : DFFS_X1 port map( D => n1943, CK => clk, SN => rst_BAR, Q
                           => n4414, QN => n_1095);
   clk_r_REG2331_S3 : DFFS_X1 port map( D => n1944, CK => clk, SN => rst_BAR, Q
                           => n4413, QN => n_1096);
   clk_r_REG2487_S45 : DFFS_X1 port map( D => n1842, CK => clk, SN => rst_BAR, 
                           Q => n4412, QN => n_1097);
   clk_r_REG2489_S45 : DFFS_X1 port map( D => n6015, CK => clk, SN => rst_BAR, 
                           Q => n4411, QN => n_1098);
   clk_r_REG2409_S46 : DFFS_X1 port map( D => n1841, CK => clk, SN => rst_BAR, 
                           Q => n4410, QN => n_1099);
   clk_r_REG69_S39 : DFFS_X1 port map( D => n1849, CK => clk, SN => rst_BAR, Q 
                           => n4409, QN => n_1100);
   clk_r_REG305_S8 : DFFS_X1 port map( D => n1855, CK => clk, SN => n6055, Q =>
                           n4408, QN => n_1101);
   clk_r_REG70_S39 : DFFS_X1 port map( D => n1848, CK => clk, SN => rst_BAR, Q 
                           => n4407, QN => n_1102);
   clk_r_REG156_S35 : DFFS_X1 port map( D => n1851, CK => clk, SN => rst_BAR, Q
                           => n4406, QN => n_1103);
   clk_r_REG2724_S38 : DFFS_X1 port map( D => n1850, CK => clk, SN => rst_BAR, 
                           Q => n4405, QN => n_1104);
   clk_r_REG2800_S36 : DFFS_X1 port map( D => n1852, CK => clk, SN => rst_BAR, 
                           Q => n4404, QN => n_1105);
   clk_r_REG153_S35 : DFFS_X1 port map( D => n1853, CK => clk, SN => rst_BAR, Q
                           => n4403, QN => n_1106);
   clk_r_REG2941_S32 : DFFS_X1 port map( D => n1854, CK => clk, SN => rst_BAR, 
                           Q => n4402, QN => n_1107);
   clk_r_REG620_S10 : DFFR_X1 port map( D => n1938, CK => clk, RN => rst_BAR, Q
                           => n4401, QN => n_1108);
   clk_r_REG3464_S7 : DFFS_X1 port map( D => n1898, CK => clk, SN => n6054, Q 
                           => n4400, QN => n_1109);
   clk_r_REG528_S4 : DFFR_X1 port map( D => n6004, CK => clk, RN => rst_BAR, Q 
                           => n4399, QN => n_1110);
   clk_r_REG531_S4 : DFFS_X1 port map( D => n5989, CK => clk, SN => n6056, Q =>
                           n4398, QN => n_1111);
   clk_r_REG2178_S4 : DFFR_X1 port map( D => DATA2_I_30_port, CK => clk, RN => 
                           rst_BAR, Q => n4397, QN => n_1112);
   clk_r_REG2177_S4 : DFFS_X1 port map( D => DATA2_I_30_port, CK => clk, SN => 
                           rst_BAR, Q => n4396, QN => n_1113);
   clk_r_REG2254_S4 : DFFR_X1 port map( D => DATA2_I_29_port, CK => clk, RN => 
                           rst_BAR, Q => n4395, QN => n_1114);
   clk_r_REG2328_S4 : DFFS_X1 port map( D => DATA2_I_28_port, CK => clk, SN => 
                           rst_BAR, Q => n4394, QN => n_1115);
   clk_r_REG2643_S4 : DFFR_X1 port map( D => DATA2_I_24_port, CK => clk, RN => 
                           rst_BAR, Q => n4393, QN => n_1116);
   clk_r_REG295_S9 : DFFS_X1 port map( D => n1865, CK => clk, SN => n6056, Q =>
                           n7809, QN => n4392);
   clk_r_REG296_S10 : DFFR_X1 port map( D => n4392, CK => clk, RN => rst_BAR, Q
                           => n4391, QN => n7811);
   clk_r_REG297_S11 : DFFR_X1 port map( D => n4391, CK => clk, RN => rst_BAR, Q
                           => n4390, QN => n7812);
   clk_r_REG298_S12 : DFFR_X1 port map( D => n4390, CK => clk, RN => rst_BAR, Q
                           => n4389, QN => n_1117);
   clk_r_REG241_S8 : DFFS_X1 port map( D => n1867, CK => clk, SN => n6054, Q =>
                           n_1118, QN => n4388);
   clk_r_REG288_S9 : DFFR_X1 port map( D => n4388, CK => clk, RN => rst_BAR, Q 
                           => n4387, QN => n_1119);
   clk_r_REG289_S10 : DFFR_X1 port map( D => n4387, CK => clk, RN => n6055, Q 
                           => n4386, QN => n_1120);
   clk_r_REG290_S11 : DFFR_X1 port map( D => n4386, CK => clk, RN => n6056, Q 
                           => n4385, QN => n_1121);
   clk_r_REG335_S8 : DFFS_X1 port map( D => n1869, CK => clk, SN => rst_BAR, Q 
                           => n_1122, QN => n4384);
   clk_r_REG341_S9 : DFFR_X1 port map( D => n4384, CK => clk, RN => rst_BAR, Q 
                           => n4383, QN => n_1123);
   clk_r_REG342_S10 : DFFR_X1 port map( D => n4383, CK => clk, RN => n6056, Q 
                           => n4382, QN => n_1124);
   clk_r_REG343_S11 : DFFR_X1 port map( D => n4382, CK => clk, RN => rst_BAR, Q
                           => n4381, QN => n_1125);
   clk_r_REG180_S8 : DFFS_X1 port map( D => n1871, CK => clk, SN => rst_BAR, Q 
                           => n_1126, QN => n4380);
   clk_r_REG1716_S9 : DFFR_X1 port map( D => n4380, CK => clk, RN => rst_BAR, Q
                           => n4379, QN => n_1127);
   clk_r_REG1717_S10 : DFFR_X1 port map( D => n4379, CK => clk, RN => rst_BAR, 
                           Q => n4378, QN => n_1128);
   clk_r_REG1718_S11 : DFFR_X1 port map( D => n4378, CK => clk, RN => rst_BAR, 
                           Q => n4377, QN => n_1129);
   clk_r_REG408_S25 : DFFS_X1 port map( D => n1873, CK => clk, SN => rst_BAR, Q
                           => n_1130, QN => n4376);
   clk_r_REG415_S26 : DFFR_X1 port map( D => n4376, CK => clk, RN => rst_BAR, Q
                           => n4375, QN => n_1131);
   clk_r_REG416_S27 : DFFR_X1 port map( D => n4375, CK => clk, RN => rst_BAR, Q
                           => n4374, QN => n_1132);
   clk_r_REG417_S28 : DFFR_X1 port map( D => n4374, CK => clk, RN => rst_BAR, Q
                           => n4373, QN => n_1133);
   clk_r_REG32_S24 : DFFS_X1 port map( D => n1875, CK => clk, SN => rst_BAR, Q 
                           => n_1134, QN => n4372);
   clk_r_REG3014_S25 : DFFR_X1 port map( D => n4372, CK => clk, RN => rst_BAR, 
                           Q => n4371, QN => n_1135);
   clk_r_REG3015_S26 : DFFR_X1 port map( D => n4371, CK => clk, RN => rst_BAR, 
                           Q => n4370, QN => n_1136);
   clk_r_REG3016_S27 : DFFR_X1 port map( D => n4370, CK => clk, RN => rst_BAR, 
                           Q => n4369, QN => n_1137);
   clk_r_REG462_S7 : DFFS_X1 port map( D => n1877, CK => clk, SN => rst_BAR, Q 
                           => n_1138, QN => n4368);
   clk_r_REG463_S8 : DFFR_X1 port map( D => n4368, CK => clk, RN => rst_BAR, Q 
                           => n4367, QN => n_1139);
   clk_r_REG464_S9 : DFFR_X1 port map( D => n4367, CK => clk, RN => rst_BAR, Q 
                           => n4366, QN => n_1140);
   clk_r_REG465_S10 : DFFR_X1 port map( D => n4366, CK => clk, RN => rst_BAR, Q
                           => n4365, QN => n_1141);
   clk_r_REG139_S8 : DFFS_X1 port map( D => n1879, CK => clk, SN => rst_BAR, Q 
                           => n_1142, QN => n4364);
   clk_r_REG2089_S9 : DFFR_X1 port map( D => n4364, CK => clk, RN => rst_BAR, Q
                           => n4363, QN => n_1143);
   clk_r_REG2090_S10 : DFFR_X1 port map( D => n4363, CK => clk, RN => rst_BAR, 
                           Q => n4362, QN => n_1144);
   clk_r_REG2091_S11 : DFFR_X1 port map( D => n4362, CK => clk, RN => rst_BAR, 
                           Q => n4361, QN => n_1145);
   clk_r_REG429_S11 : DFFS_X1 port map( D => n1881, CK => clk, SN => rst_BAR, Q
                           => n_1146, QN => n4360);
   clk_r_REG450_S12 : DFFR_X1 port map( D => n4360, CK => clk, RN => n6056, Q 
                           => n4359, QN => n_1147);
   clk_r_REG451_S13 : DFFR_X1 port map( D => n4359, CK => clk, RN => rst_BAR, Q
                           => n4358, QN => n_1148);
   clk_r_REG452_S14 : DFFR_X1 port map( D => n4358, CK => clk, RN => rst_BAR, Q
                           => n4357, QN => n_1149);
   clk_r_REG375_S8 : DFFS_X1 port map( D => n1883, CK => clk, SN => rst_BAR, Q 
                           => n_1150, QN => n4356);
   clk_r_REG1215_S9 : DFFR_X1 port map( D => n4356, CK => clk, RN => rst_BAR, Q
                           => n4355, QN => n_1151);
   clk_r_REG1216_S10 : DFFR_X1 port map( D => n4355, CK => clk, RN => rst_BAR, 
                           Q => n4354, QN => n_1152);
   clk_r_REG1217_S11 : DFFR_X1 port map( D => n4354, CK => clk, RN => rst_BAR, 
                           Q => n4353, QN => n_1153);
   clk_r_REG473_S8 : DFFS_X1 port map( D => n1885, CK => clk, SN => rst_BAR, Q 
                           => n_1154, QN => n4352);
   clk_r_REG486_S9 : DFFR_X1 port map( D => n4352, CK => clk, RN => rst_BAR, Q 
                           => n4351, QN => n_1155);
   clk_r_REG487_S10 : DFFR_X1 port map( D => n4351, CK => clk, RN => n6055, Q 
                           => n4350, QN => n_1156);
   clk_r_REG488_S11 : DFFR_X1 port map( D => n4350, CK => clk, RN => rst_BAR, Q
                           => n4349, QN => n_1157);
   clk_r_REG323_S11 : DFFS_X1 port map( D => n1887, CK => clk, SN => rst_BAR, Q
                           => n_1158, QN => n4348);
   clk_r_REG1459_S12 : DFFR_X1 port map( D => n4348, CK => clk, RN => rst_BAR, 
                           Q => n4347, QN => n_1159);
   clk_r_REG1460_S13 : DFFR_X1 port map( D => n4347, CK => clk, RN => rst_BAR, 
                           Q => n4346, QN => n_1160);
   clk_r_REG1461_S14 : DFFR_X1 port map( D => n4346, CK => clk, RN => rst_BAR, 
                           Q => n4345, QN => n_1161);
   clk_r_REG1305_S11 : DFFS_X1 port map( D => n1889, CK => clk, SN => rst_BAR, 
                           Q => n_1162, QN => n4344);
   clk_r_REG1314_S12 : DFFR_X1 port map( D => n4344, CK => clk, RN => rst_BAR, 
                           Q => n4343, QN => n_1163);
   clk_r_REG1315_S13 : DFFR_X1 port map( D => n4343, CK => clk, RN => rst_BAR, 
                           Q => n4342, QN => n_1164);
   clk_r_REG1316_S14 : DFFR_X1 port map( D => n4342, CK => clk, RN => rst_BAR, 
                           Q => n4341, QN => n_1165);
   clk_r_REG1467_S11 : DFFS_X1 port map( D => n1891, CK => clk, SN => rst_BAR, 
                           Q => n_1166, QN => n4340);
   clk_r_REG1478_S12 : DFFR_X1 port map( D => n4340, CK => clk, RN => rst_BAR, 
                           Q => n4339, QN => n_1167);
   clk_r_REG1479_S13 : DFFR_X1 port map( D => n4339, CK => clk, RN => rst_BAR, 
                           Q => n4338, QN => n_1168);
   clk_r_REG1480_S14 : DFFR_X1 port map( D => n4338, CK => clk, RN => rst_BAR, 
                           Q => n4337, QN => n_1169);
   clk_r_REG21_S15 : DFFS_X1 port map( D => n1893, CK => clk, SN => rst_BAR, Q 
                           => n_1170, QN => n4336);
   clk_r_REG3030_S16 : DFFR_X1 port map( D => n4336, CK => clk, RN => rst_BAR, 
                           Q => n4335, QN => n_1171);
   clk_r_REG3031_S17 : DFFR_X1 port map( D => n4335, CK => clk, RN => rst_BAR, 
                           Q => n4334, QN => n_1172);
   clk_r_REG3032_S18 : DFFR_X1 port map( D => n4334, CK => clk, RN => rst_BAR, 
                           Q => n4333, QN => n_1173);
   clk_r_REG3106_S13 : DFFS_X1 port map( D => n1894, CK => clk, SN => rst_BAR, 
                           Q => n7743, QN => n4332);
   clk_r_REG3107_S14 : DFFR_X1 port map( D => n4332, CK => clk, RN => rst_BAR, 
                           Q => n4331, QN => n7744);
   clk_r_REG3108_S15 : DFFR_X1 port map( D => n4331, CK => clk, RN => rst_BAR, 
                           Q => n4330, QN => n7745);
   clk_r_REG3109_S16 : DFFR_X1 port map( D => n4330, CK => clk, RN => n6054, Q 
                           => n4329, QN => n7746);
   clk_r_REG1564_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, CK 
                           => clk, RN => n6056, Q => n4328, QN => n_1174);
   clk_r_REG1565_S5 : DFFR_X1 port map( D => n4328, CK => clk, RN => rst_BAR, Q
                           => n4327, QN => n_1175);
   clk_r_REG1566_S6 : DFFR_X1 port map( D => n4327, CK => clk, RN => rst_BAR, Q
                           => n4326, QN => n_1176);
   clk_r_REG1567_S7 : DFFR_X1 port map( D => n4326, CK => clk, RN => rst_BAR, Q
                           => n4325, QN => n_1177);
   clk_r_REG1568_S8 : DFFR_X1 port map( D => n4325, CK => clk, RN => rst_BAR, Q
                           => n_1178, QN => n6007);
   clk_r_REG1640_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, CK 
                           => clk, RN => rst_BAR, Q => n4323, QN => n_1179);
   clk_r_REG1641_S5 : DFFR_X1 port map( D => n4323, CK => clk, RN => rst_BAR, Q
                           => n4322, QN => n_1180);
   clk_r_REG1642_S6 : DFFR_X1 port map( D => n4322, CK => clk, RN => rst_BAR, Q
                           => n4321, QN => n_1181);
   clk_r_REG1643_S7 : DFFR_X1 port map( D => n4321, CK => clk, RN => rst_BAR, Q
                           => n4320, QN => n_1182);
   clk_r_REG1644_S8 : DFFR_X1 port map( D => n4320, CK => clk, RN => rst_BAR, Q
                           => n4319, QN => n_1183);
   clk_r_REG1386_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => n6055, Q => n4318, QN => n_1184);
   clk_r_REG1387_S5 : DFFR_X1 port map( D => n4318, CK => clk, RN => rst_BAR, Q
                           => n4317, QN => n_1185);
   clk_r_REG1388_S6 : DFFR_X1 port map( D => n4317, CK => clk, RN => rst_BAR, Q
                           => n4316, QN => n_1186);
   clk_r_REG1389_S7 : DFFR_X1 port map( D => n4316, CK => clk, RN => rst_BAR, Q
                           => n_1187, QN => n6006);
   clk_r_REG1390_S8 : DFFS_X1 port map( D => n6006, CK => clk, SN => rst_BAR, Q
                           => n_1188, QN => n4314);
   clk_r_REG1726_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, CK 
                           => clk, RN => rst_BAR, Q => n4313, QN => n_1189);
   clk_r_REG1727_S5 : DFFR_X1 port map( D => n4313, CK => clk, RN => rst_BAR, Q
                           => n4312, QN => n_1190);
   clk_r_REG1728_S6 : DFFR_X1 port map( D => n4312, CK => clk, RN => rst_BAR, Q
                           => n4311, QN => n_1191);
   clk_r_REG1729_S7 : DFFR_X1 port map( D => n4311, CK => clk, RN => rst_BAR, Q
                           => n4310, QN => n_1192);
   clk_r_REG1005_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => rst_BAR, Q => n4309, QN => n_1193);
   clk_r_REG1006_S5 : DFFR_X1 port map( D => n4309, CK => clk, RN => rst_BAR, Q
                           => n4308, QN => n_1194);
   clk_r_REG1007_S6 : DFFR_X1 port map( D => n4308, CK => clk, RN => rst_BAR, Q
                           => n_1195, QN => n6008);
   clk_r_REG1008_S7 : DFFS_X1 port map( D => n6008, CK => clk, SN => rst_BAR, Q
                           => n_1196, QN => n4306);
   clk_r_REG1080_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, CK 
                           => clk, RN => rst_BAR, Q => n4305, QN => n_1197);
   clk_r_REG1081_S5 : DFFR_X1 port map( D => n4305, CK => clk, RN => n6054, Q 
                           => n4304, QN => n_1198);
   clk_r_REG1082_S6 : DFFR_X1 port map( D => n4304, CK => clk, RN => rst_BAR, Q
                           => n4303, QN => n_1199);
   clk_r_REG751_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => n6054, Q => n4302, QN => n_1200);
   clk_r_REG752_S5 : DFFR_X1 port map( D => n4302, CK => clk, RN => rst_BAR, Q 
                           => n_1201, QN => n6009);
   clk_r_REG753_S6 : DFFS_X1 port map( D => n6009, CK => clk, SN => rst_BAR, Q 
                           => n_1202, QN => n4300);
   clk_r_REG829_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, CK 
                           => clk, RN => rst_BAR, Q => n4299, QN => n_1203);
   clk_r_REG830_S5 : DFFR_X1 port map( D => n4299, CK => clk, RN => rst_BAR, Q 
                           => n4298, QN => n_1204);
   clk_r_REG391_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => n6055, Q => n7769, QN => n6005);
   clk_r_REG392_S5 : DFFS_X1 port map( D => n6005, CK => clk, SN => rst_BAR, Q 
                           => n_1205, QN => n4296);
   clk_r_REG1227_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, CK 
                           => clk, RN => rst_BAR, Q => n4295, QN => n_1206);
   clk_r_REG526_S4 : DFFS_X1 port map( D => n1895, CK => clk, SN => rst_BAR, Q 
                           => n_1207, QN => n4294);
   clk_r_REG127_S4 : DFFS_X1 port map( D => DATA2_I_31_port, CK => clk, SN => 
                           n6056, Q => n4293, QN => n_1208);
   clk_r_REG530_S4 : DFFS_X1 port map( D => n5989, CK => clk, SN => rst_BAR, Q 
                           => n_1209, QN => n4292);
   clk_r_REG580_S3 : DFFS_X1 port map( D => n1949, CK => clk, SN => rst_BAR, Q 
                           => n_1210, QN => n4291);
   clk_r_REG579_S3 : DFFR_X1 port map( D => n1949, CK => clk, RN => rst_BAR, Q 
                           => n7740, QN => n4290);
   clk_r_REG284_S8 : DFFS_X1 port map( D => n1863, CK => clk, SN => rst_BAR, Q 
                           => n_1211, QN => n4288);
   clk_r_REG285_S9 : DFFR_X1 port map( D => n4288, CK => clk, RN => rst_BAR, Q 
                           => n4287, QN => n_1212);
   clk_r_REG286_S10 : DFFR_X1 port map( D => n4287, CK => clk, RN => rst_BAR, Q
                           => n4286, QN => n_1213);
   clk_r_REG287_S11 : DFFR_X1 port map( D => n4286, CK => clk, RN => rst_BAR, Q
                           => n4285, QN => n_1214);
   clk_r_REG911_S5 : DFFR_X1 port map( D => dataout_mul_4_port, CK => clk, RN 
                           => rst_BAR, Q => n4284, QN => n_1215);
   clk_r_REG912_S6 : DFFR_X1 port map( D => n4284, CK => clk, RN => n6054, Q =>
                           n4283, QN => n_1216);
   clk_r_REG913_S7 : DFFR_X1 port map( D => n4283, CK => clk, RN => rst_BAR, Q 
                           => n4282, QN => n_1217);
   clk_r_REG914_S8 : DFFR_X1 port map( D => n4282, CK => clk, RN => rst_BAR, Q 
                           => n4281, QN => n_1218);
   clk_r_REG915_S9 : DFFR_X1 port map( D => n4281, CK => clk, RN => rst_BAR, Q 
                           => n4280, QN => n_1219);
   clk_r_REG365_S5 : DFFR_X1 port map( D => dataout_mul_6_port, CK => clk, RN 
                           => rst_BAR, Q => n4279, QN => n_1220);
   clk_r_REG366_S6 : DFFR_X1 port map( D => n4279, CK => clk, RN => rst_BAR, Q 
                           => n4278, QN => n_1221);
   clk_r_REG367_S7 : DFFR_X1 port map( D => n4278, CK => clk, RN => rst_BAR, Q 
                           => n4277, QN => n_1222);
   clk_r_REG368_S8 : DFFR_X1 port map( D => n4277, CK => clk, RN => rst_BAR, Q 
                           => n4276, QN => n_1223);
   clk_r_REG369_S9 : DFFR_X1 port map( D => n4276, CK => clk, RN => rst_BAR, Q 
                           => n4275, QN => n_1224);
   clk_r_REG370_S10 : DFFS_X1 port map( D => n4275, CK => clk, SN => rst_BAR, Q
                           => n4274, QN => n_1225);
   clk_r_REG754_S16 : DFFR_X1 port map( D => dataout_mul_8_port, CK => clk, RN 
                           => rst_BAR, Q => n4273, QN => n_1226);
   clk_r_REG755_S17 : DFFR_X1 port map( D => n4273, CK => clk, RN => rst_BAR, Q
                           => n4272, QN => n_1227);
   clk_r_REG756_S18 : DFFR_X1 port map( D => n4272, CK => clk, RN => rst_BAR, Q
                           => n4271, QN => n_1228);
   clk_r_REG757_S19 : DFFR_X1 port map( D => n4271, CK => clk, RN => rst_BAR, Q
                           => n4270, QN => n_1229);
   clk_r_REG401_S17 : DFFR_X1 port map( D => dataout_mul_10_port, CK => clk, RN
                           => rst_BAR, Q => n4269, QN => n_1230);
   clk_r_REG402_S18 : DFFR_X1 port map( D => n4269, CK => clk, RN => rst_BAR, Q
                           => n4268, QN => n_1231);
   clk_r_REG403_S19 : DFFR_X1 port map( D => n4268, CK => clk, RN => rst_BAR, Q
                           => n4267, QN => n_1232);
   clk_r_REG404_S20 : DFFS_X1 port map( D => n4267, CK => clk, SN => rst_BAR, Q
                           => n4266, QN => n_1233);
   clk_r_REG396_S14 : DFFR_X1 port map( D => dataout_mul_12_port, CK => clk, RN
                           => rst_BAR, Q => n4265, QN => n_1234);
   clk_r_REG397_S15 : DFFR_X1 port map( D => n4265, CK => clk, RN => rst_BAR, Q
                           => n4264, QN => n_1235);
   clk_r_REG398_S16 : DFFS_X1 port map( D => n4264, CK => clk, SN => rst_BAR, Q
                           => n4263, QN => n_1236);
   clk_r_REG1469_S11 : DFFR_X1 port map( D => dataout_mul_2_port, CK => clk, RN
                           => rst_BAR, Q => n4262, QN => n_1237);
   clk_r_REG1470_S12 : DFFR_X1 port map( D => n4262, CK => clk, RN => rst_BAR, 
                           Q => n4261, QN => n_1238);
   clk_r_REG1471_S13 : DFFR_X1 port map( D => n4261, CK => clk, RN => n6056, Q 
                           => n4260, QN => n_1239);
   clk_r_REG1472_S14 : DFFR_X1 port map( D => n4260, CK => clk, RN => rst_BAR, 
                           Q => n4259, QN => n_1240);
   clk_r_REG1473_S15 : DFFR_X1 port map( D => n4259, CK => clk, RN => rst_BAR, 
                           Q => n4258, QN => n_1241);
   clk_r_REG1474_S16 : DFFR_X1 port map( D => n4258, CK => clk, RN => rst_BAR, 
                           Q => n4257, QN => n_1242);
   clk_r_REG539_S3 : DFFR_X1 port map( D => n1959, CK => clk, RN => rst_BAR, Q 
                           => n7758, QN => n4256);
   clk_r_REG658_S3 : DFFR_X1 port map( D => n7827, CK => clk, RN => rst_BAR, Q 
                           => n_1243, QN => n4255);
   clk_r_REG3460_S7 : DFFR_X1 port map( D => n7821, CK => clk, RN => rst_BAR, Q
                           => n_1244, QN => n4254);
   clk_r_REG743_S6 : DFFS_X1 port map( D => n2520_port, CK => clk, SN => 
                           rst_BAR, Q => n4253, QN => n_1245);
   clk_r_REG927_S3 : DFFR_X1 port map( D => n1968, CK => clk, RN => rst_BAR, Q 
                           => n7813, QN => n4252);
   clk_r_REG537_S3 : DFFR_X1 port map( D => n6023, CK => clk, RN => rst_BAR, Q 
                           => n7795, QN => n4251);
   clk_r_REG552_S3 : DFFR_X1 port map( D => n1961, CK => clk, RN => n6057, Q =>
                           n7750, QN => n4250);
   clk_r_REG560_S3 : DFFR_X1 port map( D => n1963, CK => clk, RN => rst_BAR, Q 
                           => n_1246, QN => n4249);
   clk_r_REG550_S3 : DFFR_X1 port map( D => n5987, CK => clk, RN => rst_BAR, Q 
                           => n7724, QN => n4248);
   clk_r_REG650_S39 : DFFR_X1 port map( D => n1084, CK => clk, RN => rst_BAR, Q
                           => n4247, QN => n_1247);
   clk_r_REG649_S39 : DFFS_X1 port map( D => n1084, CK => clk, SN => rst_BAR, Q
                           => n4246, QN => n_1248);
   clk_r_REG574_S3 : DFFR_X1 port map( D => n5985, CK => clk, RN => rst_BAR, Q 
                           => n7765, QN => n4244);
   clk_r_REG568_S3 : DFFR_X1 port map( D => n1948, CK => clk, RN => rst_BAR, Q 
                           => n7759, QN => n4243);
   clk_r_REG654_S3 : DFFR_X1 port map( D => n1559, CK => clk, RN => rst_BAR, Q 
                           => n4242, QN => n_1249);
   clk_r_REG638_S43 : DFFS_X1 port map( D => n1546, CK => clk, SN => rst_BAR, Q
                           => n4241, QN => n_1250);
   clk_r_REG657_S45 : DFFS_X1 port map( D => n1581, CK => clk, SN => rst_BAR, Q
                           => n4240, QN => n_1251);
   clk_r_REG672_S46 : DFFS_X1 port map( D => n1677, CK => clk, SN => rst_BAR, Q
                           => n4239, QN => n7791);
   clk_r_REG634_S45 : DFFS_X1 port map( D => n1556, CK => clk, SN => rst_BAR, Q
                           => n4238, QN => n_1252);
   clk_r_REG656_S46 : DFFS_X1 port map( D => n1594, CK => clk, SN => rst_BAR, Q
                           => n4237, QN => n_1253);
   clk_r_REG671_S48 : DFFS_X1 port map( D => n1129, CK => clk, SN => rst_BAR, Q
                           => n4236, QN => n_1254);
   clk_r_REG540_S3 : DFFR_X1 port map( D => n5996, CK => clk, RN => rst_BAR, Q 
                           => n7796, QN => n4235);
   clk_r_REG562_S3 : DFFR_X1 port map( D => n5991, CK => clk, RN => rst_BAR, Q 
                           => n7733, QN => n4234);
   clk_r_REG653_S3 : DFFS_X1 port map( D => n1680, CK => clk, SN => rst_BAR, Q 
                           => n4233, QN => n_1255);
   clk_r_REG627_S46 : DFFS_X1 port map( D => n1580, CK => clk, SN => n6055, Q 
                           => n4232, QN => n_1256);
   clk_r_REG661_S45 : DFFR_X1 port map( D => n1194, CK => clk, RN => rst_BAR, Q
                           => n4231, QN => n_1257);
   clk_r_REG659_S3 : DFFR_X1 port map( D => n1203, CK => clk, RN => rst_BAR, Q 
                           => n_1258, QN => n7793);
   clk_r_REG626_S48 : DFFS_X1 port map( D => n1593, CK => clk, SN => rst_BAR, Q
                           => n4229, QN => n_1259);
   clk_r_REG900_S10 : DFFS_X1 port map( D => n1322, CK => clk, SN => rst_BAR, Q
                           => n4228, QN => n_1260);
   clk_r_REG509_S7 : DFFR_X1 port map( D => n5990, CK => clk, RN => rst_BAR, Q 
                           => n_1261, QN => n4227);
   clk_r_REG503_S10 : DFFR_X1 port map( D => n1859, CK => clk, RN => rst_BAR, Q
                           => n_1262, QN => n4226);
   clk_r_REG499_S10 : DFFR_X1 port map( D => n1860, CK => clk, RN => rst_BAR, Q
                           => n_1263, QN => n4225);
   clk_r_REG3461_S7 : DFFR_X1 port map( D => n1900, CK => clk, RN => rst_BAR, Q
                           => n_1264, QN => n4224);
   clk_r_REG3458_S7 : DFFR_X1 port map( D => n1901, CK => clk, RN => rst_BAR, Q
                           => n_1265, QN => n4223);
   clk_r_REG533_S3 : DFFR_X1 port map( D => n1902, CK => clk, RN => rst_BAR, Q 
                           => n7798, QN => n4222);
   clk_r_REG3250_S3 : DFFR_X1 port map( D => n1896, CK => clk, RN => rst_BAR, Q
                           => n_1266, QN => n4221);
   clk_r_REG497_S7 : DFFR_X1 port map( D => n1319, CK => clk, RN => rst_BAR, Q 
                           => n4220, QN => n_1267);
   clk_r_REG929_S3 : DFFR_X1 port map( D => n5986, CK => clk, RN => rst_BAR, Q 
                           => n_1268, QN => n4219);
   clk_r_REG920_S3 : DFFR_X1 port map( D => n5999, CK => clk, RN => rst_BAR, Q 
                           => n7806, QN => n4218);
   clk_r_REG925_S3 : DFFS_X1 port map( D => n5998, CK => clk, SN => rst_BAR, Q 
                           => n_1269, QN => n4217);
   clk_r_REG1302_S4 : DFFR_X1 port map( D => n1862, CK => clk, RN => rst_BAR, Q
                           => n4216, QN => n_1270);
   clk_r_REG663_S48 : DFFS_X1 port map( D => n2008, CK => clk, SN => rst_BAR, Q
                           => n4215, QN => n_1271);
   clk_r_REG1874_S4 : DFFR_X1 port map( D => n1847, CK => clk, RN => rst_BAR, Q
                           => n_1272, QN => n4214);
   clk_r_REG169_S42 : DFFR_X1 port map( D => n6018, CK => clk, RN => rst_BAR, Q
                           => n_1273, QN => n4213);
   clk_r_REG2329_S48 : DFFS_X1 port map( D => n1986, CK => clk, SN => rst_BAR, 
                           Q => n4212, QN => n_1274);
   clk_r_REG2488_S45 : DFFS_X1 port map( D => n6015, CK => clk, SN => rst_BAR, 
                           Q => n_1275, QN => n4211);
   clk_r_REG2646_S42 : DFFS_X1 port map( D => n1845, CK => clk, SN => rst_BAR, 
                           Q => n_1276, QN => n4210);
   clk_r_REG2645_S42 : DFFR_X1 port map( D => n1845, CK => clk, RN => rst_BAR, 
                           Q => n_1277, QN => n4209);
   clk_r_REG2568_S43 : DFFS_X1 port map( D => n2070, CK => clk, SN => rst_BAR, 
                           Q => n4208, QN => n_1278);
   clk_r_REG2484_S45 : DFFS_X1 port map( D => n2058, CK => clk, SN => rst_BAR, 
                           Q => n4207, QN => n_1279);
   clk_r_REG166_S42 : DFFR_X1 port map( D => n1846, CK => clk, RN => n6056, Q 
                           => n7807, QN => n4206);
   clk_r_REG532_S3 : DFFS_X1 port map( D => n2690, CK => clk, SN => rst_BAR, Q 
                           => n4205, QN => n_1280);
   clk_r_REG2411_S3 : DFFR_X1 port map( D => n2669, CK => clk, RN => rst_BAR, Q
                           => n4204, QN => n_1281);
   clk_r_REG93_S46 : DFFR_X1 port map( D => n2594, CK => clk, RN => rst_BAR, Q 
                           => n4203, QN => n_1282);
   clk_r_REG2644_S42 : DFFR_X1 port map( D => n2082, CK => clk, RN => rst_BAR, 
                           Q => n4202, QN => n_1283);
   clk_r_REG301_S8 : DFFR_X1 port map( D => n1856, CK => clk, RN => rst_BAR, Q 
                           => n_1284, QN => n4201);
   clk_r_REG1391_S12 : DFFR_X1 port map( D => n2313, CK => clk, RN => rst_BAR, 
                           Q => n4200, QN => n_1285);
   clk_r_REG420_S24 : DFFR_X1 port map( D => n2379, CK => clk, RN => n6054, Q 
                           => n4199, QN => n_1286);
   clk_r_REG500_S10 : DFFS_X1 port map( D => n2401, CK => clk, SN => rst_BAR, Q
                           => n4198, QN => n_1287);
   clk_r_REG3_S4 : DFFR_X1 port map( D => dataout_mul_0_port, CK => clk, RN => 
                           rst_BAR, Q => n4197, QN => n_1288);
   clk_r_REG4_S5 : DFFR_X1 port map( D => n4197, CK => clk, RN => rst_BAR, Q =>
                           n4196, QN => n_1289);
   clk_r_REG5_S6 : DFFR_X1 port map( D => n4196, CK => clk, RN => n6057, Q => 
                           n4195, QN => n_1290);
   clk_r_REG6_S7 : DFFR_X1 port map( D => n4195, CK => clk, RN => n6054, Q => 
                           n4194, QN => n_1291);
   clk_r_REG7_S8 : DFFR_X1 port map( D => n4194, CK => clk, RN => rst_BAR, Q =>
                           n4193, QN => n_1292);
   clk_r_REG8_S9 : DFFR_X1 port map( D => n4193, CK => clk, RN => rst_BAR, Q =>
                           n4192, QN => n_1293);
   clk_r_REG527_S4 : DFFR_X1 port map( D => n6004, CK => clk, RN => rst_BAR, Q 
                           => n_1294, QN => n4191);
   clk_r_REG336_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_3_19_port, CK => clk, 
                           RN => rst_BAR, Q => n4190, QN => n_1295);
   clk_r_REG242_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_3_20_port, CK => clk, 
                           RN => n6055, Q => n4189, QN => n_1296);
   clk_r_REG262_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_3_21_port, CK => clk, 
                           RN => rst_BAR, Q => n4188, QN => n_1297);
   clk_r_REG276_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_3_22_port, CK => clk, 
                           RN => rst_BAR, Q => n4187, QN => n_1298);
   clk_r_REG264_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_22_port, CK => clk, 
                           RN => rst_BAR, Q => n4186, QN => n_1299);
   clk_r_REG265_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_23_port, CK => clk, 
                           RN => rst_BAR, Q => n4185, QN => n_1300);
   clk_r_REG278_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_4_24_port, CK => clk, 
                           RN => rst_BAR, Q => n4184, QN => n_1301);
   clk_r_REG267_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_24_port, CK => clk, 
                           RN => rst_BAR, Q => n4183, QN => n_1302);
   clk_r_REG268_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_25_port, CK => clk, 
                           RN => rst_BAR, Q => n4182, QN => n_1303);
   clk_r_REG280_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_5_26_port, CK => clk, 
                           RN => rst_BAR, Q => n4181, QN => n_1304);
   clk_r_REG270_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_26_port, CK => clk, 
                           RN => rst_BAR, Q => n4180, QN => n_1305);
   clk_r_REG271_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_27_port, CK => clk, 
                           RN => rst_BAR, Q => n4179, QN => n_1306);
   clk_r_REG282_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_6_28_port, CK => clk, 
                           RN => rst_BAR, Q => n4178, QN => n_1307);
   clk_r_REG272_S12 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_28_port, CK => clk, 
                           RN => rst_BAR, Q => n4177, QN => n_1308);
   clk_r_REG273_S12 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_29_port, CK => clk, 
                           RN => rst_BAR, Q => n4176, QN => n_1309);
   clk_r_REG283_S12 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_7_30_port, CK => clk, 
                           RN => rst_BAR, Q => n4175, QN => n_1310);
   clk_r_REG3020_S15 : DFFS_X1 port map( D => n1892, CK => clk, SN => rst_BAR, 
                           Q => n_1311, QN => n4174);
   clk_r_REG3027_S16 : DFFR_X1 port map( D => n4174, CK => clk, RN => rst_BAR, 
                           Q => n4173, QN => n_1312);
   clk_r_REG3028_S17 : DFFR_X1 port map( D => n4173, CK => clk, RN => rst_BAR, 
                           Q => n4172, QN => n_1313);
   clk_r_REG3029_S18 : DFFR_X1 port map( D => n4172, CK => clk, RN => rst_BAR, 
                           Q => n4171, QN => n_1314);
   clk_r_REG1468_S11 : DFFS_X1 port map( D => n1890, CK => clk, SN => rst_BAR, 
                           Q => n_1315, QN => n4170);
   clk_r_REG1475_S12 : DFFR_X1 port map( D => n4170, CK => clk, RN => rst_BAR, 
                           Q => n4169, QN => n_1316);
   clk_r_REG1476_S13 : DFFR_X1 port map( D => n4169, CK => clk, RN => rst_BAR, 
                           Q => n4168, QN => n_1317);
   clk_r_REG1477_S14 : DFFR_X1 port map( D => n4168, CK => clk, RN => n6056, Q 
                           => n4167, QN => n_1318);
   clk_r_REG1306_S11 : DFFS_X1 port map( D => n1888, CK => clk, SN => rst_BAR, 
                           Q => n_1319, QN => n4166);
   clk_r_REG1307_S12 : DFFR_X1 port map( D => n4166, CK => clk, RN => rst_BAR, 
                           Q => n4165, QN => n_1320);
   clk_r_REG1308_S13 : DFFR_X1 port map( D => n4165, CK => clk, RN => rst_BAR, 
                           Q => n4164, QN => n_1321);
   clk_r_REG1309_S14 : DFFR_X1 port map( D => n4164, CK => clk, RN => rst_BAR, 
                           Q => n4163, QN => n_1322);
   clk_r_REG1310_S11 : DFFS_X1 port map( D => n1886, CK => clk, SN => rst_BAR, 
                           Q => n_1323, QN => n4162);
   clk_r_REG1311_S12 : DFFR_X1 port map( D => n4162, CK => clk, RN => rst_BAR, 
                           Q => n4161, QN => n_1324);
   clk_r_REG1312_S13 : DFFR_X1 port map( D => n4161, CK => clk, RN => n6054, Q 
                           => n4160, QN => n_1325);
   clk_r_REG1313_S14 : DFFR_X1 port map( D => n4160, CK => clk, RN => rst_BAR, 
                           Q => n4159, QN => n_1326);
   clk_r_REG474_S8 : DFFS_X1 port map( D => n1884, CK => clk, SN => rst_BAR, Q 
                           => n_1327, QN => n4158);
   clk_r_REG483_S9 : DFFR_X1 port map( D => n4158, CK => clk, RN => rst_BAR, Q 
                           => n4157, QN => n_1328);
   clk_r_REG484_S10 : DFFR_X1 port map( D => n4157, CK => clk, RN => rst_BAR, Q
                           => n4156, QN => n_1329);
   clk_r_REG485_S11 : DFFR_X1 port map( D => n4156, CK => clk, RN => rst_BAR, Q
                           => n4155, QN => n_1330);
   clk_r_REG376_S8 : DFFS_X1 port map( D => n1882, CK => clk, SN => rst_BAR, Q 
                           => n_1331, QN => n4154);
   clk_r_REG1212_S9 : DFFR_X1 port map( D => n4154, CK => clk, RN => n6056, Q 
                           => n4153, QN => n_1332);
   clk_r_REG1213_S10 : DFFR_X1 port map( D => n4153, CK => clk, RN => rst_BAR, 
                           Q => n4152, QN => n_1333);
   clk_r_REG1214_S11 : DFFR_X1 port map( D => n4152, CK => clk, RN => rst_BAR, 
                           Q => n4151, QN => n_1334);
   clk_r_REG430_S8 : DFFS_X1 port map( D => n1880, CK => clk, SN => rst_BAR, Q 
                           => n_1335, QN => n4150);
   clk_r_REG435_S9 : DFFR_X1 port map( D => n4150, CK => clk, RN => n6055, Q =>
                           n4149, QN => n_1336);
   clk_r_REG436_S10 : DFFR_X1 port map( D => n4149, CK => clk, RN => rst_BAR, Q
                           => n4148, QN => n_1337);
   clk_r_REG437_S11 : DFFR_X1 port map( D => n4148, CK => clk, RN => rst_BAR, Q
                           => n4147, QN => n_1338);
   clk_r_REG438_S8 : DFFS_X1 port map( D => n1878, CK => clk, SN => rst_BAR, Q 
                           => n_1339, QN => n4146);
   clk_r_REG439_S9 : DFFR_X1 port map( D => n4146, CK => clk, RN => rst_BAR, Q 
                           => n4145, QN => n_1340);
   clk_r_REG440_S10 : DFFR_X1 port map( D => n4145, CK => clk, RN => rst_BAR, Q
                           => n4144, QN => n_1341);
   clk_r_REG441_S11 : DFFR_X1 port map( D => n4144, CK => clk, RN => rst_BAR, Q
                           => n4143, QN => n_1342);
   clk_r_REG442_S8 : DFFS_X1 port map( D => n1876, CK => clk, SN => rst_BAR, Q 
                           => n_1343, QN => n4142);
   clk_r_REG443_S9 : DFFR_X1 port map( D => n4142, CK => clk, RN => rst_BAR, Q 
                           => n4141, QN => n_1344);
   clk_r_REG444_S10 : DFFR_X1 port map( D => n4141, CK => clk, RN => n6057, Q 
                           => n4140, QN => n_1345);
   clk_r_REG445_S11 : DFFR_X1 port map( D => n4140, CK => clk, RN => rst_BAR, Q
                           => n4139, QN => n_1346);
   clk_r_REG446_S8 : DFFS_X1 port map( D => n1874, CK => clk, SN => rst_BAR, Q 
                           => n_1347, QN => n4138);
   clk_r_REG447_S9 : DFFR_X1 port map( D => n4138, CK => clk, RN => rst_BAR, Q 
                           => n4137, QN => n_1348);
   clk_r_REG448_S10 : DFFR_X1 port map( D => n4137, CK => clk, RN => rst_BAR, Q
                           => n4136, QN => n_1349);
   clk_r_REG449_S11 : DFFR_X1 port map( D => n4136, CK => clk, RN => rst_BAR, Q
                           => n4135, QN => n_1350);
   clk_r_REG409_S25 : DFFS_X1 port map( D => n1872, CK => clk, SN => rst_BAR, Q
                           => n_1351, QN => n4134);
   clk_r_REG412_S26 : DFFR_X1 port map( D => n4134, CK => clk, RN => rst_BAR, Q
                           => n4133, QN => n_1352);
   clk_r_REG413_S27 : DFFR_X1 port map( D => n4133, CK => clk, RN => rst_BAR, Q
                           => n4132, QN => n_1353);
   clk_r_REG414_S28 : DFFR_X1 port map( D => n4132, CK => clk, RN => rst_BAR, Q
                           => n4131, QN => n_1354);
   clk_r_REG229_S8 : DFFS_X1 port map( D => n1870, CK => clk, SN => rst_BAR, Q 
                           => n_1355, QN => n4130);
   clk_r_REG1713_S9 : DFFR_X1 port map( D => n4130, CK => clk, RN => rst_BAR, Q
                           => n4129, QN => n_1356);
   clk_r_REG1714_S10 : DFFR_X1 port map( D => n4129, CK => clk, RN => rst_BAR, 
                           Q => n4128, QN => n_1357);
   clk_r_REG1715_S11 : DFFR_X1 port map( D => n4128, CK => clk, RN => rst_BAR, 
                           Q => n4127, QN => n_1358);
   clk_r_REG337_S8 : DFFS_X1 port map( D => n1868, CK => clk, SN => rst_BAR, Q 
                           => n_1359, QN => n4126);
   clk_r_REG338_S9 : DFFR_X1 port map( D => n4126, CK => clk, RN => rst_BAR, Q 
                           => n4125, QN => n_1360);
   clk_r_REG339_S10 : DFFR_X1 port map( D => n4125, CK => clk, RN => rst_BAR, Q
                           => n4124, QN => n_1361);
   clk_r_REG340_S11 : DFFR_X1 port map( D => n4124, CK => clk, RN => n6057, Q 
                           => n4123, QN => n_1362);
   clk_r_REG243_S8 : DFFS_X1 port map( D => n1866, CK => clk, SN => rst_BAR, Q 
                           => n_1363, QN => n4122);
   clk_r_REG263_S9 : DFFR_X1 port map( D => n4122, CK => clk, RN => n6057, Q =>
                           n4121, QN => n_1364);
   clk_r_REG266_S10 : DFFR_X1 port map( D => n4121, CK => clk, RN => rst_BAR, Q
                           => n4120, QN => n_1365);
   clk_r_REG269_S11 : DFFR_X1 port map( D => n4120, CK => clk, RN => rst_BAR, Q
                           => n4119, QN => n_1366);
   clk_r_REG274_S8 : DFFS_X1 port map( D => n1864, CK => clk, SN => rst_BAR, Q 
                           => n_1367, QN => n4118);
   clk_r_REG277_S9 : DFFR_X1 port map( D => n4118, CK => clk, RN => rst_BAR, Q 
                           => n4117, QN => n_1368);
   clk_r_REG279_S10 : DFFR_X1 port map( D => n4117, CK => clk, RN => rst_BAR, Q
                           => n4116, QN => n_1369);
   clk_r_REG281_S11 : DFFR_X1 port map( D => n4116, CK => clk, RN => rst_BAR, Q
                           => n4115, QN => n_1370);
   clk_r_REG542_S3 : DFFS_X1 port map( D => n6003, CK => clk, SN => rst_BAR, Q 
                           => n7802, QN => n4114);
   clk_r_REG932_S3 : DFFR_X1 port map( D => n1966, CK => clk, RN => rst_BAR, Q 
                           => n7728, QN => n4113);
   clk_r_REG910_S4 : DFFS_X1 port map( D => n2773, CK => clk, SN => rst_BAR, Q 
                           => n4111, QN => n_1371);
   clk_r_REG564_S3 : DFFS_X1 port map( D => n1962, CK => clk, SN => rst_BAR, Q 
                           => n7751, QN => n4110);
   clk_r_REG607_S3 : DFFS_X1 port map( D => n1952, CK => clk, SN => rst_BAR, Q 
                           => n_1372, QN => n4109);
   clk_r_REG606_S3 : DFFR_X1 port map( D => n1952, CK => clk, RN => rst_BAR, Q 
                           => n_1373, QN => n4108);
   clk_r_REG652_S3 : DFFR_X1 port map( D => n7828, CK => clk, RN => n6057, Q =>
                           n_1374, QN => n4107);
   clk_r_REG619_S3 : DFFR_X1 port map( D => n7826, CK => clk, RN => rst_BAR, Q 
                           => n_1375, QN => n4106);
   clk_r_REG667_S3 : DFFR_X1 port map( D => n7824, CK => clk, RN => rst_BAR, Q 
                           => n7780, QN => n_1376);
   clk_r_REG647_S41 : DFFS_X1 port map( D => n1105, CK => clk, SN => n6057, Q 
                           => n4104, QN => n7783);
   clk_r_REG586_S3 : DFFS_X1 port map( D => n1950, CK => clk, SN => rst_BAR, Q 
                           => n_1377, QN => n4103);
   clk_r_REG572_S3 : DFFR_X1 port map( D => n5997, CK => clk, RN => rst_BAR, Q 
                           => n7756, QN => n4101);
   clk_r_REG641_S35 : DFFR_X1 port map( D => n1120, CK => clk, RN => rst_BAR, Q
                           => n4100, QN => n_1378);
   clk_r_REG316_S8 : DFFS_X1 port map( D => n1178, CK => clk, SN => rst_BAR, Q 
                           => n4099, QN => n_1379);
   clk_r_REG555_S3 : DFFR_X1 port map( D => n6002, CK => clk, RN => n6057, Q =>
                           n7800, QN => n4098);
   clk_r_REG916_S10 : DFFS_X1 port map( D => n1429, CK => clk, SN => rst_BAR, Q
                           => n4097, QN => n_1380);
   clk_r_REG1219_S7 : DFFS_X1 port map( D => n1353, CK => clk, SN => rst_BAR, Q
                           => n4096, QN => n_1381);
   clk_r_REG831_S7 : DFFR_X1 port map( D => n1858, CK => clk, RN => rst_BAR, Q 
                           => n_1382, QN => n4095);
   clk_r_REG553_S3 : DFFR_X1 port map( D => n6001, CK => clk, RN => rst_BAR, Q 
                           => n_1383, QN => n4094);
   clk_r_REG468_S6 : DFFR_X1 port map( D => n1403, CK => clk, RN => rst_BAR, Q 
                           => n4093, QN => n7789);
   clk_r_REG919_S3 : DFFS_X1 port map( D => n1969, CK => clk, SN => rst_BAR, Q 
                           => n7729, QN => n4092);
   clk_r_REG923_S3 : DFFR_X1 port map( D => n5988, CK => clk, RN => rst_BAR, Q 
                           => n_1384, QN => n4091);
   clk_r_REG2799_S36 : DFFR_X1 port map( D => n1852, CK => clk, RN => rst_BAR, 
                           Q => n_1385, QN => n4090);
   clk_r_REG2940_S32 : DFFR_X1 port map( D => n1854, CK => clk, RN => rst_BAR, 
                           Q => n_1386, QN => n4089);
   clk_r_REG1645_S7 : DFFS_X1 port map( D => n2323, CK => clk, SN => rst_BAR, Q
                           => n4088, QN => n_1387);
   clk_r_REG2723_S38 : DFFR_X1 port map( D => n1850, CK => clk, RN => n6054, Q 
                           => n_1388, QN => n4087);
   clk_r_REG68_S39 : DFFR_X1 port map( D => n1849, CK => clk, RN => rst_BAR, Q 
                           => n_1389, QN => n4086);
   clk_r_REG2565_S43 : DFFS_X1 port map( D => n1844, CK => clk, SN => rst_BAR, 
                           Q => n_1390, QN => n4085);
   clk_r_REG2486_S45 : DFFS_X1 port map( D => n1842, CK => clk, SN => rst_BAR, 
                           Q => n_1391, QN => n4084);
   clk_r_REG2408_S46 : DFFS_X1 port map( D => n1841, CK => clk, SN => rst_BAR, 
                           Q => n_1392, QN => n4083);
   clk_r_REG2407_S46 : DFFR_X1 port map( D => n1841, CK => clk, RN => rst_BAR, 
                           Q => n_1393, QN => n4082);
   clk_r_REG2566_S42 : DFFR_X1 port map( D => n6017, CK => clk, RN => rst_BAR, 
                           Q => n_1394, QN => n4081);
   clk_r_REG2485_S45 : DFFR_X1 port map( D => n2031, CK => clk, RN => rst_BAR, 
                           Q => n7810, QN => n5993);
   clk_r_REG1482_S10 : DFFR_X1 port map( D => n1976, CK => clk, RN => rst_BAR, 
                           Q => n4079, QN => n_1395);
   clk_r_REG2412_S3 : DFFR_X1 port map( D => n2028, CK => clk, RN => rst_BAR, Q
                           => n4078, QN => n_1396);
   clk_r_REG96_S46 : DFFR_X1 port map( D => n2026, CK => clk, RN => n6055, Q =>
                           n4077, QN => n_1397);
   clk_r_REG2570_S3 : DFFS_X1 port map( D => n2521_port, CK => clk, SN => 
                           rst_BAR, Q => n4076, QN => n_1398);
   clk_r_REG167_S42 : DFFS_X1 port map( D => n2084, CK => clk, SN => n6054, Q 
                           => n4075, QN => n_1399);
   clk_r_REG165_S42 : DFFR_X1 port map( D => n2097, CK => clk, RN => rst_BAR, Q
                           => n4074, QN => n_1400);
   clk_r_REG1802_S3 : DFFS_X1 port map( D => n2094, CK => clk, SN => rst_BAR, Q
                           => n4073, QN => n_1401);
   clk_r_REG1951_S3 : DFFS_X1 port map( D => n2144, CK => clk, SN => rst_BAR, Q
                           => n4072, QN => n_1402);
   clk_r_REG2725_S3 : DFFR_X1 port map( D => n2161, CK => clk, RN => n6054, Q 
                           => n4071, QN => n_1403);
   clk_r_REG535_S3 : DFFR_X1 port map( D => n2204, CK => clk, RN => rst_BAR, Q 
                           => n4070, QN => n_1404);
   clk_r_REG16_S12 : DFFS_X1 port map( D => n2210, CK => clk, SN => rst_BAR, Q 
                           => n4069, QN => n_1405);
   clk_r_REG57_S36 : DFFS_X1 port map( D => n2219, CK => clk, SN => rst_BAR, Q 
                           => n4068, QN => n_1406);
   clk_r_REG2872_S3 : DFFR_X1 port map( D => n2245, CK => clk, RN => rst_BAR, Q
                           => n4067, QN => n_1407);
   clk_r_REG2949_S3 : DFFR_X1 port map( D => n2275, CK => clk, RN => rst_BAR, Q
                           => n4066, QN => n_1408);
   clk_r_REG346_S7 : DFFR_X1 port map( D => n2321, CK => clk, RN => rst_BAR, Q 
                           => n4065, QN => n_1409);
   clk_r_REG1392_S3 : DFFR_X1 port map( D => n2338, CK => clk, RN => rst_BAR, Q
                           => n4064, QN => n_1410);
   clk_r_REG344_S7 : DFFR_X1 port map( D => n2337, CK => clk, RN => rst_BAR, Q 
                           => n4063, QN => n_1411);
   clk_r_REG329_S16 : DFFS_X1 port map( D => n2381, CK => clk, SN => rst_BAR, Q
                           => n4062, QN => n_1412);
   clk_r_REG504_S10 : DFFS_X1 port map( D => n2407, CK => clk, SN => rst_BAR, Q
                           => n4061, QN => n_1413);
   clk_r_REG14_S12 : DFFS_X1 port map( D => n2694, CK => clk, SN => n6057, Q =>
                           n4060, QN => n_1414);
   clk_r_REG95_S46 : DFFR_X1 port map( D => n2671, CK => clk, RN => rst_BAR, Q 
                           => n4059, QN => n_1415);
   clk_r_REG94_S46 : DFFS_X1 port map( D => n2671, CK => clk, SN => rst_BAR, Q 
                           => n4058, QN => n_1416);
   clk_r_REG87_S45 : DFFR_X1 port map( D => n2595, CK => clk, RN => rst_BAR, Q 
                           => n4057, QN => n_1417);
   clk_r_REG899_S7 : DFFS_X1 port map( D => n2622, CK => clk, SN => rst_BAR, Q 
                           => n4056, QN => n_1418);
   clk_r_REG364_S4 : DFFS_X1 port map( D => n2806, CK => clk, SN => rst_BAR, Q 
                           => n4055, QN => n_1419);
   clk_r_REG363_S4 : DFFS_X1 port map( D => n2808, CK => clk, SN => rst_BAR, Q 
                           => n4054, QN => n_1420);
   clk_r_REG1293_S15 : DFFR_X1 port map( D => dataout_mul_3_port, CK => clk, RN
                           => rst_BAR, Q => n4053, QN => n_1421);
   clk_r_REG1294_S16 : DFFR_X1 port map( D => n4053, CK => clk, RN => rst_BAR, 
                           Q => n4052, QN => n_1422);
   clk_r_REG1295_S17 : DFFR_X1 port map( D => n4052, CK => clk, RN => n6056, Q 
                           => n4051, QN => n_1423);
   clk_r_REG1296_S18 : DFFR_X1 port map( D => n4051, CK => clk, RN => rst_BAR, 
                           Q => n4050, QN => n_1424);
   clk_r_REG1297_S19 : DFFR_X1 port map( D => n4050, CK => clk, RN => rst_BAR, 
                           Q => n4049, QN => n_1425);
   clk_r_REG1298_S20 : DFFR_X1 port map( D => n4049, CK => clk, RN => rst_BAR, 
                           Q => n4048, QN => n_1426);
   clk_r_REG1292_S4 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_4_port, CK => clk, 
                           RN => rst_BAR, Q => n_1427, QN => n7771);
   clk_r_REG476_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CK => clk, 
                           RN => rst_BAR, Q => n4046, QN => n_1428);
   clk_r_REG475_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CK => clk, 
                           RN => rst_BAR, Q => n4045, QN => n_1429);
   clk_r_REG377_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CK => clk, 
                           RN => rst_BAR, Q => n4044, QN => n_1430);
   clk_r_REG431_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CK => clk, 
                           RN => rst_BAR, Q => n4043, QN => n_1431);
   clk_r_REG433_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CK => clk, 
                           RN => rst_BAR, Q => n4042, QN => n_1432);
   clk_r_REG434_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CK => clk, 
                           RN => rst_BAR, Q => n4041, QN => n_1433);
   clk_r_REG411_S25 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CK => clk, 
                           RN => rst_BAR, Q => n4040, QN => n_1434);
   clk_r_REG410_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CK => clk, 
                           RN => rst_BAR, Q => n4039, QN => n_1435);
   clk_r_REG230_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CK => clk, 
                           RN => rst_BAR, Q => n4038, QN => n_1436);
   clk_r_REG261_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CK => clk, 
                           RN => rst_BAR, Q => n4037, QN => n_1437);
   clk_r_REG244_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CK => clk, 
                           RN => rst_BAR, Q => n4036, QN => n_1438);
   clk_r_REG257_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CK => clk, 
                           RN => rst_BAR, Q => n4035, QN => n_1439);
   clk_r_REG258_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CK => clk, 
                           RN => n6057, Q => n4034, QN => n_1440);
   clk_r_REG259_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CK => clk, 
                           RN => rst_BAR, Q => n4033, QN => n_1441);
   clk_r_REG260_S9 : DFFR_X1 port map( D => n4033, CK => clk, RN => rst_BAR, Q 
                           => n4032, QN => n_1442);
   clk_r_REG477_S9 : DFFR_X1 port map( D => dataout_mul_5_port, CK => clk, RN 
                           => n6054, Q => n4031, QN => n_1443);
   clk_r_REG478_S10 : DFFR_X1 port map( D => n4031, CK => clk, RN => rst_BAR, Q
                           => n4030, QN => n_1444);
   clk_r_REG479_S11 : DFFR_X1 port map( D => n4030, CK => clk, RN => n6055, Q 
                           => n4029, QN => n_1445);
   clk_r_REG480_S12 : DFFR_X1 port map( D => n4029, CK => clk, RN => rst_BAR, Q
                           => n4028, QN => n_1446);
   clk_r_REG481_S13 : DFFR_X1 port map( D => n4028, CK => clk, RN => rst_BAR, Q
                           => n4027, QN => n_1447);
   clk_r_REG255_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CK => clk, RN => rst_BAR, Q => n4026, QN => n_1448);
   clk_r_REG256_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CK => clk, 
                           RN => rst_BAR, Q => n4025, QN => n_1449);
   clk_r_REG378_S5 : DFFR_X1 port map( D => dataout_mul_7_port, CK => clk, RN 
                           => rst_BAR, Q => n4024, QN => n_1450);
   clk_r_REG379_S6 : DFFR_X1 port map( D => n4024, CK => clk, RN => rst_BAR, Q 
                           => n4023, QN => n_1451);
   clk_r_REG380_S7 : DFFR_X1 port map( D => n4023, CK => clk, RN => rst_BAR, Q 
                           => n4022, QN => n_1452);
   clk_r_REG381_S8 : DFFR_X1 port map( D => n4022, CK => clk, RN => rst_BAR, Q 
                           => n4021, QN => n_1453);
   clk_r_REG382_S9 : DFFR_X1 port map( D => n4021, CK => clk, RN => rst_BAR, Q 
                           => n4020, QN => n_1454);
   clk_r_REG22_S15 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_8_port, CK => clk, 
                           RN => rst_BAR, Q => n_1455, QN => n7774);
   clk_r_REG432_S15 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CK => clk, 
                           RN => rst_BAR, Q => n4018, QN => n_1456);
   clk_r_REG399_S5 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CK => clk, 
                           RN => rst_BAR, Q => n4017, QN => n_1457);
   clk_r_REG324_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CK => clk, 
                           RN => rst_BAR, Q => n4016, QN => n_1458);
   clk_r_REG393_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CK => clk, 
                           RN => n6054, Q => n4015, QN => n_1459);
   clk_r_REG231_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CK => clk, 
                           RN => n6054, Q => n4014, QN => n_1460);
   clk_r_REG140_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CK => clk, 
                           RN => rst_BAR, Q => n4013, QN => n_1461);
   clk_r_REG245_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CK => clk, 
                           RN => rst_BAR, Q => n4012, QN => n_1462);
   clk_r_REG33_S24 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CK => clk, 
                           RN => rst_BAR, Q => n4011, QN => n_1463);
   clk_r_REG249_S24 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CK => clk, 
                           RN => rst_BAR, Q => n4010, QN => n_1464);
   clk_r_REG181_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CK => clk, RN => rst_BAR, Q => n4009, QN => n_1465);
   clk_r_REG182_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CK => clk, 
                           RN => rst_BAR, Q => n4008, QN => n_1466);
   clk_r_REG228_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CK => clk, 
                           RN => rst_BAR, Q => n4007, QN => n_1467);
   clk_r_REG23_S16 : DFFR_X1 port map( D => dataout_mul_9_port, CK => clk, RN 
                           => rst_BAR, Q => n4006, QN => n_1468);
   clk_r_REG24_S17 : DFFR_X1 port map( D => n4006, CK => clk, RN => n6055, Q =>
                           n4005, QN => n_1469);
   clk_r_REG25_S18 : DFFR_X1 port map( D => n4005, CK => clk, RN => rst_BAR, Q 
                           => n4004, QN => n_1470);
   clk_r_REG26_S19 : DFFR_X1 port map( D => n4004, CK => clk, RN => rst_BAR, Q 
                           => n4003, QN => n_1471);
   clk_r_REG400_S16 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_10_port, CK => clk, 
                           RN => rst_BAR, Q => n_1472, QN => n7775);
   clk_r_REG325_S12 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CK => clk, 
                           RN => n6056, Q => n4001, QN => n_1473);
   clk_r_REG394_S12 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CK => clk, 
                           RN => rst_BAR, Q => n4000, QN => n_1474);
   clk_r_REG232_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CK => clk, 
                           RN => rst_BAR, Q => n3999, QN => n_1475);
   clk_r_REG141_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CK => clk, 
                           RN => rst_BAR, Q => n3998, QN => n_1476);
   clk_r_REG246_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CK => clk, 
                           RN => rst_BAR, Q => n3997, QN => n_1477);
   clk_r_REG34_S25 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CK => clk, 
                           RN => rst_BAR, Q => n3996, QN => n_1478);
   clk_r_REG250_S25 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CK => clk, 
                           RN => n6054, Q => n3995, QN => n_1479);
   clk_r_REG183_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CK => clk, 
                           RN => rst_BAR, Q => n3994, QN => n_1480);
   clk_r_REG223_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CK => clk, 
                           RN => rst_BAR, Q => n3993, QN => n_1481);
   clk_r_REG224_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CK => clk, 
                           RN => rst_BAR, Q => n3992, QN => n_1482);
   clk_r_REG225_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CK => clk, RN => rst_BAR, Q => n3991, QN => n_1483);
   clk_r_REG226_S9 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CK => clk, 
                           RN => rst_BAR, Q => n3990, QN => n_1484);
   clk_r_REG227_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CK => clk, 
                           RN => n6057, Q => n3989, QN => n_1485);
   clk_r_REG326_S13 : DFFR_X1 port map( D => dataout_mul_11_port, CK => clk, RN
                           => n6057, Q => n3988, QN => n_1486);
   clk_r_REG327_S14 : DFFR_X1 port map( D => n3988, CK => clk, RN => rst_BAR, Q
                           => n3987, QN => n_1487);
   clk_r_REG328_S15 : DFFR_X1 port map( D => n3987, CK => clk, RN => rst_BAR, Q
                           => n3986, QN => n_1488);
   clk_r_REG395_S13 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_12_port, CK => clk, 
                           RN => rst_BAR, Q => n_1489, QN => n7776);
   clk_r_REG233_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CK => clk, 
                           RN => rst_BAR, Q => n3984, QN => n_1490);
   clk_r_REG142_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CK => clk, 
                           RN => rst_BAR, Q => n3983, QN => n_1491);
   clk_r_REG247_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CK => clk, 
                           RN => rst_BAR, Q => n3982, QN => n_1492);
   clk_r_REG35_S26 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CK => clk, 
                           RN => rst_BAR, Q => n3981, QN => n_1493);
   clk_r_REG251_S26 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CK => clk, 
                           RN => rst_BAR, Q => n3980, QN => n_1494);
   clk_r_REG184_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CK => clk, 
                           RN => rst_BAR, Q => n3979, QN => n_1495);
   clk_r_REG216_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CK => clk, 
                           RN => rst_BAR, Q => n3978, QN => n_1496);
   clk_r_REG217_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CK => clk, 
                           RN => rst_BAR, Q => n3977, QN => n_1497);
   clk_r_REG218_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CK => clk, 
                           RN => rst_BAR, Q => n3976, QN => n_1498);
   clk_r_REG219_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CK => clk, 
                           RN => n6055, Q => n3975, QN => n_1499);
   clk_r_REG220_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CK => clk, RN => rst_BAR, Q => n3974, QN => n_1500);
   clk_r_REG221_S10 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CK => clk, 
                           RN => rst_BAR, Q => n3973, QN => n_1501);
   clk_r_REG222_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CK => clk, 
                           RN => n6057, Q => n3972, QN => n_1502);
   clk_r_REG234_S12 : DFFR_X1 port map( D => dataout_mul_13_port, CK => clk, RN
                           => n6057, Q => n3971, QN => n_1503);
   clk_r_REG235_S13 : DFFR_X1 port map( D => n3971, CK => clk, RN => rst_BAR, Q
                           => n3970, QN => n_1504);
   clk_r_REG143_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_14_port, CK => clk, 
                           RN => n6056, Q => n_1505, QN => n7777);
   clk_r_REG248_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CK => clk, 
                           RN => rst_BAR, Q => n3968, QN => n_1506);
   clk_r_REG36_S27 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CK => clk, 
                           RN => rst_BAR, Q => n3967, QN => n_1507);
   clk_r_REG252_S27 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CK => clk, 
                           RN => rst_BAR, Q => n3966, QN => n_1508);
   clk_r_REG185_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CK => clk, 
                           RN => n6057, Q => n3965, QN => n_1509);
   clk_r_REG207_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CK => clk, 
                           RN => rst_BAR, Q => n3964, QN => n_1510);
   clk_r_REG208_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CK => clk, 
                           RN => rst_BAR, Q => n3963, QN => n_1511);
   clk_r_REG209_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CK => clk, 
                           RN => rst_BAR, Q => n3962, QN => n_1512);
   clk_r_REG210_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CK => clk, 
                           RN => rst_BAR, Q => n3961, QN => n_1513);
   clk_r_REG211_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CK => clk, 
                           RN => rst_BAR, Q => n3960, QN => n_1514);
   clk_r_REG212_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CK => clk, 
                           RN => rst_BAR, Q => n3959, QN => n_1515);
   clk_r_REG213_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CK => clk, RN => rst_BAR, Q => n3958, QN => n_1516);
   clk_r_REG214_S11 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CK => clk, 
                           RN => rst_BAR, Q => n3957, QN => n_1517);
   clk_r_REG215_S12 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CK => clk, 
                           RN => rst_BAR, Q => n3956, QN => n_1518);
   clk_r_REG144_S12 : DFFR_X1 port map( D => dataout_mul_15_port, CK => clk, RN
                           => rst_BAR, Q => n3955, QN => n_1519);
   clk_r_REG145_S13 : DFFS_X1 port map( D => n3955, CK => clk, SN => rst_BAR, Q
                           => n3954, QN => n_1520);
   clk_r_REG37_S28 : DFFR_X1 port map( D => dataout_mul_16_port, CK => clk, RN 
                           => rst_BAR, Q => n3953, QN => n_1521);
   clk_r_REG253_S28 : DFFR_X1 port map( D => dataout_mul_17_port, CK => clk, RN
                           => rst_BAR, Q => n3952, QN => n_1522);
   clk_r_REG186_S12 : DFFR_X1 port map( D => dataout_mul_18_port, CK => clk, RN
                           => rst_BAR, Q => n3951, QN => n_1523);
   clk_r_REG187_S12 : DFFR_X1 port map( D => dataout_mul_19_port, CK => clk, RN
                           => rst_BAR, Q => n3950, QN => n_1524);
   clk_r_REG189_S12 : DFFR_X1 port map( D => dataout_mul_20_port, CK => clk, RN
                           => rst_BAR, Q => n3949, QN => n_1525);
   clk_r_REG190_S12 : DFFR_X1 port map( D => dataout_mul_21_port, CK => clk, RN
                           => rst_BAR, Q => n3948, QN => n_1526);
   clk_r_REG192_S12 : DFFR_X1 port map( D => dataout_mul_22_port, CK => clk, RN
                           => rst_BAR, Q => n3947, QN => n_1527);
   clk_r_REG193_S12 : DFFR_X1 port map( D => dataout_mul_23_port, CK => clk, RN
                           => rst_BAR, Q => n3946, QN => n_1528);
   clk_r_REG194_S13 : DFFS_X1 port map( D => n3946, CK => clk, SN => rst_BAR, Q
                           => n3945, QN => n_1529);
   clk_r_REG195_S12 : DFFR_X1 port map( D => dataout_mul_24_port, CK => clk, RN
                           => rst_BAR, Q => n3944, QN => n_1530);
   clk_r_REG196_S12 : DFFR_X1 port map( D => dataout_mul_25_port, CK => clk, RN
                           => rst_BAR, Q => n3943, QN => n_1531);
   clk_r_REG198_S12 : DFFR_X1 port map( D => dataout_mul_26_port, CK => clk, RN
                           => rst_BAR, Q => n3942, QN => n_1532);
   clk_r_REG199_S13 : DFFR_X1 port map( D => n3942, CK => clk, RN => rst_BAR, Q
                           => n3941, QN => n_1533);
   clk_r_REG200_S12 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CK => clk, RN => rst_BAR, Q => n3940, QN => n_1534);
   clk_r_REG201_S12 : DFFR_X1 port map( D => dataout_mul_27_port, CK => clk, RN
                           => rst_BAR, Q => n3939, QN => n_1535);
   clk_r_REG202_S13 : DFFR_X1 port map( D => n3939, CK => clk, RN => rst_BAR, Q
                           => n3938, QN => n_1536);
   clk_r_REG203_S13 : DFFR_X1 port map( D => dataout_mul_28_port, CK => clk, RN
                           => rst_BAR, Q => n3937, QN => n_1537);
   clk_r_REG204_S13 : DFFR_X1 port map( D => dataout_mul_29_port, CK => clk, RN
                           => rst_BAR, Q => n3936, QN => n_1538);
   clk_r_REG205_S13 : DFFR_X1 port map( D => dataout_mul_30_port, CK => clk, RN
                           => n6057, Q => n3935, QN => n_1539);
   clk_r_REG206_S13 : DFFS_X1 port map( D => dataout_mul_31_port, CK => clk, SN
                           => rst_BAR, Q => n3934, QN => n_1540);
   clk_r_REG529_S4 : DFFR_X1 port map( D => n2802, CK => clk, RN => rst_BAR, Q 
                           => n3933, QN => n_1541);
   clk_r_REG27_S20 : DFFS_X1 port map( D => n1256, CK => clk, SN => rst_BAR, Q 
                           => n3932, QN => n_1542);
   clk_r_REG592_S3 : DFFS_X1 port map( D => n1958, CK => clk, SN => rst_BAR, Q 
                           => n_1543, QN => n3931);
   clk_r_REG646_S43 : DFFS_X1 port map( D => n1110, CK => clk, SN => rst_BAR, Q
                           => n3930, QN => n_1544);
   clk_r_REG645_S36 : DFFS_X1 port map( D => n1095, CK => clk, SN => rst_BAR, Q
                           => n3929, QN => n_1545);
   clk_r_REG643_S38 : DFFS_X1 port map( D => n1094, CK => clk, SN => rst_BAR, Q
                           => n3928, QN => n_1546);
   clk_r_REG544_S3 : DFFS_X1 port map( D => n1965, CK => clk, SN => n6055, Q =>
                           n_1547, QN => n3927);
   clk_r_REG642_S35 : DFFR_X1 port map( D => n1142, CK => clk, RN => rst_BAR, Q
                           => n3926, QN => n_1548);
   clk_r_REG175_S42 : DFFR_X1 port map( D => n1104, CK => clk, RN => rst_BAR, Q
                           => n3925, QN => n_1549);
   clk_r_REG662_S42 : DFFS_X1 port map( D => n1109, CK => clk, SN => rst_BAR, Q
                           => n3924, QN => n_1550);
   clk_r_REG632_S7 : DFFS_X1 port map( D => n1930, CK => clk, SN => rst_BAR, Q 
                           => n_1551, QN => n3923);
   clk_r_REG356_S7 : DFFR_X1 port map( D => n1301, CK => clk, RN => rst_BAR, Q 
                           => n3922, QN => n_1552);
   clk_r_REG558_S3 : DFFS_X1 port map( D => n6000, CK => clk, SN => rst_BAR, Q 
                           => n7799, QN => n3921);
   clk_r_REG506_S10 : DFFR_X1 port map( D => n1236, CK => clk, RN => rst_BAR, Q
                           => n3920, QN => n_1553);
   clk_r_REG502_S10 : DFFR_X1 port map( D => n1235, CK => clk, RN => rst_BAR, Q
                           => n3919, QN => n_1554);
   clk_r_REG741_S6 : DFFS_X1 port map( D => n1254, CK => clk, SN => rst_BAR, Q 
                           => n3918, QN => n_1555);
   clk_r_REG508_S7 : DFFR_X1 port map( D => n1722, CK => clk, RN => rst_BAR, Q 
                           => n3917, QN => n_1556);
   clk_r_REG494_S10 : DFFR_X1 port map( D => n1720, CK => clk, RN => rst_BAR, Q
                           => n3916, QN => n_1557);
   clk_r_REG458_S10 : DFFS_X1 port map( D => n1247, CK => clk, SN => rst_BAR, Q
                           => n3915, QN => n_1558);
   clk_r_REG507_S10 : DFFS_X1 port map( D => n1249, CK => clk, SN => rst_BAR, Q
                           => n3914, QN => n_1559);
   clk_r_REG616_S14 : DFFR_X1 port map( D => n1394, CK => clk, RN => rst_BAR, Q
                           => n3913, QN => n_1560);
   clk_r_REG625_S6 : DFFR_X1 port map( D => n1334, CK => clk, RN => rst_BAR, Q 
                           => n3912, QN => n7787);
   clk_r_REG518_S10 : DFFS_X1 port map( D => n1278, CK => clk, SN => n6056, Q 
                           => n3911, QN => n_1561);
   clk_r_REG833_S7 : DFFS_X1 port map( D => n1277, CK => clk, SN => rst_BAR, Q 
                           => n3910, QN => n_1562);
   clk_r_REG383_S10 : DFFS_X1 port map( D => n1324, CK => clk, SN => rst_BAR, Q
                           => n_1563, QN => n7819);
   clk_r_REG498_S7 : DFFR_X1 port map( D => n1321, CK => clk, RN => rst_BAR, Q 
                           => n3908, QN => n_1564);
   clk_r_REG424_S24 : DFFR_X1 port map( D => n1366, CK => clk, RN => rst_BAR, Q
                           => n3907, QN => n7786);
   clk_r_REG928_S3 : DFFR_X1 port map( D => n1967, CK => clk, RN => n6056, Q =>
                           n_1565, QN => n3906);
   clk_r_REG496_S7 : DFFS_X1 port map( D => n1354, CK => clk, SN => rst_BAR, Q 
                           => n3905, QN => n_1566);
   clk_r_REG1218_S7 : DFFR_X1 port map( D => n1328, CK => clk, RN => rst_BAR, Q
                           => n3904, QN => n_1567);
   clk_r_REG495_S7 : DFFR_X1 port map( D => n1349, CK => clk, RN => rst_BAR, Q 
                           => n3903, QN => n_1568);
   clk_r_REG492_S7 : DFFS_X1 port map( D => n1393, CK => clk, SN => n6055, Q =>
                           n3902, QN => n_1569);
   clk_r_REG490_S7 : DFFS_X1 port map( D => n2519_port, CK => clk, SN => 
                           rst_BAR, Q => n3901, QN => n_1570);
   clk_r_REG482_S14 : DFFS_X1 port map( D => n1392, CK => clk, SN => rst_BAR, Q
                           => n3900, QN => n_1571);
   clk_r_REG918_S10 : DFFR_X1 port map( D => n1389, CK => clk, RN => rst_BAR, Q
                           => n3899, QN => n_1572);
   clk_r_REG466_S6 : DFFR_X1 port map( D => n1441, CK => clk, RN => n6055, Q =>
                           n3898, QN => n_1573);
   clk_r_REG1300_S4 : DFFS_X1 port map( D => n1430, CK => clk, SN => rst_BAR, Q
                           => n3897, QN => n_1574);
   clk_r_REG517_S10 : DFFS_X1 port map( D => n1428, CK => clk, SN => rst_BAR, Q
                           => n3896, QN => n_1575);
   clk_r_REG1299_S4 : DFFR_X1 port map( D => n1425, CK => clk, RN => rst_BAR, Q
                           => n3895, QN => n_1576);
   clk_r_REG536_S3 : DFFS_X1 port map( D => n1470, CK => clk, SN => rst_BAR, Q 
                           => n3894, QN => n_1577);
   clk_r_REG513_S3 : DFFS_X1 port map( D => n1469, CK => clk, SN => rst_BAR, Q 
                           => n3893, QN => n_1578);
   clk_r_REG1301_S4 : DFFS_X1 port map( D => n1467, CK => clk, SN => rst_BAR, Q
                           => n3892, QN => n_1579);
   clk_r_REG423_S7 : DFFR_X1 port map( D => n1615, CK => clk, RN => rst_BAR, Q 
                           => n3891, QN => n_1580);
   clk_r_REG614_S42 : DFFR_X1 port map( D => n1550, CK => clk, RN => rst_BAR, Q
                           => n3890, QN => n_1581);
   clk_r_REG640_S43 : DFFR_X1 port map( D => n1560, CK => clk, RN => rst_BAR, Q
                           => n3889, QN => n7782);
   clk_r_REG313_S32 : DFFS_X1 port map( D => n1531, CK => clk, SN => rst_BAR, Q
                           => n3888, QN => n_1582);
   clk_r_REG174_S42 : DFFR_X1 port map( D => n1535, CK => clk, RN => n6055, Q 
                           => n3887, QN => n_1583);
   clk_r_REG310_S32 : DFFR_X1 port map( D => n1534, CK => clk, RN => rst_BAR, Q
                           => n3886, QN => n_1584);
   clk_r_REG309_S32 : DFFS_X1 port map( D => n1537, CK => clk, SN => n6056, Q 
                           => n3885, QN => n_1585);
   clk_r_REG308_S32 : DFFS_X1 port map( D => n1542, CK => clk, SN => rst_BAR, Q
                           => n3884, QN => n_1586);
   clk_r_REG639_S45 : DFFS_X1 port map( D => n1584, CK => clk, SN => rst_BAR, Q
                           => n3883, QN => n_1587);
   clk_r_REG635_S46 : DFFR_X1 port map( D => n1908, CK => clk, RN => rst_BAR, Q
                           => n_1588, QN => n3882);
   clk_r_REG631_S7 : DFFR_X1 port map( D => n1633, CK => clk, RN => rst_BAR, Q 
                           => n3881, QN => n_1589);
   clk_r_REG629_S46 : DFFR_X1 port map( D => n1682, CK => clk, RN => rst_BAR, Q
                           => n_1590, QN => n6021);
   clk_r_REG628_S46 : DFFS_X1 port map( D => n1682, CK => clk, SN => rst_BAR, Q
                           => n3879, QN => n_1591);
   clk_r_REG666_S43 : DFFS_X1 port map( D => n1595, CK => clk, SN => rst_BAR, Q
                           => n3878, QN => n_1592);
   clk_r_REG624_S7 : DFFR_X1 port map( D => n1724, CK => clk, RN => n6056, Q =>
                           n3877, QN => n_1593);
   clk_r_REG665_S46 : DFFS_X1 port map( D => n1803, CK => clk, SN => n6055, Q 
                           => n3876, QN => n_1594);
   clk_r_REG621_S12 : DFFS_X1 port map( D => n1979, CK => clk, SN => n6054, Q 
                           => n3875, QN => n_1595);
   clk_r_REG516_S10 : DFFS_X1 port map( D => n1978, CK => clk, SN => rst_BAR, Q
                           => n_1596, QN => n7820);
   clk_r_REG493_S7 : DFFR_X1 port map( D => n2433, CK => clk, RN => n6055, Q =>
                           n3873, QN => n_1597);
   clk_r_REG1481_S10 : DFFR_X1 port map( D => n1974, CK => clk, RN => rst_BAR, 
                           Q => n3872, QN => n_1598);
   clk_r_REG2330_S48 : DFFS_X1 port map( D => n2670, CK => clk, SN => rst_BAR, 
                           Q => n3871, QN => n_1599);
   clk_r_REG102_S48 : DFFS_X1 port map( D => n2011, CK => clk, SN => rst_BAR, Q
                           => n3870, QN => n_1600);
   clk_r_REG2490_S45 : DFFR_X1 port map( D => n1909, CK => clk, RN => rst_BAR, 
                           Q => n_1601, QN => n3869);
   clk_r_REG88_S45 : DFFS_X1 port map( D => n2052, CK => clk, SN => rst_BAR, Q 
                           => n3868, QN => n_1602);
   clk_r_REG197_S13 : DFFS_X1 port map( D => n2078, CK => clk, SN => rst_BAR, Q
                           => n3867, QN => n_1603);
   clk_r_REG81_S43 : DFFS_X1 port map( D => n2075, CK => clk, SN => rst_BAR, Q 
                           => n3866, QN => n_1604);
   clk_r_REG76_S42 : DFFS_X1 port map( D => n2085, CK => clk, SN => rst_BAR, Q 
                           => n3865, QN => n_1605);
   clk_r_REG304_S39 : DFFS_X1 port map( D => n2134, CK => clk, SN => rst_BAR, Q
                           => n3864, QN => n_1606);
   clk_r_REG71_S39 : DFFS_X1 port map( D => n2116, CK => clk, SN => rst_BAR, Q 
                           => n3863, QN => n_1607);
   clk_r_REG1876_S3 : DFFR_X1 port map( D => n2131, CK => clk, RN => rst_BAR, Q
                           => n3862, QN => n_1608);
   clk_r_REG161_S41 : DFFS_X1 port map( D => n2127, CK => clk, SN => rst_BAR, Q
                           => n3861, QN => n_1609);
   clk_r_REG303_S35 : DFFS_X1 port map( D => n2150, CK => clk, SN => rst_BAR, Q
                           => n3860, QN => n_1610);
   clk_r_REG191_S13 : DFFS_X1 port map( D => n2143, CK => clk, SN => n6057, Q 
                           => n3859, QN => n_1611);
   clk_r_REG154_S35 : DFFS_X1 port map( D => n2165, CK => clk, SN => rst_BAR, Q
                           => n3858, QN => n_1612);
   clk_r_REG155_S35 : DFFS_X1 port map( D => n2163, CK => clk, SN => rst_BAR, Q
                           => n3857, QN => n_1613);
   clk_r_REG64_S38 : DFFS_X1 port map( D => n2157, CK => clk, SN => rst_BAR, Q 
                           => n3856, QN => n_1614);
   clk_r_REG3033_S14 : DFFS_X1 port map( D => n2513, CK => clk, SN => rst_BAR, 
                           Q => n3855, QN => n_1615);
   clk_r_REG515_S10 : DFFS_X1 port map( D => n2212, CK => clk, SN => rst_BAR, Q
                           => n3854, QN => n_1616);
   clk_r_REG489_S7 : DFFR_X1 port map( D => n2435, CK => clk, RN => rst_BAR, Q 
                           => n3853, QN => n_1617);
   clk_r_REG152_S35 : DFFS_X1 port map( D => n2226, CK => clk, SN => rst_BAR, Q
                           => n3852, QN => n_1618);
   clk_r_REG188_S36 : DFFS_X1 port map( D => n2220, CK => clk, SN => rst_BAR, Q
                           => n3851, QN => n_1619);
   clk_r_REG151_S35 : DFFR_X1 port map( D => n2244, CK => clk, RN => n6057, Q 
                           => n3850, QN => n_1620);
   clk_r_REG53_S35 : DFFS_X1 port map( D => n2240, CK => clk, SN => rst_BAR, Q 
                           => n3849, QN => n_1621);
   clk_r_REG302_S8 : DFFS_X1 port map( D => n2250, CK => clk, SN => rst_BAR, Q 
                           => n3848, QN => n_1622);
   clk_r_REG254_S29 : DFFS_X1 port map( D => n2267, CK => clk, SN => rst_BAR, Q
                           => n3847, QN => n_1623);
   clk_r_REG46_S32 : DFFR_X1 port map( D => n2262, CK => clk, RN => rst_BAR, Q 
                           => n3846, QN => n_1624);
   clk_r_REG306_S8 : DFFR_X1 port map( D => n2261, CK => clk, RN => rst_BAR, Q 
                           => n3845, QN => n_1625);
   clk_r_REG150_S35 : DFFS_X1 port map( D => n2264, CK => clk, SN => rst_BAR, Q
                           => n3844, QN => n_1626);
   clk_r_REG38_S29 : DFFS_X1 port map( D => n2271, CK => clk, SN => rst_BAR, Q 
                           => n3843, QN => n_1627);
   clk_r_REG299_S8 : DFFR_X1 port map( D => n2294, CK => clk, RN => rst_BAR, Q 
                           => n3842, QN => n_1628);
   clk_r_REG347_S7 : DFFR_X1 port map( D => n2322, CK => clk, RN => n6056, Q =>
                           n3841, QN => n_1629);
   clk_r_REG291_S7 : DFFS_X1 port map( D => n2635, CK => clk, SN => rst_BAR, Q 
                           => n3840, QN => n_1630);
   clk_r_REG512_S10 : DFFS_X1 port map( D => n2319, CK => clk, SN => rst_BAR, Q
                           => n3839, QN => n_1631);
   clk_r_REG345_S7 : DFFS_X1 port map( D => n2340, CK => clk, SN => rst_BAR, Q 
                           => n3838, QN => n_1632);
   clk_r_REG236_S14 : DFFS_X1 port map( D => n2333, CK => clk, SN => rst_BAR, Q
                           => n3837, QN => n_1633);
   clk_r_REG421_S24 : DFFR_X1 port map( D => n2355, CK => clk, RN => rst_BAR, Q
                           => n3836, QN => n_1634);
   clk_r_REG418_S24 : DFFS_X1 port map( D => n2361, CK => clk, SN => n6057, Q 
                           => n3835, QN => n_1635);
   clk_r_REG501_S10 : DFFR_X1 port map( D => n2403, CK => clk, RN => rst_BAR, Q
                           => n3834, QN => n_1636);
   clk_r_REG1083_S23 : DFFS_X1 port map( D => n2399, CK => clk, SN => rst_BAR, 
                           Q => n3833, QN => n_1637);
   clk_r_REG15_S3 : DFFR_X1 port map( D => n1940, CK => clk, RN => rst_BAR, Q 
                           => n_1638, QN => n3832);
   clk_r_REG9_S10 : DFFS_X1 port map( D => n2693, CK => clk, SN => rst_BAR, Q 
                           => n3831, QN => n_1639);
   clk_r_REG52_S35 : DFFS_X1 port map( D => n2529_port, CK => clk, SN => 
                           rst_BAR, Q => n3830, QN => n_1640);
   clk_r_REG354_S7 : DFFS_X1 port map( D => n2527_port, CK => clk, SN => 
                           rst_BAR, Q => n3829, QN => n_1641);
   clk_r_REG45_S32 : DFFS_X1 port map( D => n2542_port, CK => clk, SN => 
                           rst_BAR, Q => n3828, QN => n_1642);
   clk_r_REG834_S7 : DFFS_X1 port map( D => n2541_port, CK => clk, SN => 
                           rst_BAR, Q => n3827, QN => n_1643);
   clk_r_REG63_S38 : DFFS_X1 port map( D => n2539_port, CK => clk, SN => 
                           rst_BAR, Q => n3826, QN => n_1644);
   clk_r_REG13_S12 : DFFR_X1 port map( D => n2596, CK => clk, RN => rst_BAR, Q 
                           => n3825, QN => n_1645);
   clk_r_REG44_S32 : DFFR_X1 port map( D => n2672, CK => clk, RN => rst_BAR, Q 
                           => n3824, QN => n_1646);
   clk_r_REG457_S10 : DFFR_X1 port map( D => n1286, CK => clk, RN => rst_BAR, Q
                           => n3823, QN => n_1647);
   clk_r_REG3034_S14 : DFFS_X1 port map( D => n2209, CK => clk, SN => rst_BAR, 
                           Q => n3822, QN => n_1648);
   clk_r_REG300_S8 : DFFS_X1 port map( D => n2300, CK => clk, SN => rst_BAR, Q 
                           => n3821, QN => n_1649);
   clk_r_REG419_S24 : DFFR_X1 port map( D => n2378, CK => clk, RN => rst_BAR, Q
                           => n3820, QN => n_1650);
   clk_r_REG600_S3 : DFFR_X1 port map( D => n1167, CK => clk, RN => n6056, Q =>
                           n3819, QN => n7779);
   clk_r_REG599_S3 : DFFR_X1 port map( D => n1157, CK => clk, RN => n6056, Q =>
                           n_1651, QN => n6019);
   clk_r_REG598_S3 : DFFS_X1 port map( D => n1157, CK => clk, SN => rst_BAR, Q 
                           => n3817, QN => n_1652);
   clk_r_REG317_S8 : DFFS_X1 port map( D => n1302, CK => clk, SN => rst_BAR, Q 
                           => n3816, QN => n7773);
   clk_r_REG455_S10 : DFFR_X1 port map( D => n2445, CK => clk, RN => rst_BAR, Q
                           => n3815, QN => n_1653);
   clk_r_REG314_S32 : DFFR_X1 port map( D => n1924, CK => clk, RN => rst_BAR, Q
                           => n_1654, QN => n3814);
   clk_r_REG312_S32 : DFFS_X1 port map( D => n1920, CK => clk, SN => rst_BAR, Q
                           => n_1655, QN => n3813);
   clk_r_REG311_S32 : DFFR_X1 port map( D => n1920, CK => clk, RN => rst_BAR, Q
                           => n_1656, QN => n3812);
   clk_r_REG307_S32 : DFFR_X1 port map( D => n1923, CK => clk, RN => rst_BAR, Q
                           => n_1657, QN => n3811);
   clk_r_REG172_S42 : DFFR_X1 port map( D => n1916, CK => clk, RN => rst_BAR, Q
                           => n_1658, QN => n3810);
   clk_r_REG595_S3 : DFFR_X1 port map( D => n1919, CK => clk, RN => n6057, Q =>
                           n_1659, QN => n3809);
   clk_r_REG353_S7 : DFFR_X1 port map( D => n1708, CK => clk, RN => rst_BAR, Q 
                           => n_1660, QN => n6011);
   clk_r_REG352_S7 : DFFS_X1 port map( D => n1708, CK => clk, SN => rst_BAR, Q 
                           => n3807, QN => n7781);
   clk_r_REG351_S7 : DFFR_X1 port map( D => n1728, CK => clk, RN => rst_BAR, Q 
                           => n_1661, QN => n6012);
   clk_r_REG350_S7 : DFFS_X1 port map( D => n1728, CK => clk, SN => rst_BAR, Q 
                           => n3805, QN => n7792);
   clk_r_REG349_S7 : DFFR_X1 port map( D => n1655, CK => clk, RN => rst_BAR, Q 
                           => n3804, QN => n_1662);
   clk_r_REG348_S7 : DFFS_X1 port map( D => n1655, CK => clk, SN => n6056, Q =>
                           n_1663, QN => n6013);
   clk_r_REG454_S10 : DFFS_X1 port map( D => n2441, CK => clk, SN => n6056, Q 
                           => n3802, QN => n_1664);
   clk_r_REG453_S10 : DFFR_X1 port map( D => n2425, CK => clk, RN => rst_BAR, Q
                           => n7778, QN => n6010);
   clk_r_REG275_S8 : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_mux_out_2_20_port, CK => clk, 
                           RN => rst_BAR, Q => n3800, QN => n_1665);
   clk_r_REG3021_S15 : DFFR_X1 port map( D => dataout_mul_1_port, CK => clk, RN
                           => rst_BAR, Q => n3799, QN => n_1666);
   clk_r_REG3022_S16 : DFFR_X1 port map( D => n3799, CK => clk, RN => rst_BAR, 
                           Q => n3798, QN => n_1667);
   clk_r_REG3023_S17 : DFFR_X1 port map( D => n3798, CK => clk, RN => rst_BAR, 
                           Q => n3797, QN => n_1668);
   clk_r_REG3024_S18 : DFFR_X1 port map( D => n3797, CK => clk, RN => rst_BAR, 
                           Q => n3796, QN => n_1669);
   clk_r_REG3025_S19 : DFFR_X1 port map( D => n3796, CK => clk, RN => rst_BAR, 
                           Q => n3795, QN => n_1670);
   clk_r_REG3026_S20 : DFFR_X1 port map( D => n3795, CK => clk, RN => rst_BAR, 
                           Q => n3794, QN => n_1671);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n554, Q => 
                           DATA2_I_30_port);
   clk_r_REG581_S3 : DFFR_X1 port map( D => n5992, CK => clk, RN => rst_BAR, Q 
                           => n7764, QN => n4102);
   clk_r_REG575_S3 : DFFR_X1 port map( D => n5985, CK => clk, RN => rst_BAR, Q 
                           => n4518, QN => n7755);
   clk_r_REG576_S3 : DFFR_X1 port map( D => n5994, CK => clk, RN => rst_BAR, Q 
                           => n7739, QN => n4245);
   clk_r_REG673_S3 : DFFR_X1 port map( D => n1960, CK => clk, RN => n6054, Q =>
                           n7738, QN => n4112);
   clk_r_REG603_S3 : DFFR_X1 port map( D => n1068, CK => clk, RN => rst_BAR, Q 
                           => n7737, QN => n4521);
   clk_r_REG546_S3 : DFFS_X1 port map( D => n1965, CK => clk, SN => rst_BAR, Q 
                           => n4478, QN => n7735);
   clk_r_REG588_S3 : DFFR_X1 port map( D => n1951, CK => clk, RN => rst_BAR, Q 
                           => n7732, QN => n4289);
   clk_r_REG589_S3 : DFFR_X1 port map( D => n1951, CK => clk, RN => rst_BAR, Q 
                           => n4477, QN => n7721);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n7822, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port);
   clk_r_REG590_S3 : DFFS_X1 port map( D => n1950, CK => clk, SN => rst_BAR, Q 
                           => n4519, QN => n7760);
   U3 : CLKBUF_X1 port map( A => n6056, Z => n6054);
   U4 : CLKBUF_X1 port map( A => rst_BAR, Z => n6055);
   U5 : CLKBUF_X1 port map( A => rst_BAR, Z => n6056);
   U6 : CLKBUF_X1 port map( A => rst_BAR, Z => n6057);
   U7 : NOR2_X2 port map( A1 => n6009, A2 => n7488, ZN => n7521);
   U8 : NOR2_X2 port map( A1 => n6008, A2 => n7528, ZN => n7561);
   U9 : NOR2_X2 port map( A1 => n6006, A2 => n7568, ZN => n7601);
   U10 : NOR2_X2 port map( A1 => n6007, A2 => n7607, ZN => n7641);
   U11 : NOR2_X2 port map( A1 => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , A2 => n7379, ZN => n7410);
   U12 : NOR2_X2 port map( A1 => n7486, A2 => n6009, ZN => n7522);
   U13 : NOR2_X2 port map( A1 => n7526, A2 => n6008, ZN => n7562);
   U14 : NOR2_X2 port map( A1 => n7566, A2 => n6006, ZN => n7602);
   U15 : NOR2_X2 port map( A1 => n6005, A2 => n7449, ZN => n7480);
   U16 : NOR3_X4 port map( A1 => n6007, A2 => n4319, A3 => n4314, ZN => n7642);
   U17 : NOR2_X1 port map( A1 => n7829, A2 => n4523, ZN => n7166);
   U18 : INV_X1 port map( A => n554, ZN => n7350);
   U19 : NOR3_X1 port map( A1 => DATA2(0), A2 => n7374, A3 => n7709, ZN => 
                           n7691);
   U20 : NOR2_X1 port map( A1 => n7709, A2 => n7669, ZN => n6101);
   U21 : AND2_X1 port map( A1 => n6444, A2 => n1970, ZN => n7688);
   U22 : CLKBUF_X1 port map( A => n7375, Z => n7370);
   U23 : INV_X1 port map( A => data1_mul_0_port, ZN => n1894);
   U24 : INV_X1 port map( A => data1_mul_15_port, ZN => n1865);
   U25 : NOR2_X1 port map( A1 => FUNC(1), A2 => n7672, ZN => n1901);
   U26 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_5_port, 
                           ZN => n1895);
   U27 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           ZN => n7418);
   U28 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n7418, ZN => n2773);
   U29 : OR2_X1 port map( A1 => n1895, A2 => n2773, ZN => n5989);
   U30 : INV_X1 port map( A => DATA2(31), ZN => n1941);
   U31 : INV_X1 port map( A => DATA2(30), ZN => n1942);
   U32 : INV_X1 port map( A => DATA2(29), ZN => n1943);
   U33 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n1866);
   U34 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n1870);
   U35 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n1868);
   U36 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n1864);
   U37 : NOR2_X1 port map( A1 => DATA2(2), A2 => DATA2(1), ZN => n7662);
   U38 : NAND2_X1 port map( A1 => DATA2(4), A2 => DATA2(3), ZN => n7653);
   U39 : NOR2_X1 port map( A1 => n7662, A2 => n7653, ZN => n7654);
   U40 : INV_X1 port map( A => n7654, ZN => n1967);
   U41 : NAND2_X1 port map( A1 => DATA2(2), A2 => DATA2(0), ZN => n6102);
   U42 : NOR2_X1 port map( A1 => DATA2(1), A2 => n6102, ZN => n6103);
   U43 : INV_X1 port map( A => DATA2(3), ZN => n7661);
   U44 : AND3_X1 port map( A1 => DATA2(4), A2 => n6103, A3 => n7661, ZN => 
                           n6002);
   U45 : NOR2_X1 port map( A1 => DATA2(5), A2 => DATA2(4), ZN => n1959);
   U46 : INV_X1 port map( A => DATA2(1), ZN => n7374);
   U47 : INV_X1 port map( A => DATA2(0), ZN => n7658);
   U48 : NAND2_X1 port map( A1 => n7374, A2 => n7658, ZN => n7666);
   U49 : NOR2_X1 port map( A1 => DATA2(2), A2 => n7666, ZN => n6058);
   U50 : AOI21_X1 port map( B1 => n6058, B2 => n7661, A => n1959, ZN => n1960);
   U51 : INV_X1 port map( A => DATA2(2), ZN => n1970);
   U52 : NAND2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n7669);
   U53 : NOR2_X1 port map( A1 => n7661, A2 => n7669, ZN => n7667);
   U54 : INV_X1 port map( A => n7667, ZN => n7674);
   U55 : OAI21_X1 port map( B1 => n1970, B2 => n7674, A => n1959, ZN => n1964);
   U56 : INV_X1 port map( A => n1964, ZN => n1219);
   U57 : NOR2_X1 port map( A1 => n1959, A2 => n7661, ZN => n1961);
   U58 : NAND2_X1 port map( A1 => DATA2(4), A2 => DATA2(2), ZN => n7677);
   U59 : OR4_X1 port map( A1 => n7374, A2 => n7677, A3 => n1961, A4 => DATA2(0)
                           , ZN => n6000);
   U60 : INV_X1 port map( A => n1961, ZN => n7676);
   U61 : NAND2_X1 port map( A1 => n7676, A2 => n7677, ZN => n7659);
   U62 : INV_X1 port map( A => n7659, ZN => n1963);
   U63 : INV_X1 port map( A => n1959, ZN => n7656);
   U64 : AOI21_X1 port map( B1 => DATA2(2), B2 => DATA2(3), A => n7656, ZN => 
                           n7664);
   U65 : INV_X1 port map( A => n7664, ZN => n7660);
   U66 : OAI21_X1 port map( B1 => DATA2(1), B2 => n7656, A => n7660, ZN => 
                           n1947);
   U67 : NOR2_X1 port map( A1 => n7661, A2 => n6102, ZN => n7665);
   U68 : NAND2_X1 port map( A1 => n7665, A2 => n1947, ZN => n1948);
   U69 : INV_X1 port map( A => n1948, ZN => n2332);
   U70 : INV_X1 port map( A => n1947, ZN => n1102);
   U71 : NOR2_X1 port map( A1 => DATA2(3), A2 => n7656, ZN => n6444);
   U72 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n6069);
   U73 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n6069, 
                           ZN => n1429);
   U74 : INV_X1 port map( A => FUNC(1), ZN => n1903);
   U75 : INV_X1 port map( A => FUNC(0), ZN => n1898);
   U76 : INV_X1 port map( A => FUNC(2), ZN => n1904);
   U77 : NAND3_X1 port map( A1 => n1903, A2 => n1898, A3 => n1904, ZN => n554);
   U78 : INV_X1 port map( A => n7350, ZN => n7829);
   U79 : AND2_X1 port map( A1 => DATA1(3), A2 => DATA2_I_3_port, ZN => n6066);
   U80 : NAND2_X1 port map( A1 => DATA1(2), A2 => DATA2_I_2_port, ZN => n6063);
   U81 : OAI21_X1 port map( B1 => DATA1(2), B2 => DATA2_I_2_port, A => n6063, 
                           ZN => n6810);
   U82 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n6973);
   U83 : INV_X1 port map( A => n6973, ZN => n7160);
   U84 : NAND2_X1 port map( A1 => DATA1(1), A2 => DATA2_I_1_port, ZN => n6065);
   U85 : OAI21_X1 port map( B1 => DATA1(1), B2 => DATA2_I_1_port, A => n6065, 
                           ZN => n6972);
   U86 : INV_X1 port map( A => n6972, ZN => n6974);
   U87 : INV_X1 port map( A => n6065, ZN => n6060);
   U88 : AOI21_X1 port map( B1 => n7160, B2 => n6974, A => n6060, ZN => n6809);
   U89 : OAI21_X1 port map( B1 => n6810, B2 => n6809, A => n6063, ZN => n6059);
   U90 : INV_X1 port map( A => n6059, ZN => n7714);
   U91 : XOR2_X1 port map( A => DATA1(3), B => DATA2_I_3_port, Z => n6068);
   U92 : INV_X1 port map( A => n6068, ZN => n7713);
   U93 : NOR2_X1 port map( A1 => n7714, A2 => n7713, ZN => n7712);
   U94 : NOR2_X1 port map( A1 => n6066, A2 => n7712, ZN => n6374);
   U95 : OAI21_X1 port map( B1 => n6374, B2 => n1429, A => n6069, ZN => n6347);
   U96 : NOR2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n7159);
   U97 : NOR2_X1 port map( A1 => n7159, A2 => n6972, ZN => n6962);
   U98 : NOR2_X1 port map( A1 => n6060, A2 => n6962, ZN => n6807);
   U99 : OAI21_X1 port map( B1 => n6810, B2 => n6807, A => n6063, ZN => n6061);
   U100 : INV_X1 port map( A => n6061, ZN => n6415);
   U101 : NOR2_X1 port map( A1 => n6415, A2 => n7713, ZN => n6414);
   U102 : NOR2_X1 port map( A1 => n6066, A2 => n6414, ZN => n6373);
   U103 : OAI21_X1 port map( B1 => n6373, B2 => n1429, A => n6069, ZN => n6346)
                           ;
   U104 : NAND2_X1 port map( A1 => n7350, A2 => n4523, ZN => n7162);
   U105 : INV_X1 port map( A => n7162, ZN => n6808);
   U106 : AOI22_X1 port map( A1 => n6347, A2 => n7166, B1 => n6346, B2 => n6808
                           , ZN => n6062);
   U107 : INV_X1 port map( A => n6062, ZN => n1861);
   U108 : XOR2_X1 port map( A => DATA1(7), B => DATA2_I_7_port, Z => n1322);
   U109 : XOR2_X1 port map( A => DATA1(5), B => DATA2_I_5_port, Z => n5990);
   U110 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n6286)
                           ;
   U111 : OAI21_X1 port map( B1 => DATA1(6), B2 => DATA2_I_6_port, A => n6286, 
                           ZN => n1353);
   U112 : OAI21_X1 port map( B1 => n4523, B2 => n7160, A => n6962, ZN => n6064)
                           ;
   U113 : OAI221_X1 port map( B1 => n6810, B2 => n6065, C1 => n6810, C2 => 
                           n6064, A => n6063, ZN => n6067);
   U114 : AOI21_X1 port map( B1 => n6068, B2 => n6067, A => n6066, ZN => n6070)
                           ;
   U115 : OAI21_X1 port map( B1 => n6070, B2 => n1429, A => n6069, ZN => n6071)
                           ;
   U116 : AND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n6285);
   U117 : AOI21_X1 port map( B1 => n5990, B2 => n6071, A => n6285, ZN => n6072)
                           ;
   U118 : OAI21_X1 port map( B1 => n6072, B2 => n1353, A => n6286, ZN => n6073)
                           ;
   U119 : AOI22_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, B1 => n1322,
                           B2 => n6073, ZN => n7091);
   U120 : NOR2_X1 port map( A1 => n7829, A2 => n7091, ZN => n7147);
   U121 : INV_X1 port map( A => n7147, ZN => n1859);
   U122 : NAND2_X1 port map( A1 => n7350, A2 => n7091, ZN => n7129);
   U123 : INV_X1 port map( A => n7129, ZN => n1860);
   U124 : INV_X1 port map( A => DATA1(16), ZN => n1929);
   U125 : INV_X1 port map( A => DATA2(14), ZN => n7363);
   U126 : NOR2_X1 port map( A1 => DATA1(14), A2 => n7363, ZN => n7201);
   U127 : INV_X1 port map( A => DATA2(12), ZN => n7365);
   U128 : INV_X1 port map( A => DATA1(12), ZN => n7687);
   U129 : AOI22_X1 port map( A1 => DATA1(12), A2 => n7365, B1 => DATA2(12), B2 
                           => n7687, ZN => n7247);
   U130 : INV_X1 port map( A => n7247, ZN => n6074);
   U131 : INV_X1 port map( A => DATA2(10), ZN => n7367);
   U132 : INV_X1 port map( A => DATA1(11), ZN => n7125);
   U133 : NAND2_X1 port map( A1 => DATA2(11), A2 => n7125, ZN => n7246);
   U134 : OAI21_X1 port map( B1 => DATA1(10), B2 => n7367, A => n7246, ZN => 
                           n7197);
   U135 : INV_X1 port map( A => DATA2(16), ZN => n7361);
   U136 : OAI22_X1 port map( A1 => n1929, A2 => DATA2(16), B1 => n7361, B2 => 
                           DATA1(16), ZN => n7041);
   U137 : INV_X1 port map( A => DATA1(15), ZN => n7695);
   U138 : NAND2_X1 port map( A1 => DATA2(15), A2 => n7695, ZN => n7204);
   U139 : INV_X1 port map( A => n7204, ZN => n7059);
   U140 : OR2_X1 port map( A1 => n7041, A2 => n7059, ZN => n7257);
   U141 : OR4_X1 port map( A1 => n7201, A2 => n6074, A3 => n7197, A4 => n7257, 
                           ZN => n2542_port);
   U142 : NOR2_X1 port map( A1 => FUNC(0), A2 => n1904, ZN => n6497);
   U143 : NAND2_X1 port map( A1 => FUNC(3), A2 => n6497, ZN => n7672);
   U144 : NOR3_X1 port map( A1 => FUNC(0), A2 => FUNC(2), A3 => n1903, ZN => 
                           n6100);
   U145 : INV_X1 port map( A => n6100, ZN => n7161);
   U146 : NOR2_X1 port map( A1 => FUNC(3), A2 => n7161, ZN => n1900);
   U147 : INV_X1 port map( A => n1901, ZN => n7158);
   U148 : INV_X1 port map( A => n1900, ZN => n7143);
   U149 : NAND2_X1 port map( A1 => n7158, A2 => n7143, ZN => n7105);
   U150 : AND3_X1 port map( A1 => n7105, A2 => DATA2(22), A3 => DATA1(22), ZN 
                           => n2131);
   U151 : NAND2_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, ZN => 
                           n7057);
   U152 : OAI21_X1 port map( B1 => DATA1(14), B2 => DATA2_I_14_port, A => n7057
                           , ZN => n2323);
   U153 : NOR2_X1 port map( A1 => DATA2_I_8_port, A2 => DATA1(8), ZN => n6152);
   U154 : AOI21_X1 port map( B1 => DATA1(8), B2 => DATA2_I_8_port, A => n6152, 
                           ZN => n1858);
   U155 : XOR2_X1 port map( A => DATA1(9), B => DATA2_I_9_port, Z => n6151);
   U156 : NAND3_X1 port map( A1 => DATA2_I_8_port, A2 => DATA1(8), A3 => n6151,
                           ZN => n1857);
   U157 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n7052);
   U158 : OAI21_X1 port map( B1 => DATA1(10), B2 => DATA2_I_10_port, A => n7052
                           , ZN => n7145);
   U159 : NAND2_X1 port map( A1 => DATA2_I_13_port, A2 => DATA1(13), ZN => 
                           n7074);
   U160 : OAI21_X1 port map( B1 => DATA2_I_13_port, B2 => DATA1(13), A => n7074
                           , ZN => n7095);
   U161 : NAND2_X1 port map( A1 => DATA1(12), A2 => DATA2_I_12_port, ZN => 
                           n7094);
   U162 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => n7094
                           , ZN => n7111);
   U163 : NOR2_X1 port map( A1 => n7095, A2 => n7111, ZN => n7056);
   U164 : NOR2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => n6076
                           );
   U165 : AOI21_X1 port map( B1 => DATA2_I_11_port, B2 => DATA1(11), A => n6076
                           , ZN => n7133);
   U166 : NAND4_X1 port map( A1 => n1858, A2 => n6151, A3 => n7056, A4 => n7133
                           , ZN => n6075);
   U167 : NOR4_X1 port map( A1 => n7091, A2 => n2323, A3 => n7145, A4 => n6075,
                           ZN => n6079);
   U168 : XOR2_X1 port map( A => DATA1(15), B => DATA2_I_15_port, Z => n7063);
   U169 : INV_X1 port map( A => n6076, ZN => n6077);
   U170 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n7142)
                           ;
   U171 : INV_X1 port map( A => n7142, ZN => n7051);
   U172 : INV_X1 port map( A => n1857, ZN => n6153);
   U173 : INV_X1 port map( A => n7145, ZN => n7050);
   U174 : OAI21_X1 port map( B1 => n7051, B2 => n6153, A => n7050, ZN => n7139)
                           ;
   U175 : NAND2_X1 port map( A1 => n7052, A2 => n7139, ZN => n7132);
   U176 : AOI22_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, B1 => 
                           n6077, B2 => n7132, ZN => n7110);
   U177 : INV_X1 port map( A => n7110, ZN => n7112);
   U178 : INV_X1 port map( A => n7095, ZN => n7090);
   U179 : AND3_X1 port map( A1 => n7090, A2 => DATA1(12), A3 => DATA2_I_12_port
                           , ZN => n7055);
   U180 : AOI21_X1 port map( B1 => n7112, B2 => n7056, A => n7055, ZN => n7076)
                           ;
   U181 : AND2_X1 port map( A1 => n7074, A2 => n7076, ZN => n7073);
   U182 : OAI21_X1 port map( B1 => n7073, B2 => n2323, A => n7057, ZN => n7064)
                           ;
   U183 : AND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => n6078
                           );
   U184 : AOI221_X1 port map( B1 => n6079, B2 => n7063, C1 => n7064, C2 => 
                           n7063, A => n6078, ZN => n6110);
   U185 : NOR2_X1 port map( A1 => n6110, A2 => n7829, ZN => n1856);
   U186 : NAND2_X1 port map( A1 => n7350, A2 => n6110, ZN => n1855);
   U187 : INV_X1 port map( A => n1856, ZN => n7029);
   U188 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n6082);
   U189 : NAND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n7012);
   U190 : NOR2_X1 port map( A1 => DATA2_I_16_port, A2 => DATA1(16), ZN => n7031
                           );
   U191 : OAI21_X1 port map( B1 => DATA1(17), B2 => DATA2_I_17_port, A => n7012
                           , ZN => n7034);
   U192 : NOR2_X1 port map( A1 => n7031, A2 => n7034, ZN => n7030);
   U193 : INV_X1 port map( A => n7030, ZN => n6080);
   U194 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => n6082
                           , ZN => n7011);
   U195 : AOI21_X1 port map( B1 => n7012, B2 => n6080, A => n7011, ZN => n6081)
                           ;
   U196 : INV_X1 port map( A => n6081, ZN => n7015);
   U197 : AND2_X1 port map( A1 => n6082, A2 => n7015, ZN => n6997);
   U198 : INV_X1 port map( A => n7034, ZN => n6083);
   U199 : NAND3_X1 port map( A1 => DATA2_I_16_port, A2 => DATA1(16), A3 => 
                           n6083, ZN => n7032);
   U200 : AOI21_X1 port map( B1 => n7012, B2 => n7032, A => n7011, ZN => n7013)
                           ;
   U201 : AOI21_X1 port map( B1 => DATA2_I_18_port, B2 => DATA1(18), A => n7013
                           , ZN => n6998);
   U202 : OAI22_X1 port map( A1 => n7029, A2 => n6997, B1 => n1855, B2 => n6998
                           , ZN => n6084);
   U203 : INV_X1 port map( A => n6084, ZN => n1853);
   U204 : INV_X1 port map( A => n7166, ZN => n1896);
   U205 : INV_X1 port map( A => DATA1(9), ZN => n6402);
   U206 : NOR2_X1 port map( A1 => DATA2(9), A2 => n6402, ZN => n7242);
   U207 : NAND2_X1 port map( A1 => DATA2(9), A2 => n6402, ZN => n7194);
   U208 : INV_X1 port map( A => n7194, ZN => n7245);
   U209 : OR2_X1 port map( A1 => n7242, A2 => n7245, ZN => n2520_port);
   U210 : NOR2_X1 port map( A1 => DATA2_I_19_port, A2 => DATA1(19), ZN => n6108
                           );
   U211 : NAND2_X1 port map( A1 => DATA2_I_19_port, A2 => DATA1(19), ZN => 
                           n6085);
   U212 : OAI21_X1 port map( B1 => n6108, B2 => n6998, A => n6085, ZN => n6953)
                           ;
   U213 : OAI21_X1 port map( B1 => n6108, B2 => n6997, A => n6085, ZN => n6954)
                           ;
   U214 : OAI22_X1 port map( A1 => n6953, A2 => n1855, B1 => n7029, B2 => n6954
                           , ZN => n6086);
   U215 : INV_X1 port map( A => n6086, ZN => n2163);
   U216 : INV_X1 port map( A => DATA1(13), ZN => n1933);
   U217 : INV_X1 port map( A => FUNC(3), ZN => n1905);
   U218 : NAND2_X1 port map( A1 => n6497, A2 => n1905, ZN => n6096);
   U219 : OR2_X1 port map( A1 => FUNC(1), A2 => n6096, ZN => n7822);
   U220 : NOR4_X1 port map( A1 => DATA2(9), A2 => DATA2(8), A3 => DATA2(7), A4 
                           => DATA2(6), ZN => n6094);
   U221 : INV_X1 port map( A => n7688, ZN => n7709);
   U222 : OR2_X1 port map( A1 => n7709, A2 => n7666, ZN => n7707);
   U223 : INV_X1 port map( A => DATA2(13), ZN => n7364);
   U224 : INV_X1 port map( A => DATA2(11), ZN => n7366);
   U225 : NAND4_X1 port map( A1 => n7364, A2 => n7365, A3 => n7366, A4 => n7367
                           , ZN => n6087);
   U226 : NOR4_X1 port map( A1 => DATA2(15), A2 => DATA2(14), A3 => n7707, A4 
                           => n6087, ZN => n6093);
   U227 : INV_X1 port map( A => DATA1(8), ZN => n7191);
   U228 : INV_X1 port map( A => DATA1(14), ZN => n7080);
   U229 : NAND4_X1 port map( A1 => n7695, A2 => n7191, A3 => n6402, A4 => n7080
                           , ZN => n6091);
   U230 : INV_X1 port map( A => DATA1(10), ZN => n7167);
   U231 : NAND4_X1 port map( A1 => n7167, A2 => n1933, A3 => n7687, A4 => n7125
                           , ZN => n6090);
   U232 : INV_X1 port map( A => DATA1(7), ZN => n7174);
   U233 : INV_X1 port map( A => DATA1(6), ZN => n7175);
   U234 : INV_X1 port map( A => DATA1(5), ZN => n6806);
   U235 : INV_X1 port map( A => DATA1(4), ZN => n7183);
   U236 : NAND4_X1 port map( A1 => n7174, A2 => n7175, A3 => n6806, A4 => n7183
                           , ZN => n6089);
   U237 : OR4_X1 port map( A1 => DATA1(3), A2 => DATA1(2), A3 => DATA1(1), A4 
                           => DATA1(0), ZN => n6088);
   U238 : NOR4_X1 port map( A1 => n6091, A2 => n6090, A3 => n6089, A4 => n6088,
                           ZN => n6092);
   U239 : AOI211_X1 port map( C1 => n6094, C2 => n6093, A => n6092, B => n7822,
                           ZN => n6095);
   U240 : CLKBUF_X1 port map( A => n6095, Z => n7823);
   U241 : NOR2_X1 port map( A1 => n1970, A2 => n7653, ZN => n7657);
   U242 : NAND2_X1 port map( A1 => DATA2(1), A2 => n7657, ZN => n1968);
   U243 : INV_X1 port map( A => DATA2(5), ZN => n7373);
   U244 : OAI211_X1 port map( C1 => n7658, C2 => n1968, A => FUNC(1), B => 
                           n7373, ZN => n7671);
   U245 : NOR2_X1 port map( A1 => n7671, A2 => n6096, ZN => n1902);
   U246 : OR3_X1 port map( A1 => DATA2(1), A2 => n7658, A3 => n7709, ZN => 
                           n7696);
   U247 : INV_X1 port map( A => n7696, ZN => n7825);
   U248 : NOR2_X1 port map( A1 => n7125, A2 => n7707, ZN => n6098);
   U249 : INV_X1 port map( A => n6101, ZN => n7711);
   U250 : NAND2_X1 port map( A1 => DATA1(7), A2 => n7709, ZN => n6410);
   U251 : NAND2_X1 port map( A1 => DATA1(10), A2 => n7825, ZN => n6149);
   U252 : OAI211_X1 port map( C1 => n7711, C2 => n7191, A => n6410, B => n6149,
                           ZN => n6097);
   U253 : AOI211_X1 port map( C1 => n7691, C2 => DATA1(9), A => n6098, B => 
                           n6097, ZN => n1935);
   U254 : NOR2_X1 port map( A1 => n7687, A2 => n7707, ZN => n6146);
   U255 : NOR2_X1 port map( A1 => n7688, A2 => n7191, ZN => n6406);
   U256 : NOR2_X1 port map( A1 => n7125, A2 => n7696, ZN => n7684);
   U257 : INV_X1 port map( A => n7691, ZN => n7708);
   U258 : OAI22_X1 port map( A1 => n6402, A2 => n7711, B1 => n7167, B2 => n7708
                           , ZN => n6099);
   U259 : NOR4_X1 port map( A1 => n6146, A2 => n6406, A3 => n7684, A4 => n6099,
                           ZN => n1934);
   U260 : INV_X1 port map( A => DATA1(25), ZN => n1911);
   U261 : NOR2_X1 port map( A1 => DATA2(25), A2 => n1911, ZN => n7221);
   U262 : INV_X1 port map( A => DATA2(25), ZN => n7353);
   U263 : NOR2_X1 port map( A1 => DATA1(25), A2 => n7353, ZN => n7275);
   U264 : OR2_X1 port map( A1 => n7221, A2 => n7275, ZN => n2521_port);
   U265 : CLKBUF_X1 port map( A => n6100, Z => n7821);
   U266 : CLKBUF_X1 port map( A => n6101, Z => n7824);
   U267 : NAND2_X1 port map( A1 => n7824, A2 => DATA1(28), ZN => n1129);
   U268 : NAND2_X1 port map( A1 => DATA1(27), A2 => n7709, ZN => n6138);
   U269 : AND2_X1 port map( A1 => n6138, A2 => n1129, ZN => n1803);
   U270 : INV_X1 port map( A => DATA1(23), ZN => n1914);
   U271 : INV_X1 port map( A => DATA2(7), ZN => n1946);
   U272 : INV_X1 port map( A => DATA2(24), ZN => n1945);
   U273 : XOR2_X1 port map( A => DATA1(22), B => DATA2_I_22_port, Z => n1847);
   U274 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_116_port, ZN =>
                           n1892);
   U275 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_115_port, ZN =>
                           n1890);
   U276 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_114_port, ZN =>
                           n1888);
   U277 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_113_port, ZN =>
                           n1886);
   U278 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_112_port, ZN =>
                           n1884);
   U279 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_111_port, ZN =>
                           n1882);
   U280 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_110_port, ZN =>
                           n1880);
   U281 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_109_port, ZN =>
                           n1878);
   U282 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_108_port, ZN =>
                           n1876);
   U283 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_107_port, ZN =>
                           n1874);
   U284 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_0_106_port, ZN =>
                           n1872);
   U285 : INV_X1 port map( A => DATA1(28), ZN => n1906);
   U286 : INV_X1 port map( A => DATA2(28), ZN => n1944);
   U287 : OAI21_X1 port map( B1 => n1970, B2 => n7374, A => n6444, ZN => n1068)
                           ;
   U288 : INV_X1 port map( A => n1068, ZN => n6466);
   U289 : NAND2_X1 port map( A1 => n6466, A2 => n6102, ZN => n1952);
   U290 : INV_X1 port map( A => DATA1(1), ZN => n1939);
   U291 : NAND2_X1 port map( A1 => n6444, A2 => n6103, ZN => n1958);
   U292 : INV_X1 port map( A => DATA2_I_25_port, ZN => n6104);
   U293 : NOR2_X1 port map( A1 => n1911, A2 => n6104, ZN => n1843);
   U294 : AOI21_X1 port map( B1 => n1911, B2 => n6104, A => n1843, ZN => n1844)
                           ;
   U295 : NOR2_X1 port map( A1 => DATA2_I_24_port, A2 => DATA1(24), ZN => n6107
                           );
   U296 : INV_X1 port map( A => n1844, ZN => n6496);
   U297 : NOR2_X1 port map( A1 => n6107, A2 => n6496, ZN => n2070);
   U298 : INV_X1 port map( A => DATA1(26), ZN => n1910);
   U299 : INV_X1 port map( A => DATA2_I_26_port, ZN => n6105);
   U300 : NOR2_X1 port map( A1 => n1910, A2 => n6105, ZN => n6015);
   U301 : AOI21_X1 port map( B1 => n1910, B2 => n6105, A => n6015, ZN => n2058)
                           ;
   U302 : OAI21_X1 port map( B1 => n1843, B2 => n2070, A => n2058, ZN => n6106)
                           ;
   U303 : INV_X1 port map( A => n6106, ZN => n1842);
   U304 : INV_X1 port map( A => n6107, ZN => n1845);
   U305 : AOI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => n6108
                           , ZN => n1852);
   U306 : AOI21_X1 port map( B1 => DATA1(16), B2 => DATA2_I_16_port, A => n7031
                           , ZN => n1854);
   U307 : INV_X1 port map( A => DATA1(20), ZN => n1922);
   U308 : XNOR2_X1 port map( A => DATA2_I_20_port, B => n1922, ZN => n1850);
   U309 : INV_X1 port map( A => DATA1(21), ZN => n1921);
   U310 : XNOR2_X1 port map( A => DATA2_I_21_port, B => n1921, ZN => n1849);
   U311 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n6917);
   U312 : NAND4_X1 port map( A1 => n1852, A2 => n1854, A3 => n1850, A4 => n1849
                           , ZN => n6109);
   U313 : NOR4_X1 port map( A1 => n6110, A2 => n7034, A3 => n7011, A4 => n6109,
                           ZN => n6111);
   U314 : AOI22_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, B1 => 
                           n1850, B2 => n6953, ZN => n7717);
   U315 : INV_X1 port map( A => n7717, ZN => n6946);
   U316 : AND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => n6911
                           );
   U317 : AOI21_X1 port map( B1 => n6946, B2 => n1849, A => n6911, ZN => n6912)
                           ;
   U318 : INV_X1 port map( A => n6912, ZN => n6914);
   U319 : OAI21_X1 port map( B1 => n6111, B2 => n6914, A => n1847, ZN => n6113)
                           ;
   U320 : NAND2_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, ZN => 
                           n6112);
   U321 : OAI21_X1 port map( B1 => DATA1(23), B2 => DATA2_I_23_port, A => n6112
                           , ZN => n6919);
   U322 : AOI21_X1 port map( B1 => n6917, B2 => n6113, A => n6919, ZN => n6114)
                           ;
   U323 : AOI21_X1 port map( B1 => DATA2_I_23_port, B2 => DATA1(23), A => n6114
                           , ZN => n7670);
   U324 : NAND2_X1 port map( A1 => n7350, A2 => n7670, ZN => n1846);
   U325 : AOI21_X1 port map( B1 => n6444, B2 => n7658, A => n6466, ZN => n1950)
                           ;
   U326 : INV_X1 port map( A => n7666, ZN => n7678);
   U327 : NAND4_X1 port map( A1 => DATA2(3), A2 => n1959, A3 => n7678, A4 => 
                           n1970, ZN => n1965);
   U328 : INV_X1 port map( A => DATA1(18), ZN => n1925);
   U329 : NAND2_X1 port map( A1 => n6444, A2 => n1950, ZN => n1951);
   U330 : INV_X1 port map( A => n7707, ZN => n7827);
   U331 : INV_X1 port map( A => n7708, ZN => n7828);
   U332 : AOI22_X1 port map( A1 => DATA1(14), A2 => n7709, B1 => DATA1(18), B2 
                           => n7827, ZN => n6115);
   U333 : NAND2_X1 port map( A1 => DATA1(15), A2 => n7824, ZN => n6144);
   U334 : NAND2_X1 port map( A1 => DATA1(17), A2 => n7825, ZN => n6135);
   U335 : NAND2_X1 port map( A1 => DATA1(16), A2 => n7828, ZN => n6133);
   U336 : NAND4_X1 port map( A1 => n6115, A2 => n6144, A3 => n6135, A4 => n6133
                           , ZN => n1926);
   U337 : INV_X1 port map( A => n7696, ZN => n7826);
   U338 : INV_X1 port map( A => DATA1(27), ZN => n1907);
   U339 : INV_X1 port map( A => DATA1(24), ZN => n1912);
   U340 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_27_port, ZN => 
                           n1867);
   U341 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_28_port, ZN => 
                           n1869);
   U342 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_64_port, ZN => 
                           n1893);
   U343 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_63_port, ZN => 
                           n1891);
   U344 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_62_port, ZN => 
                           n1889);
   U345 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_61_port, ZN => 
                           n1887);
   U346 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_60_port, ZN => 
                           n1885);
   U347 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_59_port, ZN => 
                           n1883);
   U348 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_34_port, ZN => 
                           n1881);
   U349 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_33_port, ZN => 
                           n1879);
   U350 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_32_port, ZN => 
                           n1877);
   U351 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_31_port, ZN => 
                           n1875);
   U352 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_30_port, ZN => 
                           n1873);
   U353 : INV_X1 port map( A => boothmul_pipelined_i_muxes_in_4_29_port, ZN => 
                           n1871);
   U354 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n1895, ZN => n2808);
   U355 : AOI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, A
                           => n2808, ZN => n2802);
   U356 : NOR3_X1 port map( A1 => n4111, A2 => n1894, A3 => n7771, ZN => n3026)
                           ;
   U357 : AOI221_X1 port map( B1 => n4111, B2 => n7771, C1 => n1894, C2 => 
                           n7771, A => n3026, ZN => dataout_mul_4_port);
   U358 : NAND2_X1 port map( A1 => n4294, A2 => n4295, ZN => n6116);
   U359 : OAI21_X1 port map( B1 => n4294, B2 => n4295, A => n6116, ZN => n7449)
                           ;
   U360 : INV_X1 port map( A => boothmul_pipelined_i_sum_B_in_3_6_port, ZN => 
                           n6117);
   U361 : NOR3_X1 port map( A1 => n1894, A2 => n7449, A3 => n6117, ZN => n3030)
                           ;
   U362 : OR2_X1 port map( A1 => n1894, A2 => n7449, ZN => n6118);
   U363 : AOI21_X1 port map( B1 => n6118, B2 => n6117, A => n3030, ZN => 
                           dataout_mul_6_port);
   U364 : NAND2_X1 port map( A1 => n4296, A2 => n4298, ZN => n6119);
   U365 : OAI21_X1 port map( B1 => n4296, B2 => n4298, A => n6119, ZN => n7488)
                           ;
   U366 : NOR3_X1 port map( A1 => n7488, A2 => n7743, A3 => n7774, ZN => n3029)
                           ;
   U367 : INV_X1 port map( A => n7488, ZN => n7487);
   U368 : NAND2_X1 port map( A1 => n7487, A2 => n4332, ZN => n6120);
   U369 : AOI21_X1 port map( B1 => n6120, B2 => n7774, A => n3029, ZN => 
                           dataout_mul_8_port);
   U370 : NAND2_X1 port map( A1 => n4300, A2 => n4303, ZN => n6121);
   U371 : OAI21_X1 port map( B1 => n4300, B2 => n4303, A => n6121, ZN => n7528)
                           ;
   U372 : NOR3_X1 port map( A1 => n7528, A2 => n7744, A3 => n7775, ZN => n3028)
                           ;
   U373 : INV_X1 port map( A => n7528, ZN => n7527);
   U374 : NAND2_X1 port map( A1 => n7527, A2 => n4331, ZN => n6122);
   U375 : AOI21_X1 port map( B1 => n6122, B2 => n7775, A => n3028, ZN => 
                           dataout_mul_10_port);
   U376 : NAND2_X1 port map( A1 => n4306, A2 => n4310, ZN => n6123);
   U377 : OAI21_X1 port map( B1 => n4306, B2 => n4310, A => n6123, ZN => n7568)
                           ;
   U378 : NOR3_X1 port map( A1 => n7568, A2 => n7745, A3 => n7776, ZN => n3027)
                           ;
   U379 : INV_X1 port map( A => n7568, ZN => n7567);
   U380 : NAND2_X1 port map( A1 => n7567, A2 => n4330, ZN => n6124);
   U381 : AOI21_X1 port map( B1 => n6124, B2 => n7776, A => n3027, ZN => 
                           dataout_mul_12_port);
   U382 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n7652);
   U383 : INV_X1 port map( A => n7652, ZN => n7646);
   U384 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN 
                           => n7377);
   U385 : NAND2_X1 port map( A1 => n7377, A2 => data2_mul_1_port, ZN => n7645);
   U386 : INV_X1 port map( A => n7645, ZN => n7650);
   U387 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => n7377, ZN => n7649);
   U388 : AOI222_X1 port map( A1 => n7646, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           n7650, B2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, C1 => 
                           n7649, C2 => boothmul_pipelined_i_muxes_in_4_63_port
                           , ZN => n6126);
   U389 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n7413);
   U390 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n7413, ZN => n7380);
   U391 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n7380, ZN => n6125);
   U392 : NOR2_X1 port map( A1 => n6126, A2 => n6125, ZN => n3036);
   U393 : AOI21_X1 port map( B1 => n6126, B2 => n6125, A => n3036, ZN => 
                           dataout_mul_2_port);
   U394 : AOI22_X1 port map( A1 => n7821, A2 => n2520_port, B1 => n7823, B2 => 
                           n4003, ZN => n1256);
   U395 : NOR2_X1 port map( A1 => n1914, A2 => n7711, ZN => n6474);
   U396 : NAND2_X1 port map( A1 => DATA1(21), A2 => n7825, ZN => n6445);
   U397 : NAND2_X1 port map( A1 => DATA1(22), A2 => n7828, ZN => n6439);
   U398 : OAI211_X1 port map( C1 => n7688, C2 => n1912, A => n6445, B => n6439,
                           ZN => n6127);
   U399 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(20), A => n6474, B => 
                           n6127, ZN => n1084);
   U400 : NOR2_X1 port map( A1 => n7688, A2 => n1911, ZN => n6477);
   U401 : INV_X1 port map( A => n7707, ZN => n7692);
   U402 : NAND2_X1 port map( A1 => DATA1(21), A2 => n7692, ZN => n6448);
   U403 : NAND2_X1 port map( A1 => DATA1(22), A2 => n7825, ZN => n6457);
   U404 : OAI211_X1 port map( C1 => n7708, C2 => n1914, A => n6448, B => n6457,
                           ZN => n6128);
   U405 : AOI211_X1 port map( C1 => n7824, C2 => DATA1(24), A => n6477, B => 
                           n6128, ZN => n1105);
   U406 : NOR2_X1 port map( A1 => n1911, A2 => n7711, ZN => n6475);
   U407 : NAND2_X1 port map( A1 => DATA1(22), A2 => n7692, ZN => n6129);
   U408 : NAND2_X1 port map( A1 => DATA1(23), A2 => n7825, ZN => n6438);
   U409 : OAI211_X1 port map( C1 => n7688, C2 => n1910, A => n6129, B => n6438,
                           ZN => n6130);
   U410 : AOI211_X1 port map( C1 => n7828, C2 => DATA1(24), A => n6475, B => 
                           n6130, ZN => n1110);
   U411 : NOR2_X1 port map( A1 => n1925, A2 => n7711, ZN => n6450);
   U412 : INV_X1 port map( A => DATA1(19), ZN => n7000);
   U413 : NAND2_X1 port map( A1 => DATA1(17), A2 => n7828, ZN => n6131);
   U414 : NAND2_X1 port map( A1 => DATA1(16), A2 => n7825, ZN => n6462);
   U415 : OAI211_X1 port map( C1 => n7688, C2 => n7000, A => n6131, B => n6462,
                           ZN => n6132);
   U416 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(15), A => n6450, B => 
                           n6132, ZN => n1120);
   U417 : INV_X1 port map( A => DATA1(17), ZN => n7027);
   U418 : NOR2_X1 port map( A1 => n7027, A2 => n7711, ZN => n6453);
   U419 : NAND2_X1 port map( A1 => DATA1(14), A2 => n7692, ZN => n6480);
   U420 : OAI211_X1 port map( C1 => n7688, C2 => n1925, A => n6133, B => n6480,
                           ZN => n6134);
   U421 : AOI211_X1 port map( C1 => n7826, C2 => DATA1(15), A => n6453, B => 
                           n6134, ZN => n1142);
   U422 : NOR2_X1 port map( A1 => n7000, A2 => n7711, ZN => n6447);
   U423 : NAND2_X1 port map( A1 => DATA1(18), A2 => n7828, ZN => n6451);
   U424 : OAI211_X1 port map( C1 => n7707, C2 => n1929, A => n6451, B => n6135,
                           ZN => n6136);
   U425 : AOI211_X1 port map( C1 => DATA1(20), C2 => n7709, A => n6447, B => 
                           n6136, ZN => n1095);
   U426 : OAI222_X1 port map( A1 => n1958, A2 => n1120, B1 => n1952, B2 => 
                           n1142, C1 => n1095, C2 => n6466, ZN => n1167);
   U427 : NOR2_X1 port map( A1 => n1922, A2 => n7711, ZN => n6459);
   U428 : NAND2_X1 port map( A1 => DATA1(18), A2 => n7825, ZN => n6454);
   U429 : NAND2_X1 port map( A1 => DATA1(17), A2 => n7692, ZN => n6463);
   U430 : OAI211_X1 port map( C1 => n7708, C2 => n7000, A => n6454, B => n6463,
                           ZN => n6137);
   U431 : AOI211_X1 port map( C1 => DATA1(21), C2 => n7709, A => n6459, B => 
                           n6137, ZN => n1094);
   U432 : OAI222_X1 port map( A1 => n1958, A2 => n1095, B1 => n1952, B2 => 
                           n1120, C1 => n1094, C2 => n6466, ZN => n1157);
   U433 : NAND2_X1 port map( A1 => DATA1(23), A2 => n7692, ZN => n6139);
   U434 : OAI211_X1 port map( C1 => n7696, C2 => n1912, A => n6139, B => n6138,
                           ZN => n1104);
   U435 : AOI22_X1 port map( A1 => DATA1(24), A2 => n7692, B1 => DATA1(28), B2 
                           => n7709, ZN => n1109);
   U436 : NAND2_X1 port map( A1 => n7824, A2 => DATA1(27), ZN => n1677);
   U437 : NAND2_X1 port map( A1 => n7828, A2 => DATA1(27), ZN => n1594);
   U438 : NOR2_X1 port map( A1 => n7688, A2 => n7695, ZN => n6140);
   U439 : NOR2_X1 port map( A1 => n1933, A2 => n7708, ZN => n6483);
   U440 : AOI211_X1 port map( C1 => n7824, C2 => DATA1(14), A => n6140, B => 
                           n6483, ZN => n6141);
   U441 : NAND2_X1 port map( A1 => DATA1(12), A2 => n7825, ZN => n6488);
   U442 : OAI211_X1 port map( C1 => n7707, C2 => n7125, A => n6141, B => n6488,
                           ZN => n1178);
   U443 : NOR2_X1 port map( A1 => n1929, A2 => n7711, ZN => n6456);
   U444 : NAND2_X1 port map( A1 => DATA1(17), A2 => n7709, ZN => n6142);
   U445 : NAND2_X1 port map( A1 => DATA1(15), A2 => n7828, ZN => n6461);
   U446 : OAI211_X1 port map( C1 => n7707, C2 => n1933, A => n6142, B => n6461,
                           ZN => n6143);
   U447 : AOI211_X1 port map( C1 => n7826, C2 => DATA1(14), A => n6456, B => 
                           n6143, ZN => n1927);
   U448 : NAND2_X1 port map( A1 => DATA1(13), A2 => n7825, ZN => n6479);
   U449 : OAI211_X1 port map( C1 => n7688, C2 => n1929, A => n6144, B => n6479,
                           ZN => n6145);
   U450 : AOI211_X1 port map( C1 => n7691, C2 => DATA1(14), A => n6146, B => 
                           n6145, ZN => n1930);
   U451 : INV_X1 port map( A => n1952, ZN => n6969);
   U452 : OAI22_X1 port map( A1 => n6466, A2 => n1927, B1 => n1930, B2 => n1958
                           , ZN => n6147);
   U453 : AOI21_X1 port map( B1 => n6969, B2 => n1178, A => n6147, ZN => n1302)
                           ;
   U454 : NOR2_X1 port map( A1 => n7125, A2 => n7708, ZN => n6486);
   U455 : NOR2_X1 port map( A1 => n7687, A2 => n7711, ZN => n6148);
   U456 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(9), A => n6486, B => 
                           n6148, ZN => n6150);
   U457 : OAI211_X1 port map( C1 => n7688, C2 => n1933, A => n6150, B => n6149,
                           ZN => n1301);
   U458 : NOR2_X1 port map( A1 => n7708, A2 => n1906, ZN => n1680);
   U459 : NAND2_X1 port map( A1 => n7825, A2 => DATA1(28), ZN => n1593);
   U460 : INV_X1 port map( A => n6151, ZN => n6154);
   U461 : NOR2_X1 port map( A1 => n6152, A2 => n6154, ZN => n7146);
   U462 : AOI211_X1 port map( C1 => n6152, C2 => n6154, A => n7146, B => n1859,
                           ZN => n1236);
   U463 : NAND2_X1 port map( A1 => DATA2_I_8_port, A2 => DATA1(8), ZN => n6155)
                           ;
   U464 : AOI211_X1 port map( C1 => n6155, C2 => n6154, A => n6153, B => n7129,
                           ZN => n1235);
   U465 : NAND3_X1 port map( A1 => DATA2(9), A2 => DATA1(9), A3 => n7105, ZN =>
                           n1254);
   U466 : NOR2_X1 port map( A1 => n7175, A2 => n7711, ZN => n6158);
   U467 : NOR2_X1 port map( A1 => n7174, A2 => n7708, ZN => n6157);
   U468 : NOR2_X1 port map( A1 => n7688, A2 => n6806, ZN => n6965);
   U469 : OAI22_X1 port map( A1 => n7191, A2 => n7696, B1 => n6402, B2 => n7707
                           , ZN => n6156);
   U470 : NOR4_X1 port map( A1 => n6158, A2 => n6157, A3 => n6965, A4 => n6156,
                           ZN => n1722);
   U471 : NOR2_X1 port map( A1 => n7175, A2 => n7708, ZN => n6407);
   U472 : NAND2_X1 port map( A1 => DATA1(8), A2 => n7692, ZN => n6264);
   U473 : NAND2_X1 port map( A1 => DATA1(4), A2 => n7709, ZN => n7682);
   U474 : OAI211_X1 port map( C1 => n7711, C2 => n6806, A => n6264, B => n7682,
                           ZN => n6159);
   U475 : AOI211_X1 port map( C1 => n7825, C2 => DATA1(7), A => n6407, B => 
                           n6159, ZN => n1720);
   U476 : NOR2_X1 port map( A1 => n7183, A2 => n7711, ZN => n6162);
   U477 : INV_X1 port map( A => DATA1(3), ZN => n6400);
   U478 : NAND2_X1 port map( A1 => DATA1(5), A2 => n7828, ZN => n6160);
   U479 : NAND2_X1 port map( A1 => DATA1(6), A2 => n7826, ZN => n6404);
   U480 : OAI211_X1 port map( C1 => n7688, C2 => n6400, A => n6160, B => n6404,
                           ZN => n6161);
   U481 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(7), A => n6162, B => 
                           n6161, ZN => n1247);
   U482 : NOR2_X1 port map( A1 => n7183, A2 => n7708, ZN => n6803);
   U483 : INV_X1 port map( A => DATA1(2), ZN => n7227);
   U484 : NAND2_X1 port map( A1 => DATA1(6), A2 => n7692, ZN => n6317);
   U485 : NAND2_X1 port map( A1 => DATA1(3), A2 => n7824, ZN => n7681);
   U486 : OAI211_X1 port map( C1 => n7688, C2 => n7227, A => n6317, B => n7681,
                           ZN => n6163);
   U487 : AOI211_X1 port map( C1 => n7826, C2 => DATA1(5), A => n6803, B => 
                           n6163, ZN => n1249);
   U488 : OAI211_X1 port map( C1 => n4511, C2 => n6022, A => n4232, B => n4231,
                           ZN => n6164);
   U489 : AOI211_X1 port map( C1 => n4499, C2 => n7762, A => n4233, B => n6164,
                           ZN => n6880);
   U490 : NAND4_X1 port map( A1 => n4241, A2 => n3924, A3 => n4239, A4 => n4240
                           , ZN => n6169);
   U491 : INV_X1 port map( A => n6169, ZN => n6166);
   U492 : AOI22_X1 port map( A1 => n4522, A2 => n4536, B1 => n4515, B2 => n7762
                           , ZN => n6165);
   U493 : AND4_X1 port map( A1 => n4236, A2 => n4238, A3 => n4237, A4 => n6165,
                           ZN => n6179);
   U494 : OAI222_X1 port map( A1 => n4521, A2 => n6880, B1 => n4483, B2 => 
                           n6166, C1 => n4496, C2 => n6179, ZN => n6939);
   U495 : INV_X1 port map( A => n6939, ZN => n6926);
   U496 : OAI222_X1 port map( A1 => n4521, A2 => n3930, B1 => n4504, B2 => 
                           n4247, C1 => n4496, C2 => n4104, ZN => n6198);
   U497 : AOI211_X1 port map( C1 => n4492, C2 => n4537, A => n4242, B => n3925,
                           ZN => n6167);
   U498 : OAI222_X1 port map( A1 => n4521, A2 => n6167, B1 => n4483, B2 => 
                           n4104, C1 => n4482, C2 => n3930, ZN => n6187);
   U499 : AOI22_X1 port map( A1 => n6198, A2 => n4489, B1 => n6187, B2 => n4289
                           , ZN => n6171);
   U500 : OAI222_X1 port map( A1 => n6167, A2 => n4503, B1 => n6179, B2 => 
                           n4521, C1 => n6166, C2 => n4482, ZN => n6938);
   U501 : OAI22_X1 port map( A1 => n4482, A2 => n6167, B1 => n3930, B2 => n4503
                           , ZN => n6168);
   U502 : AOI21_X1 port map( B1 => n7737, B2 => n6169, A => n6168, ZN => n6184)
                           ;
   U503 : INV_X1 port map( A => n6184, ZN => n6937);
   U504 : AOI22_X1 port map( A1 => n7764, A2 => n6938, B1 => n6937, B2 => n4480
                           , ZN => n6170);
   U505 : OAI211_X1 port map( C1 => n7772, C2 => n6926, A => n6171, B => n6170,
                           ZN => n7020);
   U506 : INV_X1 port map( A => n7020, ZN => n7001);
   U507 : OAI22_X1 port map( A1 => n4482, A2 => n4246, B1 => n4504, B2 => n4481
                           , ZN => n6172);
   U508 : AOI21_X1 port map( B1 => n7737, B2 => n7783, A => n6172, ZN => n6194)
                           ;
   U509 : INV_X1 port map( A => n6194, ZN => n6182);
   U510 : OAI222_X1 port map( A1 => n4521, A2 => n4247, B1 => n4483, B2 => 
                           n4487, C1 => n4482, C2 => n4481, ZN => n6209);
   U511 : AOI22_X1 port map( A1 => n4289, A2 => n6182, B1 => n4489, B2 => n6209
                           , ZN => n6174);
   U512 : AOI22_X1 port map( A1 => n4474, A2 => n6187, B1 => n4480, B2 => n6198
                           , ZN => n6173);
   U513 : OAI211_X1 port map( C1 => n4290, C2 => n6184, A => n6174, B => n6173,
                           ZN => n7017);
   U514 : OAI22_X1 port map( A1 => n4487, A2 => n4496, B1 => n4504, B2 => n3928
                           , ZN => n6175);
   U515 : AOI21_X1 port map( B1 => n7737, B2 => n7784, A => n6175, ZN => n6206)
                           ;
   U516 : AOI22_X1 port map( A1 => n4474, A2 => n6198, B1 => n4480, B2 => n6182
                           , ZN => n6177);
   U517 : AOI22_X1 port map( A1 => n4505, A2 => n6187, B1 => n4289, B2 => n6209
                           , ZN => n6176);
   U518 : OAI211_X1 port map( C1 => n4519, C2 => n6206, A => n6177, B => n6176,
                           ZN => n6225);
   U519 : AOI22_X1 port map( A1 => n4518, A2 => n7017, B1 => n4475, B2 => n6225
                           , ZN => n6189);
   U520 : AOI22_X1 port map( A1 => n4289, A2 => n6937, B1 => n4489, B2 => n6187
                           , ZN => n6181);
   U521 : NAND2_X1 port map( A1 => n7762, A2 => n4488, ZN => n6674);
   U522 : AOI22_X1 port map( A1 => n7742, A2 => n7780, B1 => n7726, B2 => n4515
                           , ZN => n6178);
   U523 : AND4_X1 port map( A1 => n6674, A2 => n7793, A3 => n4229, A4 => n6178,
                           ZN => n6881);
   U524 : OAI222_X1 port map( A1 => n4521, A2 => n6881, B1 => n4483, B2 => 
                           n6179, C1 => n4496, C2 => n6880, ZN => n6940);
   U525 : AOI22_X1 port map( A1 => n4480, A2 => n6938, B1 => n4459, B2 => n6940
                           , ZN => n6180);
   U526 : OAI211_X1 port map( C1 => n4102, C2 => n6926, A => n6181, B => n6180,
                           ZN => n7019);
   U527 : AOI22_X1 port map( A1 => n7760, A2 => n6182, B1 => n6198, B2 => n4289
                           , ZN => n6183);
   U528 : INV_X1 port map( A => n6183, ZN => n6186);
   U529 : INV_X1 port map( A => n6938, ZN => n6925);
   U530 : OAI22_X1 port map( A1 => n4290, A2 => n6925, B1 => n4102, B2 => n6184
                           , ZN => n6185);
   U531 : AOI211_X1 port map( C1 => n7735, C2 => n6187, A => n6186, B => n6185,
                           ZN => n7002);
   U532 : INV_X1 port map( A => n7002, ZN => n7018);
   U533 : AOI22_X1 port map( A1 => n4473, A2 => n7019, B1 => n4468, B2 => n7018
                           , ZN => n6188);
   U534 : OAI211_X1 port map( C1 => n4472, C2 => n7001, A => n6189, B => n6188,
                           ZN => n7043);
   U535 : OAI22_X1 port map( A1 => n3929, A2 => n4504, B1 => n3928, B2 => n4496
                           , ZN => n6190);
   U536 : AOI21_X1 port map( B1 => n7737, B2 => n7785, A => n6190, ZN => n6216)
                           ;
   U537 : INV_X1 port map( A => n6216, ZN => n6203);
   U538 : INV_X1 port map( A => n6209, ZN => n6195);
   U539 : OAI22_X1 port map( A1 => n4519, A2 => n6019, B1 => n6195, B2 => n7767
                           , ZN => n6192);
   U540 : OAI22_X1 port map( A1 => n4478, A2 => n6206, B1 => n4290, B2 => n6194
                           , ZN => n6191);
   U541 : AOI211_X1 port map( C1 => n7721, C2 => n6203, A => n6192, B => n6191,
                           ZN => n6228);
   U542 : INV_X1 port map( A => n6225, ZN => n6193);
   U543 : OAI22_X1 port map( A1 => n4245, A2 => n6228, B1 => n6193, B2 => n7719
                           , ZN => n6200);
   U544 : OAI22_X1 port map( A1 => n4519, A2 => n6216, B1 => n4102, B2 => n6194
                           , ZN => n6197);
   U545 : OAI22_X1 port map( A1 => n4478, A2 => n6195, B1 => n4477, B2 => n6206
                           , ZN => n6196);
   U546 : AOI211_X1 port map( C1 => n4505, C2 => n6198, A => n6197, B => n6196,
                           ZN => n6220);
   U547 : OAI22_X1 port map( A1 => n4476, A2 => n7002, B1 => n4244, B2 => n6220
                           , ZN => n6199);
   U548 : AOI211_X1 port map( C1 => n7727, C2 => n7017, A => n6200, B => n6199,
                           ZN => n6233);
   U549 : INV_X1 port map( A => n6233, ZN => n6229);
   U550 : INV_X1 port map( A => n6220, ZN => n6224);
   U551 : AOI22_X1 port map( A1 => n4518, A2 => n6225, B1 => n7739, B2 => n6224
                           , ZN => n6202);
   U552 : AOI22_X1 port map( A1 => n4243, A2 => n7018, B1 => n7756, B2 => n7017
                           , ZN => n6201);
   U553 : OAI211_X1 port map( C1 => n4476, C2 => n7001, A => n6202, B => n6201,
                           ZN => n7042);
   U554 : AOI222_X1 port map( A1 => n7043, A2 => n4256, B1 => n6229, B2 => 
                           n4455, C1 => n7042, C2 => n4456, ZN => n7082);
   U555 : AOI22_X1 port map( A1 => n3927, A2 => n3817, B1 => n3819, B2 => n7721
                           , ZN => n6205);
   U556 : OAI222_X1 port map( A1 => n4521, A2 => n4100, B1 => n3926, B2 => 
                           n4482, C1 => n4483, C2 => n4470, ZN => n6239);
   U557 : AOI22_X1 port map( A1 => n4103, A2 => n6239, B1 => n4469, B2 => n6203
                           , ZN => n6204);
   U558 : OAI211_X1 port map( C1 => n6206, C2 => n7770, A => n6205, B => n6204,
                           ZN => n6244);
   U559 : INV_X1 port map( A => n6244, ZN => n6219);
   U560 : OAI22_X1 port map( A1 => n4519, A2 => n7779, B1 => n4477, B2 => n6019
                           , ZN => n6208);
   U561 : OAI22_X1 port map( A1 => n4478, A2 => n6216, B1 => n4102, B2 => n6206
                           , ZN => n6207);
   U562 : AOI211_X1 port map( C1 => n4505, C2 => n6209, A => n6208, B => n6207,
                           ZN => n6223);
   U563 : OAI22_X1 port map( A1 => n4245, A2 => n6219, B1 => n4244, B2 => n6223
                           , ZN => n6211);
   U564 : OAI22_X1 port map( A1 => n4472, A2 => n6220, B1 => n4101, B2 => n6228
                           , ZN => n6210);
   U565 : AOI211_X1 port map( C1 => n4473, C2 => n6225, A => n6211, B => n6210,
                           ZN => n6232);
   U566 : AOI22_X1 port map( A1 => n4505, A2 => n3817, B1 => n4469, B2 => n3819
                           , ZN => n6213);
   U567 : OAI222_X1 port map( A1 => n4521, A2 => n3926, B1 => n4483, B2 => 
                           n4467, C1 => n4470, C2 => n4482, ZN => n6273);
   U568 : AOI22_X1 port map( A1 => n4480, A2 => n6239, B1 => n7721, B2 => n6273
                           , ZN => n6212);
   U569 : OAI211_X1 port map( C1 => n4519, C2 => n3816, A => n6213, B => n6212,
                           ZN => n6295);
   U570 : AOI22_X1 port map( A1 => n4474, A2 => n3817, B1 => n4480, B2 => n3819
                           , ZN => n6215);
   U571 : AOI22_X1 port map( A1 => n4289, A2 => n6239, B1 => n4103, B2 => n6273
                           , ZN => n6214);
   U572 : OAI211_X1 port map( C1 => n4290, C2 => n6216, A => n6215, B => n6214,
                           ZN => n6270);
   U573 : INV_X1 port map( A => n6270, ZN => n6248);
   U574 : OAI22_X1 port map( A1 => n4101, A2 => n6219, B1 => n6248, B2 => n7755
                           , ZN => n6218);
   U575 : OAI22_X1 port map( A1 => n6223, A2 => n7759, B1 => n6228, B2 => n7734
                           , ZN => n6217);
   U576 : AOI211_X1 port map( C1 => n4466, C2 => n6295, A => n6218, B => n6217,
                           ZN => n6236);
   U577 : OAI22_X1 port map( A1 => n6223, A2 => n7719, B1 => n6219, B2 => n7755
                           , ZN => n6222);
   U578 : OAI22_X1 port map( A1 => n4476, A2 => n6220, B1 => n6228, B2 => n7759
                           , ZN => n6221);
   U579 : AOI211_X1 port map( C1 => n4475, C2 => n6270, A => n6222, B => n6221,
                           ZN => n6249);
   U580 : OAI222_X1 port map( A1 => n4512, A2 => n6232, B1 => n4506, B2 => 
                           n6236, C1 => n4248, C2 => n6249, ZN => n6305);
   U581 : INV_X1 port map( A => n6223, ZN => n6245);
   U582 : AOI22_X1 port map( A1 => n4475, A2 => n6245, B1 => n7756, B2 => n6224
                           , ZN => n6227);
   U583 : AOI22_X1 port map( A1 => n4471, A2 => n6225, B1 => n4473, B2 => n7017
                           , ZN => n6226);
   U584 : OAI211_X1 port map( C1 => n6228, C2 => n7755, A => n6227, B => n6226,
                           ZN => n6230);
   U585 : INV_X1 port map( A => n6230, ZN => n6231);
   U586 : OAI222_X1 port map( A1 => n4248, A2 => n6232, B1 => n6231, B2 => 
                           n4512, C1 => n6249, C2 => n4506, ZN => n7117);
   U587 : AOI22_X1 port map( A1 => n4112, A2 => n6305, B1 => n4454, B2 => n7117
                           , ZN => n6235);
   U588 : AOI222_X1 port map( A1 => n7042, A2 => n4256, B1 => n6230, B2 => 
                           n4455, C1 => n6229, C2 => n4456, ZN => n6254);
   U589 : INV_X1 port map( A => n6254, ZN => n7118);
   U590 : OAI222_X1 port map( A1 => n4512, A2 => n6233, B1 => n4506, B2 => 
                           n6232, C1 => n4248, C2 => n6231, ZN => n7116);
   U591 : AOI22_X1 port map( A1 => n4453, A2 => n7118, B1 => n4114, B2 => n7116
                           , ZN => n6234);
   U592 : OAI211_X1 port map( C1 => n4462, C2 => n7082, A => n6235, B => n6234,
                           ZN => n6311);
   U593 : INV_X1 port map( A => n6311, ZN => n7148);
   U594 : INV_X1 port map( A => n6236, ZN => n6250);
   U595 : AOI222_X1 port map( A1 => n4498, A2 => n4465, B1 => n4099, B2 => 
                           n4516, C1 => n4109, C2 => n3922, ZN => n6351);
   U596 : AOI222_X1 port map( A1 => n4517, A2 => n3923, B1 => n4498, B2 => 
                           n4099, C1 => n4465, C2 => n4109, ZN => n6323);
   U597 : INV_X1 port map( A => n6323, ZN => n6300);
   U598 : AOI22_X1 port map( A1 => n6300, A2 => n7721, B1 => n7735, B2 => n7773
                           , ZN => n6238);
   U599 : AOI22_X1 port map( A1 => n4505, A2 => n6239, B1 => n6273, B2 => n7764
                           , ZN => n6237);
   U600 : OAI211_X1 port map( C1 => n6351, C2 => n4519, A => n6238, B => n6237,
                           ZN => n6327);
   U601 : INV_X1 port map( A => n6327, ZN => n6354);
   U602 : AOI22_X1 port map( A1 => n4471, A2 => n6270, B1 => n7756, B2 => n6295
                           , ZN => n6243);
   U603 : AOI22_X1 port map( A1 => n3819, A2 => n4505, B1 => n7721, B2 => n7773
                           , ZN => n6241);
   U604 : AOI22_X1 port map( A1 => n4469, A2 => n6239, B1 => n4480, B2 => n6273
                           , ZN => n6240);
   U605 : OAI211_X1 port map( C1 => n6323, C2 => n7725, A => n6241, B => n6240,
                           ZN => n6321);
   U606 : AOI22_X1 port map( A1 => n4518, A2 => n6321, B1 => n4473, B2 => n6244
                           , ZN => n6242);
   U607 : OAI211_X1 port map( C1 => n4245, C2 => n6354, A => n6243, B => n6242,
                           ZN => n6303);
   U608 : AOI22_X1 port map( A1 => n6295, A2 => n4518, B1 => n6244, B2 => n4243
                           , ZN => n6247);
   U609 : AOI22_X1 port map( A1 => n6321, A2 => n4475, B1 => n7761, B2 => n6245
                           , ZN => n6246);
   U610 : OAI211_X1 port map( C1 => n7719, C2 => n6248, A => n6247, B => n6246,
                           ZN => n6277);
   U611 : AOI222_X1 port map( A1 => n7731, A2 => n6250, B1 => n7757, B2 => 
                           n6303, C1 => n7724, C2 => n6277, ZN => n6304);
   U612 : INV_X1 port map( A => n7117, ZN => n6278);
   U613 : OAI22_X1 port map( A1 => n4464, A2 => n6304, B1 => n4234, B2 => n6278
                           , ZN => n6253);
   U614 : INV_X1 port map( A => n6305, ZN => n6269);
   U615 : INV_X1 port map( A => n6249, ZN => n6251);
   U616 : AOI222_X1 port map( A1 => n7731, A2 => n6251, B1 => n7757, B2 => 
                           n6277, C1 => n7724, C2 => n6250, ZN => n6308);
   U617 : OAI22_X1 port map( A1 => n4463, A2 => n6269, B1 => n6308, B2 => n4235
                           , ZN => n6252);
   U618 : AOI211_X1 port map( C1 => n4249, C2 => n7116, A => n6253, B => n6252,
                           ZN => n6362);
   U619 : OAI22_X1 port map( A1 => n6308, A2 => n7738, B1 => n6278, B2 => n7802
                           , ZN => n6256);
   U620 : OAI22_X1 port map( A1 => n4462, A2 => n6254, B1 => n6269, B2 => n7801
                           , ZN => n6255);
   U621 : AOI211_X1 port map( C1 => n4453, C2 => n7116, A => n6256, B => n6255,
                           ZN => n7149);
   U622 : OAI222_X1 port map( A1 => n4460, A2 => n7148, B1 => n4507, B2 => 
                           n6362, C1 => n4098, C2 => n7149, ZN => n6257);
   U623 : AOI211_X1 port map( C1 => n4508, C2 => n6257, A => n3920, B => n3919,
                           ZN => n6263);
   U624 : OAI222_X1 port map( A1 => n4521, A2 => n3915, B1 => n4483, B2 => 
                           n3917, C1 => n4495, C2 => n3916, ZN => n6718);
   U625 : INV_X1 port map( A => n6718, ZN => n6761);
   U626 : OAI222_X1 port map( A1 => n4521, A2 => n3913, B1 => n4483, B2 => 
                           n3914, C1 => n4495, C2 => n4448, ZN => n6764);
   U627 : INV_X1 port map( A => n6764, ZN => n6293);
   U628 : OAI22_X1 port map( A1 => n4519, A2 => n6761, B1 => n4102, B2 => n6293
                           , ZN => n6261);
   U629 : OAI22_X1 port map( A1 => n4521, A2 => n4448, B1 => n4504, B2 => n3915
                           , ZN => n6258);
   U630 : INV_X1 port map( A => n6258, ZN => n6259);
   U631 : OAI21_X1 port map( B1 => n4482, B2 => n3914, A => n6259, ZN => n6713)
                           ;
   U632 : INV_X1 port map( A => n6713, ZN => n6760);
   U633 : OAI222_X1 port map( A1 => n4521, A2 => n3914, B1 => n4483, B2 => 
                           n3916, C1 => n4495, C2 => n3915, ZN => n6714);
   U634 : INV_X1 port map( A => n6714, ZN => n6758);
   U635 : OAI22_X1 port map( A1 => n4478, A2 => n6760, B1 => n4477, B2 => n6758
                           , ZN => n6260);
   U636 : OAI21_X1 port map( B1 => n6261, B2 => n6260, A => n4447, ZN => n6262)
                           ;
   U637 : NAND4_X1 port map( A1 => n3932, A2 => n3918, A3 => n6263, A4 => n6262
                           , ZN => OUTALU(9));
   U638 : AOI22_X1 port map( A1 => DATA1(9), A2 => n7825, B1 => DATA1(12), B2 
                           => n7709, ZN => n6266);
   U639 : NAND2_X1 port map( A1 => DATA1(11), A2 => n7824, ZN => n6478);
   U640 : NAND2_X1 port map( A1 => DATA1(10), A2 => n7828, ZN => n6265);
   U641 : NAND4_X1 port map( A1 => n6266, A2 => n6478, A3 => n6265, A4 => n6264
                           , ZN => n1334);
   U642 : INV_X1 port map( A => DATA2(8), ZN => n7369);
   U643 : AOI22_X1 port map( A1 => DATA1(8), A2 => DATA2(8), B1 => n7369, B2 =>
                           n7191, ZN => n7238);
   U644 : AOI22_X1 port map( A1 => n4270, A2 => n7823, B1 => n7821, B2 => n7238
                           , ZN => n1278);
   U645 : NAND3_X1 port map( A1 => DATA2(8), A2 => DATA1(8), A3 => n7105, ZN =>
                           n1277);
   U646 : OAI222_X1 port map( A1 => n7732, A2 => n6760, B1 => n7725, B2 => 
                           n6758, C1 => n7763, C2 => n6293, ZN => n6268);
   U647 : OAI22_X1 port map( A1 => n4446, A2 => n4451, B1 => n4095, B2 => n4225
                           , ZN => n6267);
   U648 : AOI21_X1 port map( B1 => n7798, B2 => n6268, A => n6267, ZN => n6284)
                           ;
   U649 : OAI22_X1 port map( A1 => n4460, A2 => n7149, B1 => n4098, B2 => n6362
                           , ZN => n6282);
   U650 : INV_X1 port map( A => n6308, ZN => n6331);
   U651 : OAI22_X1 port map( A1 => n4234, A2 => n6269, B1 => n6304, B2 => n4235
                           , ZN => n6280);
   U652 : AOI22_X1 port map( A1 => n4471, A2 => n6295, B1 => n4473, B2 => n6270
                           , ZN => n6276);
   U653 : AOI222_X1 port map( A1 => n4517, A2 => n4465, B1 => n4498, B2 => 
                           n3922, C1 => n4109, C2 => n3912, ZN => n6380);
   U654 : OAI22_X1 port map( A1 => n6380, A2 => n4519, B1 => n3816, B2 => n4102
                           , ZN => n6272);
   U655 : OAI22_X1 port map( A1 => n6323, A2 => n4478, B1 => n6351, B2 => n4477
                           , ZN => n6271);
   U656 : AOI211_X1 port map( C1 => n4505, C2 => n6273, A => n6272, B => n6271,
                           ZN => n6381);
   U657 : INV_X1 port map( A => n6381, ZN => n6274);
   U658 : AOI22_X1 port map( A1 => n4468, A2 => n6321, B1 => n4475, B2 => n6274
                           , ZN => n6275);
   U659 : OAI211_X1 port map( C1 => n6354, C2 => n4244, A => n6276, B => n6275,
                           ZN => n6330);
   U660 : AOI222_X1 port map( A1 => n7731, A2 => n6277, B1 => n7757, B2 => 
                           n6330, C1 => n7724, C2 => n6303, ZN => n6388);
   U661 : OAI22_X1 port map( A1 => n4462, A2 => n6278, B1 => n6388, B2 => n4464
                           , ZN => n6279);
   U662 : AOI211_X1 port map( C1 => n4114, C2 => n6331, A => n6280, B => n6279,
                           ZN => n6389);
   U663 : OAI22_X1 port map( A1 => n4094, A2 => n7148, B1 => n4507, B2 => n6389
                           , ZN => n6281);
   U664 : OAI21_X1 port map( B1 => n6282, B2 => n6281, A => n4508, ZN => n6283)
                           ;
   U665 : NAND4_X1 port map( A1 => n3911, A2 => n3910, A3 => n6284, A4 => n6283
                           , ZN => OUTALU(8));
   U666 : OAI221_X1 port map( B1 => DATA1(7), B2 => n7161, C1 => n7174, C2 => 
                           n7158, A => n7143, ZN => n1286);
   U667 : NAND2_X1 port map( A1 => DATA1(7), A2 => n1946, ZN => n7192);
   U668 : INV_X1 port map( A => n7192, ZN => n7220);
   U669 : AOI22_X1 port map( A1 => n7220, A2 => n7821, B1 => n7823, B2 => n4020
                           , ZN => n1324);
   U670 : AOI21_X1 port map( B1 => n5990, B2 => n6347, A => n6285, ZN => n6320)
                           ;
   U671 : OAI21_X1 port map( B1 => n6320, B2 => n1353, A => n6286, ZN => n6291)
                           ;
   U672 : AOI21_X1 port map( B1 => n5990, B2 => n6346, A => n6285, ZN => n6319)
                           ;
   U673 : OAI21_X1 port map( B1 => n6319, B2 => n1353, A => n6286, ZN => n6290)
                           ;
   U674 : OAI22_X1 port map( A1 => n1896, A2 => n6291, B1 => n7162, B2 => n6290
                           , ZN => n1321);
   U675 : NOR2_X1 port map( A1 => n7688, A2 => n7125, ZN => n6482);
   U676 : NOR2_X1 port map( A1 => n6402, A2 => n7708, ZN => n6287);
   U677 : AOI211_X1 port map( C1 => n7825, C2 => DATA1(8), A => n6482, B => 
                           n6287, ZN => n6289);
   U678 : NAND2_X1 port map( A1 => DATA1(10), A2 => n7824, ZN => n6288);
   U679 : OAI211_X1 port map( C1 => n7707, C2 => n7174, A => n6289, B => n6288,
                           ZN => n1366);
   U680 : AOI22_X1 port map( A1 => n7166, A2 => n6291, B1 => n6808, B2 => n6290
                           , ZN => n6292);
   U681 : NOR2_X1 port map( A1 => n1322, A2 => n6292, ZN => n1319);
   U682 : AOI22_X1 port map( A1 => n3908, A2 => n4228, B1 => n3823, B2 => n4525
                           , ZN => n6314);
   U683 : OAI22_X1 port map( A1 => n4477, A2 => n6293, B1 => n4519, B2 => n6760
                           , ZN => n6294);
   U684 : AOI211_X1 port map( C1 => n4447, C2 => n6294, A => n4220, B => n7819,
                           ZN => n6313);
   U685 : AOI22_X1 port map( A1 => n4471, A2 => n6321, B1 => n7761, B2 => n6295
                           , ZN => n6302);
   U686 : AOI22_X1 port map( A1 => n4498, A2 => n3912, B1 => n3907, B2 => n4485
                           , ZN => n6296);
   U687 : INV_X1 port map( A => n6296, ZN => n6297);
   U688 : AOI21_X1 port map( B1 => n4517, B2 => n3922, A => n6297, ZN => n6377)
                           ;
   U689 : OAI22_X1 port map( A1 => n4519, A2 => n6377, B1 => n3816, B2 => n4290
                           , ZN => n6299);
   U690 : OAI22_X1 port map( A1 => n4478, A2 => n6351, B1 => n4477, B2 => n6380
                           , ZN => n6298);
   U691 : AOI211_X1 port map( C1 => n4474, C2 => n6300, A => n6299, B => n6298,
                           ZN => n6422);
   U692 : INV_X1 port map( A => n6422, ZN => n6357);
   U693 : AOI22_X1 port map( A1 => n6357, A2 => n7739, B1 => n7756, B2 => n6327
                           , ZN => n6301);
   U694 : OAI211_X1 port map( C1 => n6381, C2 => n4244, A => n6302, B => n6301,
                           ZN => n6358);
   U695 : AOI222_X1 port map( A1 => n7724, A2 => n6330, B1 => n6303, B2 => 
                           n7731, C1 => n6358, C2 => n7757, ZN => n6361);
   U696 : INV_X1 port map( A => n6361, ZN => n6417);
   U697 : INV_X1 port map( A => n6304, ZN => n6348);
   U698 : AOI22_X1 port map( A1 => n4112, A2 => n6417, B1 => n4114, B2 => n6348
                           , ZN => n6307);
   U699 : INV_X1 port map( A => n6388, ZN => n6349);
   U700 : AOI22_X1 port map( A1 => n4454, A2 => n6349, B1 => n4249, B2 => n6305
                           , ZN => n6306);
   U701 : OAI211_X1 port map( C1 => n4234, C2 => n6308, A => n6307, B => n6306,
                           ZN => n6430);
   U702 : INV_X1 port map( A => n6430, ZN => n6390);
   U703 : OAI22_X1 port map( A1 => n6390, A2 => n4507, B1 => n6389, B2 => n4098
                           , ZN => n6310);
   U704 : OAI22_X1 port map( A1 => n4460, A2 => n6362, B1 => n4094, B2 => n7149
                           , ZN => n6309);
   U705 : AOI211_X1 port map( C1 => n4461, C2 => n6311, A => n6310, B => n6309,
                           ZN => n6365);
   U706 : OR3_X1 port map( A1 => n4113, A2 => n6365, A3 => n4251, ZN => n6312);
   U707 : NAND3_X1 port map( A1 => n6314, A2 => n6313, A3 => n6312, ZN => 
                           OUTALU(7));
   U708 : AOI22_X1 port map( A1 => n7166, A2 => n6320, B1 => n6808, B2 => n6319
                           , ZN => n1354);
   U709 : INV_X1 port map( A => DATA2(6), ZN => n7372);
   U710 : AOI22_X1 port map( A1 => DATA1(6), A2 => n7372, B1 => DATA2(6), B2 =>
                           n7175, ZN => n7235);
   U711 : AOI21_X1 port map( B1 => n1901, B2 => DATA1(6), A => n1900, ZN => 
                           n6315);
   U712 : OAI22_X1 port map( A1 => n7235, A2 => n7161, B1 => n6315, B2 => n7372
                           , ZN => n1328);
   U713 : NOR2_X1 port map( A1 => n7688, A2 => n7167, ZN => n6316);
   U714 : NOR2_X1 port map( A1 => n7191, A2 => n7708, ZN => n6495);
   U715 : AOI211_X1 port map( C1 => n7826, C2 => DATA1(7), A => n6316, B => 
                           n6495, ZN => n6318);
   U716 : OAI211_X1 port map( C1 => n7711, C2 => n6402, A => n6318, B => n6317,
                           ZN => n1403);
   U717 : OAI22_X1 port map( A1 => n6320, A2 => n1896, B1 => n6319, B2 => n7162
                           , ZN => n1349);
   U718 : NAND2_X1 port map( A1 => n7760, A2 => n6764, ZN => n6338);
   U719 : AOI22_X1 port map( A1 => n4473, A2 => n6321, B1 => n6357, B2 => n7765
                           , ZN => n6329);
   U720 : AOI22_X1 port map( A1 => n4109, A2 => n4093, B1 => n3907, B2 => n3931
                           , ZN => n6322);
   U721 : OAI21_X1 port map( B1 => n7741, B2 => n7787, A => n6322, ZN => n6376)
                           ;
   U722 : OAI22_X1 port map( A1 => n6351, A2 => n4102, B1 => n6323, B2 => n7770
                           , ZN => n6325);
   U723 : OAI22_X1 port map( A1 => n4478, A2 => n6380, B1 => n4477, B2 => n6377
                           , ZN => n6324);
   U724 : AOI211_X1 port map( C1 => n7760, C2 => n6376, A => n6325, B => n6324,
                           ZN => n6820);
   U725 : INV_X1 port map( A => n6820, ZN => n6326);
   U726 : AOI22_X1 port map( A1 => n7727, A2 => n6327, B1 => n7739, B2 => n6326
                           , ZN => n6328);
   U727 : OAI211_X1 port map( C1 => n6381, C2 => n4101, A => n6329, B => n6328,
                           ZN => n6384);
   U728 : AOI222_X1 port map( A1 => n7724, A2 => n6358, B1 => n6330, B2 => 
                           n7731, C1 => n6384, C2 => n7757, ZN => n6825);
   U729 : INV_X1 port map( A => n6825, ZN => n6418);
   U730 : AOI22_X1 port map( A1 => n4112, A2 => n6418, B1 => n4453, B2 => n6348
                           , ZN => n6333);
   U731 : AOI22_X1 port map( A1 => n4114, A2 => n6349, B1 => n4249, B2 => n6331
                           , ZN => n6332);
   U732 : OAI211_X1 port map( C1 => n6361, C2 => n4235, A => n6333, B => n6332,
                           ZN => n6814);
   U733 : INV_X1 port map( A => n6814, ZN => n6391);
   U734 : OAI22_X1 port map( A1 => n6391, A2 => n4507, B1 => n7149, B2 => n7808
                           , ZN => n6335);
   U735 : OAI22_X1 port map( A1 => n4460, A2 => n6389, B1 => n4094, B2 => n6362
                           , ZN => n6334);
   U736 : AOI211_X1 port map( C1 => n6430, C2 => n7800, A => n6335, B => n6334,
                           ZN => n6394);
   U737 : OAI22_X1 port map( A1 => n4113, A2 => n6394, B1 => n4443, B2 => n6365
                           , ZN => n6336);
   U738 : INV_X1 port map( A => n6336, ZN => n6337);
   U739 : OAI22_X1 port map( A1 => n4222, A2 => n6338, B1 => n6337, B2 => n7748
                           , ZN => n6339);
   U740 : AOI211_X1 port map( C1 => n4274, C2 => n4510, A => n3904, B => n6339,
                           ZN => n6341);
   U741 : NAND2_X1 port map( A1 => n4096, A2 => n3903, ZN => n6340);
   U742 : OAI211_X1 port map( C1 => n4096, C2 => n3905, A => n6341, B => n6340,
                           ZN => OUTALU(6));
   U743 : NOR2_X1 port map( A1 => n6806, A2 => n7707, ZN => n6403);
   U744 : NAND2_X1 port map( A1 => DATA1(3), A2 => n7828, ZN => n6967);
   U745 : NAND2_X1 port map( A1 => DATA1(4), A2 => n7826, ZN => n6412);
   U746 : OAI211_X1 port map( C1 => n7688, C2 => n1939, A => n6967, B => n6412,
                           ZN => n6342);
   U747 : AOI211_X1 port map( C1 => n7824, C2 => DATA1(2), A => n6403, B => 
                           n6342, ZN => n1937);
   U748 : NOR2_X1 port map( A1 => n7227, A2 => n7708, ZN => n7680);
   U749 : NAND2_X1 port map( A1 => DATA1(3), A2 => n7826, ZN => n6804);
   U750 : NAND2_X1 port map( A1 => DATA1(4), A2 => n7692, ZN => n6408);
   U751 : OAI211_X1 port map( C1 => n7711, C2 => n1939, A => n6804, B => n6408,
                           ZN => n6343);
   U752 : AOI211_X1 port map( C1 => DATA1(0), C2 => n7709, A => n7680, B => 
                           n6343, ZN => n1394);
   U753 : OAI21_X1 port map( B1 => n7158, B2 => n6806, A => n7143, ZN => n6345)
                           ;
   U754 : OAI22_X1 port map( A1 => n1937, A2 => n1952, B1 => n1394, B2 => n1958
                           , ZN => n6344);
   U755 : AOI22_X1 port map( A1 => DATA2(5), A2 => n6345, B1 => n1902, B2 => 
                           n6344, ZN => n1393);
   U756 : NAND2_X1 port map( A1 => DATA1(5), A2 => n7373, ZN => n7231);
   U757 : NAND2_X1 port map( A1 => DATA2(5), A2 => n6806, ZN => n7234);
   U758 : NAND2_X1 port map( A1 => n7231, A2 => n7234, ZN => n2519_port);
   U759 : AOI22_X1 port map( A1 => n7821, A2 => n2519_port, B1 => n7823, B2 => 
                           n4027, ZN => n1392);
   U760 : OAI22_X1 port map( A1 => n1896, A2 => n6347, B1 => n7162, B2 => n6346
                           , ZN => n1389);
   U761 : AOI22_X1 port map( A1 => n3899, A2 => n4452, B1 => n4442, B2 => n4227
                           , ZN => n6367);
   U762 : AOI22_X1 port map( A1 => n4453, A2 => n6349, B1 => n4249, B2 => n6348
                           , ZN => n6360);
   U763 : AOI22_X1 port map( A1 => n4498, A2 => n4093, B1 => n4485, B2 => n3898
                           , ZN => n6350);
   U764 : OAI21_X1 port map( B1 => n7741, B2 => n7786, A => n6350, ZN => n6818)
                           ;
   U765 : INV_X1 port map( A => n6376, ZN => n6815);
   U766 : OAI22_X1 port map( A1 => n6815, A2 => n7732, B1 => n4478, B2 => n6377
                           , ZN => n6353);
   U767 : OAI22_X1 port map( A1 => n6351, A2 => n4290, B1 => n6380, B2 => n4102
                           , ZN => n6352);
   U768 : AOI211_X1 port map( C1 => n7760, C2 => n6818, A => n6353, B => n6352,
                           ZN => n6980);
   U769 : OAI22_X1 port map( A1 => n4245, A2 => n6980, B1 => n6820, B2 => n4244
                           , ZN => n6356);
   U770 : OAI22_X1 port map( A1 => n7766, A2 => n6381, B1 => n4476, B2 => n6354
                           , ZN => n6355);
   U771 : AOI211_X1 port map( C1 => n6357, C2 => n7756, A => n6356, B => n6355,
                           ZN => n6425);
   U772 : INV_X1 port map( A => n6425, ZN => n6385);
   U773 : AOI222_X1 port map( A1 => n7724, A2 => n6384, B1 => n6358, B2 => 
                           n7731, C1 => n6385, C2 => n7757, ZN => n6826);
   U774 : INV_X1 port map( A => n6826, ZN => n6985);
   U775 : AOI22_X1 port map( A1 => n4112, A2 => n6985, B1 => n4454, B2 => n6418
                           , ZN => n6359);
   U776 : OAI211_X1 port map( C1 => n4463, C2 => n6361, A => n6360, B => n6359,
                           ZN => n6975);
   U777 : OAI22_X1 port map( A1 => n6391, A2 => n4098, B1 => n6390, B2 => n7799
                           , ZN => n6364);
   U778 : OAI22_X1 port map( A1 => n4250, A2 => n6362, B1 => n4094, B2 => n6389
                           , ZN => n6363);
   U779 : AOI211_X1 port map( C1 => n6975, C2 => n7804, A => n6364, B => n6363,
                           ZN => n6433);
   U780 : OAI222_X1 port map( A1 => n4113, A2 => n6433, B1 => n4445, B2 => 
                           n6365, C1 => n4443, C2 => n6394, ZN => n6993);
   U781 : INV_X1 port map( A => n6993, ZN => n6812);
   U782 : OR3_X1 port map( A1 => n6812, A2 => n4441, A3 => n4251, ZN => n6366);
   U783 : NAND4_X1 port map( A1 => n3902, A2 => n3900, A3 => n6367, A4 => n6366
                           , ZN => OUTALU(5));
   U784 : AOI22_X1 port map( A1 => n7166, A2 => n6374, B1 => n6808, B2 => n6373
                           , ZN => n1430);
   U785 : INV_X1 port map( A => n1902, ZN => n6368);
   U786 : NOR3_X1 port map( A1 => n1394, A2 => n6368, A3 => n1952, ZN => n6372)
                           ;
   U787 : NAND2_X1 port map( A1 => DATA2(4), A2 => n7183, ZN => n7228);
   U788 : OAI21_X1 port map( B1 => n7183, B2 => DATA2(4), A => n7228, ZN => 
                           n6369);
   U789 : INV_X1 port map( A => n6369, ZN => n7176);
   U790 : AOI21_X1 port map( B1 => n1901, B2 => DATA1(4), A => n1900, ZN => 
                           n6370);
   U791 : INV_X1 port map( A => DATA2(4), ZN => n7675);
   U792 : OAI22_X1 port map( A1 => n7176, A2 => n7161, B1 => n6370, B2 => n7675
                           , ZN => n6371);
   U793 : AOI211_X1 port map( C1 => n7823, C2 => n4280, A => n6372, B => n6371,
                           ZN => n1428);
   U794 : OAI22_X1 port map( A1 => n6374, A2 => n1896, B1 => n6373, B2 => n7162
                           , ZN => n1425);
   U795 : AOI22_X1 port map( A1 => n6418, A2 => n7723, B1 => n6417, B2 => n7733
                           , ZN => n6387);
   U796 : AOI22_X1 port map( A1 => n4498, A2 => n3898, B1 => n4438, B2 => n4108
                           , ZN => n6375);
   U797 : OAI21_X1 port map( B1 => n7741, B2 => n7789, A => n6375, ZN => n7283)
                           ;
   U798 : AOI22_X1 port map( A1 => n4103, A2 => n7283, B1 => n4480, B2 => n6376
                           , ZN => n6379);
   U799 : INV_X1 port map( A => n6377, ZN => n6421);
   U800 : AOI22_X1 port map( A1 => n7721, A2 => n6818, B1 => n6421, B2 => n7764
                           , ZN => n6378);
   U801 : OAI211_X1 port map( C1 => n6380, C2 => n4290, A => n6379, B => n6378,
                           ZN => n7290);
   U802 : OAI22_X1 port map( A1 => n6820, A2 => n4101, B1 => n6980, B2 => n7755
                           , ZN => n6383);
   U803 : OAI22_X1 port map( A1 => n6422, A2 => n4472, B1 => n6381, B2 => n4476
                           , ZN => n6382);
   U804 : AOI211_X1 port map( C1 => n7739, C2 => n7290, A => n6383, B => n6382,
                           ZN => n6824);
   U805 : INV_X1 port map( A => n6824, ZN => n6427);
   U806 : AOI222_X1 port map( A1 => n7724, A2 => n6385, B1 => n6384, B2 => 
                           n7731, C1 => n7757, C2 => n6427, ZN => n6988);
   U807 : INV_X1 port map( A => n6988, ZN => n7296);
   U808 : AOI22_X1 port map( A1 => n4454, A2 => n6985, B1 => n7296, B2 => n7736
                           , ZN => n6386);
   U809 : OAI211_X1 port map( C1 => n4462, C2 => n6388, A => n6387, B => n6386,
                           ZN => n7278);
   U810 : INV_X1 port map( A => n7278, ZN => n6832);
   U811 : OAI22_X1 port map( A1 => n6832, A2 => n4507, B1 => n4250, B2 => n6389
                           , ZN => n6393);
   U812 : OAI22_X1 port map( A1 => n6391, A2 => n4460, B1 => n6390, B2 => n4094
                           , ZN => n6392);
   U813 : AOI211_X1 port map( C1 => n4439, C2 => n6975, A => n6393, B => n6392,
                           ZN => n6434);
   U814 : OAI222_X1 port map( A1 => n4113, A2 => n6434, B1 => n4445, B2 => 
                           n6394, C1 => n4443, C2 => n6433, ZN => n7313);
   U815 : INV_X1 port map( A => n7313, ZN => n6813);
   U816 : OAI22_X1 port map( A1 => n6813, A2 => n4441, B1 => n6812, B2 => n4440
                           , ZN => n6395);
   U817 : AOI22_X1 port map( A1 => n4508, A2 => n6395, B1 => n3895, B2 => n4097
                           , ZN => n6396);
   U818 : OAI211_X1 port map( C1 => n4097, C2 => n3897, A => n3896, B => n6396,
                           ZN => OUTALU(4));
   U819 : NAND2_X1 port map( A1 => DATA1(3), A2 => n7661, ZN => n7226);
   U820 : NOR2_X1 port map( A1 => DATA1(3), A2 => n7661, ZN => n7233);
   U821 : INV_X1 port map( A => n7233, ZN => n6397);
   U822 : NAND2_X1 port map( A1 => n7226, A2 => n6397, ZN => n7173);
   U823 : NOR2_X1 port map( A1 => n7227, A2 => n7696, ZN => n6966);
   U824 : AOI21_X1 port map( B1 => n7824, B2 => DATA1(0), A => n6966, ZN => 
                           n6398);
   U825 : NAND2_X1 port map( A1 => DATA1(3), A2 => n7827, ZN => n6411);
   U826 : OAI211_X1 port map( C1 => n7708, C2 => n1939, A => n6398, B => n6411,
                           ZN => n6399);
   U827 : AOI22_X1 port map( A1 => n7821, A2 => n7173, B1 => n1902, B2 => n6399
                           , ZN => n1470);
   U828 : OAI21_X1 port map( B1 => n7158, B2 => n6400, A => n7143, ZN => n6401)
                           ;
   U829 : AOI22_X1 port map( A1 => DATA2(3), A2 => n6401, B1 => n7823, B2 => 
                           n4048, ZN => n1469);
   U830 : NOR2_X1 port map( A1 => n7688, A2 => n6402, ZN => n6487);
   U831 : AOI211_X1 port map( C1 => n7824, C2 => DATA1(8), A => n6403, B => 
                           n6487, ZN => n6405);
   U832 : OAI211_X1 port map( C1 => n7708, C2 => n7174, A => n6405, B => n6404,
                           ZN => n1441);
   U833 : AOI211_X1 port map( C1 => n7826, C2 => DATA1(5), A => n6407, B => 
                           n6406, ZN => n6409);
   U834 : OAI211_X1 port map( C1 => n7711, C2 => n7174, A => n6409, B => n6408,
                           ZN => n1936);
   U835 : INV_X1 port map( A => n1958, ZN => n6970);
   U836 : AOI22_X1 port map( A1 => DATA1(6), A2 => n7824, B1 => DATA1(5), B2 =>
                           n7691, ZN => n6413);
   U837 : NAND4_X1 port map( A1 => n6413, A2 => n6412, A3 => n6411, A4 => n6410
                           , ZN => n6971);
   U838 : AOI222_X1 port map( A1 => n1441, A2 => n1068, B1 => n1936, B2 => 
                           n6970, C1 => n6971, C2 => n6969, ZN => n2445);
   U839 : AOI21_X1 port map( B1 => n7713, B2 => n6415, A => n6414, ZN => n6416)
                           ;
   U840 : NAND2_X1 port map( A1 => n6808, A2 => n6416, ZN => n1467);
   U841 : AOI22_X1 port map( A1 => n4453, A2 => n6418, B1 => n7794, B2 => n6417
                           , ZN => n6429);
   U842 : INV_X1 port map( A => n6818, ZN => n6977);
   U843 : OAI22_X1 port map( A1 => n4478, A2 => n6977, B1 => n4519, B2 => n3815
                           , ZN => n6420);
   U844 : INV_X1 port map( A => n7283, ZN => n6976);
   U845 : OAI22_X1 port map( A1 => n7732, A2 => n6976, B1 => n4102, B2 => n6815
                           , ZN => n6419);
   U846 : AOI211_X1 port map( C1 => n6421, C2 => n7740, A => n6420, B => n6419,
                           ZN => n7287);
   U847 : OAI22_X1 port map( A1 => n4245, A2 => n7287, B1 => n4101, B2 => n6980
                           , ZN => n6424);
   U848 : OAI22_X1 port map( A1 => n6422, A2 => n4476, B1 => n4472, B2 => n6820
                           , ZN => n6423);
   U849 : AOI211_X1 port map( C1 => n4518, C2 => n7290, A => n6424, B => n6423,
                           ZN => n6983);
   U850 : OAI22_X1 port map( A1 => n4512, A2 => n6425, B1 => n4506, B2 => n6983
                           , ZN => n6426);
   U851 : AOI21_X1 port map( B1 => n6427, B2 => n7724, A => n6426, ZN => n7300)
                           ;
   U852 : INV_X1 port map( A => n7300, ZN => n6984);
   U853 : AOI22_X1 port map( A1 => n4112, A2 => n6984, B1 => n4454, B2 => n7296
                           , ZN => n6428);
   U854 : OAI211_X1 port map( C1 => n6826, C2 => n7802, A => n6429, B => n6428,
                           ZN => n7279);
   U855 : AOI22_X1 port map( A1 => n4110, A2 => n7279, B1 => n4436, B2 => n6814
                           , ZN => n6432);
   U856 : AOI22_X1 port map( A1 => n3921, A2 => n6975, B1 => n4461, B2 => n6430
                           , ZN => n6431);
   U857 : OAI211_X1 port map( C1 => n6832, C2 => n4098, A => n6432, B => n6431,
                           ZN => n6991);
   U858 : INV_X1 port map( A => n6433, ZN => n6435);
   U859 : INV_X1 port map( A => n6434, ZN => n6833);
   U860 : AOI222_X1 port map( A1 => n7728, A2 => n6991, B1 => n7797, B2 => 
                           n6435, C1 => n6833, C2 => n7747, ZN => n7312);
   U861 : OAI222_X1 port map( A1 => n6813, A2 => n4440, B1 => n6812, B2 => 
                           n4217, C1 => n7312, C2 => n4441, ZN => n6436);
   U862 : AOI22_X1 port map( A1 => n4508, A2 => n6436, B1 => n4216, B2 => n4221
                           , ZN => n6437);
   U863 : NAND4_X1 port map( A1 => n3893, A2 => n3892, A3 => n3894, A4 => n6437
                           , ZN => OUTALU(3));
   U864 : NOR2_X1 port map( A1 => n1921, A2 => n7711, ZN => n7700);
   U865 : OAI211_X1 port map( C1 => n7707, C2 => n1912, A => n6439, B => n6438,
                           ZN => n6440);
   U866 : AOI211_X1 port map( C1 => DATA1(20), C2 => n7709, A => n7700, B => 
                           n6440, ZN => n1550);
   U867 : NOR2_X1 port map( A1 => n1914, A2 => n7708, ZN => n6443);
   U868 : NAND2_X1 port map( A1 => DATA1(21), A2 => n7709, ZN => n6441);
   U869 : NAND2_X1 port map( A1 => DATA1(22), A2 => n7824, ZN => n7702);
   U870 : OAI211_X1 port map( C1 => n7707, C2 => n1911, A => n6441, B => n7702,
                           ZN => n6442);
   U871 : AOI211_X1 port map( C1 => n7826, C2 => DATA1(24), A => n6443, B => 
                           n6442, ZN => n1560);
   U872 : OAI21_X1 port map( B1 => n7374, B2 => n7661, A => n7664, ZN => n1949)
                           ;
   U873 : NOR3_X1 port map( A1 => n6444, A2 => n7678, A3 => n1949, ZN => n5992)
                           ;
   U874 : NAND2_X1 port map( A1 => DATA1(20), A2 => n7828, ZN => n7698);
   U875 : OAI211_X1 port map( C1 => n7688, C2 => n1925, A => n6445, B => n7698,
                           ZN => n6446);
   U876 : AOI211_X1 port map( C1 => DATA1(22), C2 => n7692, A => n6447, B => 
                           n6446, ZN => n1918);
   U877 : NAND2_X1 port map( A1 => DATA1(20), A2 => n7826, ZN => n7701);
   U878 : OAI211_X1 port map( C1 => n7688, C2 => n7027, A => n6448, B => n7701,
                           ZN => n6449);
   U879 : AOI211_X1 port map( C1 => n7828, C2 => DATA1(19), A => n6450, B => 
                           n6449, ZN => n6460);
   U880 : NAND2_X1 port map( A1 => DATA1(19), A2 => n7826, ZN => n7697);
   U881 : OAI211_X1 port map( C1 => n7688, C2 => n1929, A => n6451, B => n7697,
                           ZN => n6452);
   U882 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(20), A => n6453, B => 
                           n6452, ZN => n6469);
   U883 : OAI222_X1 port map( A1 => n1952, A2 => n1918, B1 => n1958, B2 => 
                           n6460, C1 => n6469, C2 => n6466, ZN => n1919);
   U884 : NAND2_X1 port map( A1 => DATA1(19), A2 => n7827, ZN => n7704);
   U885 : OAI211_X1 port map( C1 => n7688, C2 => n7695, A => n6454, B => n7704,
                           ZN => n6455);
   U886 : AOI211_X1 port map( C1 => n7828, C2 => DATA1(17), A => n6456, B => 
                           n6455, ZN => n6468);
   U887 : OAI222_X1 port map( A1 => n1958, A2 => n6469, B1 => n1952, B2 => 
                           n6460, C1 => n6468, C2 => n6466, ZN => n1920);
   U888 : AOI22_X1 port map( A1 => n5992, A2 => n1919, B1 => n1949, B2 => n1920
                           , ZN => n1531);
   U889 : NAND2_X1 port map( A1 => DATA1(21), A2 => n7828, ZN => n7703);
   U890 : OAI211_X1 port map( C1 => n7688, C2 => n7000, A => n6457, B => n7703,
                           ZN => n6458);
   U891 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(23), A => n6459, B => 
                           n6458, ZN => n1915);
   U892 : OAI222_X1 port map( A1 => n1958, A2 => n1918, B1 => n1952, B2 => 
                           n1915, C1 => n6460, C2 => n6466, ZN => n1916);
   U893 : AOI22_X1 port map( A1 => DATA1(14), A2 => n7824, B1 => DATA1(13), B2 
                           => n7709, ZN => n6464);
   U894 : NAND4_X1 port map( A1 => n6464, A2 => n6463, A3 => n6462, A4 => n6461
                           , ZN => n1928);
   U895 : AOI22_X1 port map( A1 => n6970, A2 => n1926, B1 => n1068, B2 => n1928
                           , ZN => n6465);
   U896 : OAI21_X1 port map( B1 => n6468, B2 => n1952, A => n6465, ZN => n1924)
                           ;
   U897 : INV_X1 port map( A => n1950, ZN => n6471);
   U898 : AOI22_X1 port map( A1 => n1949, A2 => n1924, B1 => n6471, B2 => n1916
                           , ZN => n1535);
   U899 : INV_X1 port map( A => n1926, ZN => n6467);
   U900 : OAI222_X1 port map( A1 => n1952, A2 => n6469, B1 => n1958, B2 => 
                           n6468, C1 => n6467, C2 => n6466, ZN => n1923);
   U901 : INV_X1 port map( A => n1951, ZN => n6470);
   U902 : AOI22_X1 port map( A1 => n5992, A2 => n1923, B1 => n6470, B2 => n1919
                           , ZN => n1534);
   U903 : AOI22_X1 port map( A1 => n5992, A2 => n1920, B1 => n1949, B2 => n1923
                           , ZN => n1537);
   U904 : INV_X1 port map( A => n1965, ZN => n6472);
   U905 : AOI22_X1 port map( A1 => n6472, A2 => n1923, B1 => n1919, B2 => n6471
                           , ZN => n1542);
   U906 : NAND2_X1 port map( A1 => DATA1(26), A2 => n7827, ZN => n1194);
   U907 : NAND2_X1 port map( A1 => DATA1(25), A2 => n7826, ZN => n1546);
   U908 : INV_X1 port map( A => DATA1(22), ZN => n7168);
   U909 : OAI211_X1 port map( C1 => n7688, C2 => n7168, A => n1194, B => n1546,
                           ZN => n6473);
   U910 : AOI211_X1 port map( C1 => n7691, C2 => DATA1(24), A => n6474, B => 
                           n6473, ZN => n1584);
   U911 : NAND2_X1 port map( A1 => n7692, A2 => DATA1(28), ZN => n2008);
   U912 : NAND2_X1 port map( A1 => n7825, A2 => DATA1(27), ZN => n1580);
   U913 : NAND2_X1 port map( A1 => DATA1(26), A2 => n7828, ZN => n1581);
   U914 : AOI21_X1 port map( B1 => DATA1(24), B2 => n7709, A => n6475, ZN => 
                           n6476);
   U915 : NAND4_X1 port map( A1 => n6476, A2 => n2008, A3 => n1581, A4 => n1580
                           , ZN => n1682);
   U916 : AOI21_X1 port map( B1 => n7824, B2 => DATA1(26), A => n6477, ZN => 
                           n1595);
   U917 : AOI22_X1 port map( A1 => DATA1(10), A2 => n7709, B1 => DATA1(12), B2 
                           => n7828, ZN => n6481);
   U918 : NAND4_X1 port map( A1 => n6481, A2 => n6480, A3 => n6479, A4 => n6478
                           , ZN => n1633);
   U919 : AOI211_X1 port map( C1 => n7824, C2 => DATA1(12), A => n6483, B => 
                           n6482, ZN => n6485);
   U920 : NAND2_X1 port map( A1 => DATA1(14), A2 => n7825, ZN => n6484);
   U921 : OAI211_X1 port map( C1 => n7707, C2 => n7695, A => n6485, B => n6484,
                           ZN => n1615);
   U922 : AOI211_X1 port map( C1 => n7824, C2 => DATA1(10), A => n6487, B => 
                           n6486, ZN => n6489);
   U923 : OAI211_X1 port map( C1 => n7707, C2 => n1933, A => n6489, B => n6488,
                           ZN => n6490);
   U924 : AOI222_X1 port map( A1 => n6490, A2 => n1068, B1 => n1633, B2 => 
                           n6970, C1 => n1615, C2 => n6969, ZN => n1708);
   U925 : INV_X1 port map( A => n1934, ZN => n6491);
   U926 : AOI222_X1 port map( A1 => n6491, A2 => n1068, B1 => n6490, B2 => 
                           n6970, C1 => n1633, C2 => n6969, ZN => n1728);
   U927 : INV_X1 port map( A => n1935, ZN => n6492);
   U928 : AOI222_X1 port map( A1 => n6492, A2 => n1068, B1 => n6491, B2 => 
                           n6970, C1 => n6490, C2 => n6969, ZN => n1655);
   U929 : NAND2_X1 port map( A1 => DATA1(9), A2 => n7826, ZN => n6493);
   U930 : NAND2_X1 port map( A1 => DATA1(10), A2 => n7692, ZN => n7685);
   U931 : OAI211_X1 port map( C1 => n7688, C2 => n7175, A => n6493, B => n7685,
                           ZN => n6494);
   U932 : AOI211_X1 port map( C1 => n7824, C2 => DATA1(7), A => n6495, B => 
                           n6494, ZN => n1724);
   U933 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n1986);
   U934 : NAND2_X1 port map( A1 => DATA2_I_24_port, A2 => DATA1(24), ZN => 
                           n2082);
   U935 : NOR2_X1 port map( A1 => n2082, A2 => n6496, ZN => n6017);
   U936 : OAI21_X1 port map( B1 => n1843, B2 => n6017, A => n2058, ZN => n2031)
                           ;
   U937 : INV_X1 port map( A => n6497, ZN => n6499);
   U938 : NAND2_X1 port map( A1 => FUNC(1), A2 => n7373, ZN => n6498);
   U939 : NOR4_X1 port map( A1 => n7658, A2 => n6499, A3 => n1968, A4 => n6498,
                           ZN => n2690);
   U940 : OAI222_X1 port map( A1 => n4521, A2 => n4431, B1 => n4496, B2 => 
                           n4432, C1 => n4484, C2 => n3890, ZN => n6516);
   U941 : OAI222_X1 port map( A1 => n4521, A2 => n3890, B1 => n4483, B2 => 
                           n3883, C1 => n4482, C2 => n3889, ZN => n6570);
   U942 : OAI222_X1 port map( A1 => n4521, A2 => n4432, B1 => n4483, B2 => 
                           n3889, C1 => n3890, C2 => n4495, ZN => n6539);
   U943 : AOI22_X1 port map( A1 => n4489, A2 => n6570, B1 => n7721, B2 => n6539
                           , ZN => n6501);
   U944 : AOI22_X1 port map( A1 => n4469, A2 => n4429, B1 => n4459, B2 => n4430
                           , ZN => n6500);
   U945 : NAND2_X1 port map( A1 => n6501, A2 => n6500, ZN => n6502);
   U946 : AOI21_X1 port map( B1 => n4480, B2 => n6516, A => n6502, ZN => n6513)
                           ;
   U947 : AOI22_X1 port map( A1 => n4498, A2 => n4434, B1 => n4109, B2 => n4435
                           , ZN => n6503);
   U948 : OAI21_X1 port map( B1 => n7741, B2 => n7788, A => n6503, ZN => n6561)
                           ;
   U949 : AOI22_X1 port map( A1 => n4469, A2 => n4428, B1 => n4459, B2 => n6561
                           , ZN => n6504);
   U950 : OAI211_X1 port map( C1 => n4477, C2 => n3812, A => n3884, B => n6504,
                           ZN => n6533);
   U951 : OAI211_X1 port map( C1 => n3813, C2 => n4479, A => n3887, B => n3886,
                           ZN => n6523);
   U952 : AOI22_X1 port map( A1 => n4473, A2 => n6533, B1 => n4243, B2 => n6523
                           , ZN => n6508);
   U953 : AOI22_X1 port map( A1 => n4103, A2 => n6516, B1 => n4289, B2 => n4429
                           , ZN => n6505);
   U954 : OAI211_X1 port map( C1 => n4478, C2 => n3809, A => n3885, B => n6505,
                           ZN => n6522);
   U955 : AOI22_X1 port map( A1 => n4103, A2 => n6539, B1 => n4289, B2 => n6516
                           , ZN => n6506);
   U956 : OAI211_X1 port map( C1 => n4478, C2 => n3810, A => n3888, B => n6506,
                           ZN => n6542);
   U957 : AOI22_X1 port map( A1 => n4468, A2 => n6522, B1 => n7765, B2 => n6542
                           , ZN => n6507);
   U958 : OAI211_X1 port map( C1 => n6513, C2 => n7768, A => n6508, B => n6507,
                           ZN => n6538);
   U959 : AOI22_X1 port map( A1 => n6539, A2 => n4480, B1 => n4505, B2 => n4429
                           , ZN => n6509);
   U960 : INV_X1 port map( A => n6509, ZN => n6512);
   U961 : INV_X1 port map( A => n6570, ZN => n6519);
   U962 : OAI22_X1 port map( A1 => n4483, A2 => n3882, B1 => n4495, B2 => n3883
                           , ZN => n6510);
   U963 : AOI21_X1 port map( B1 => n7737, B2 => n7782, A => n6510, ZN => n6672)
                           ;
   U964 : OAI22_X1 port map( A1 => n4477, A2 => n6519, B1 => n6672, B2 => n7725
                           , ZN => n6511);
   U965 : AOI211_X1 port map( C1 => n4469, C2 => n6516, A => n6512, B => n6511,
                           ZN => n6543);
   U966 : AOI22_X1 port map( A1 => n4471, A2 => n6522, B1 => n4473, B2 => n6523
                           , ZN => n6515);
   U967 : INV_X1 port map( A => n6513, ZN => n6568);
   U968 : AOI22_X1 port map( A1 => n4468, A2 => n6542, B1 => n7765, B2 => n6568
                           , ZN => n6514);
   U969 : OAI211_X1 port map( C1 => n6543, C2 => n7768, A => n6515, B => n6514,
                           ZN => n6547);
   U970 : AOI22_X1 port map( A1 => n4473, A2 => n6522, B1 => n4468, B2 => n6568
                           , ZN => n6521);
   U971 : INV_X1 port map( A => n6672, ZN => n6571);
   U972 : OAI222_X1 port map( A1 => n4521, A2 => n3883, B1 => n4482, B2 => 
                           n3882, C1 => n4503, C2 => n6021, ZN => n6671);
   U973 : AOI22_X1 port map( A1 => n4289, A2 => n6571, B1 => n4489, B2 => n6671
                           , ZN => n6518);
   U974 : AOI22_X1 port map( A1 => n4505, A2 => n6516, B1 => n7764, B2 => n6539
                           , ZN => n6517);
   U975 : OAI211_X1 port map( C1 => n6519, C2 => n7763, A => n6518, B => n6517,
                           ZN => n6684);
   U976 : AOI22_X1 port map( A1 => n4471, A2 => n6542, B1 => n4475, B2 => n6684
                           , ZN => n6520);
   U977 : OAI211_X1 port map( C1 => n4244, C2 => n6543, A => n6521, B => n6520,
                           ZN => n6578);
   U978 : AOI222_X1 port map( A1 => n6538, A2 => n4256, B1 => n6547, B2 => 
                           n4456, C1 => n6578, C2 => n4455, ZN => n6565);
   U979 : INV_X1 port map( A => n6565, ZN => n6697);
   U980 : INV_X1 port map( A => n6522, ZN => n6528);
   U981 : INV_X1 port map( A => n6523, ZN => n6551);
   U982 : OAI22_X1 port map( A1 => n6528, A2 => n7755, B1 => n6551, B2 => n7719
                           , ZN => n6527);
   U983 : OAI22_X1 port map( A1 => n4477, A2 => n3811, B1 => n4520, B2 => n3813
                           , ZN => n6525);
   U984 : AOI222_X1 port map( A1 => n4517, A2 => n3891, B1 => n4498, B2 => 
                           n4433, C1 => n4485, C2 => n4434, ZN => n6582);
   U985 : OAI22_X1 port map( A1 => n4478, A2 => n3814, B1 => n4290, B2 => n6582
                           , ZN => n6524);
   U986 : AOI211_X1 port map( C1 => n4474, C2 => n6561, A => n6525, B => n6524,
                           ZN => n6585);
   U987 : INV_X1 port map( A => n6533, ZN => n6558);
   U988 : OAI22_X1 port map( A1 => n4476, A2 => n6585, B1 => n6558, B2 => n7759
                           , ZN => n6526);
   U989 : AOI211_X1 port map( C1 => n4475, C2 => n6542, A => n6527, B => n6526,
                           ZN => n6554);
   U990 : INV_X1 port map( A => n6538, ZN => n6534);
   U991 : OAI22_X1 port map( A1 => n4245, A2 => n6528, B1 => n6551, B2 => n7755
                           , ZN => n6532);
   U992 : OAI22_X1 port map( A1 => n4477, A2 => n3814, B1 => n4519, B2 => n3811
                           , ZN => n6530);
   U993 : AOI222_X1 port map( A1 => n4517, A2 => n3881, B1 => n4485, B2 => 
                           n4433, C1 => n3931, C2 => n3891, ZN => n6590);
   U994 : OAI22_X1 port map( A1 => n4290, A2 => n6590, B1 => n4102, B2 => n6582
                           , ZN => n6529);
   U995 : AOI211_X1 port map( C1 => n4480, C2 => n6561, A => n6530, B => n6529,
                           ZN => n6591);
   U996 : OAI22_X1 port map( A1 => n6585, A2 => n7766, B1 => n6591, B2 => n7734
                           , ZN => n6531);
   U997 : AOI211_X1 port map( C1 => n4468, C2 => n6533, A => n6532, B => n6531,
                           ZN => n6564);
   U998 : OAI222_X1 port map( A1 => n7730, A2 => n6554, B1 => n7720, B2 => 
                           n6534, C1 => n7758, C2 => n6564, ZN => n6535);
   U999 : INV_X1 port map( A => n6535, ZN => n6599);
   U1000 : INV_X1 port map( A => n6547, ZN => n6536);
   U1001 : OAI22_X1 port map( A1 => n7758, A2 => n6554, B1 => n7720, B2 => 
                           n6536, ZN => n6537);
   U1002 : AOI21_X1 port map( B1 => n6538, B2 => n4456, A => n6537, ZN => n6670
                           );
   U1003 : OAI22_X1 port map( A1 => n7749, A2 => n6599, B1 => n4463, B2 => 
                           n6670, ZN => n6557);
   U1004 : NAND2_X1 port map( A1 => n4522, A2 => n4540, ZN => n6839);
   U1005 : NAND4_X1 port map( A1 => n4229, A2 => n4237, A3 => n3878, A4 => 
                           n6839, ZN => n6677);
   U1006 : AOI222_X1 port map( A1 => n6677, A2 => n4485, B1 => n4497, B2 => 
                           n3879, C1 => n4516, C2 => n4427, ZN => n6572);
   U1007 : AOI22_X1 port map( A1 => n4474, A2 => n6570, B1 => n7740, B2 => 
                           n6539, ZN => n6541);
   U1008 : AOI22_X1 port map( A1 => n7735, A2 => n6571, B1 => n7721, B2 => 
                           n6671, ZN => n6540);
   U1009 : OAI211_X1 port map( C1 => n4519, C2 => n6572, A => n6541, B => n6540
                           , ZN => n6685);
   U1010 : INV_X1 port map( A => n6685, ZN => n6546);
   U1011 : AOI22_X1 port map( A1 => n7727, A2 => n6568, B1 => n7761, B2 => 
                           n6542, ZN => n6545);
   U1012 : INV_X1 port map( A => n6543, ZN => n6683);
   U1013 : AOI22_X1 port map( A1 => n7756, A2 => n6683, B1 => n6684, B2 => 
                           n4518, ZN => n6544);
   U1014 : OAI211_X1 port map( C1 => n4245, C2 => n6546, A => n6545, B => n6544
                           , ZN => n6691);
   U1015 : AOI222_X1 port map( A1 => n4456, A2 => n6578, B1 => n4455, B2 => 
                           n6691, C1 => n4256, C2 => n6547, ZN => n6669);
   U1016 : AOI22_X1 port map( A1 => n4428, A2 => n4489, B1 => n7740, B2 => 
                           n7781, ZN => n6550);
   U1017 : INV_X1 port map( A => n6582, ZN => n6548);
   U1018 : AOI22_X1 port map( A1 => n7735, A2 => n6548, B1 => n7721, B2 => 
                           n6561, ZN => n6549);
   U1019 : OAI211_X1 port map( C1 => n4102, C2 => n6590, A => n6550, B => n6549
                           , ZN => n6614);
   U1020 : OAI22_X1 port map( A1 => n4244, A2 => n6558, B1 => n6551, B2 => 
                           n7768, ZN => n6553);
   U1021 : OAI22_X1 port map( A1 => n6585, A2 => n7719, B1 => n6591, B2 => 
                           n7766, ZN => n6552);
   U1022 : AOI211_X1 port map( C1 => n4473, C2 => n6614, A => n6553, B => n6552
                           , ZN => n6595);
   U1023 : OAI222_X1 port map( A1 => n7730, A2 => n6564, B1 => n7720, B2 => 
                           n6554, C1 => n7758, C2 => n6595, ZN => n6555);
   U1024 : INV_X1 port map( A => n6555, ZN => n6626);
   U1025 : OAI22_X1 port map( A1 => n7738, A2 => n6669, B1 => n4462, B2 => 
                           n6626, ZN => n6556);
   U1026 : AOI211_X1 port map( C1 => n7796, C2 => n6697, A => n6557, B => n6556
                           , ZN => n6702);
   U1027 : OAI22_X1 port map( A1 => n4244, A2 => n6585, B1 => n6558, B2 => 
                           n7768, ZN => n6563);
   U1028 : OAI22_X1 port map( A1 => n4290, A2 => n3805, B1 => n4102, B2 => 
                           n3807, ZN => n6560);
   U1029 : OAI22_X1 port map( A1 => n4478, A2 => n6590, B1 => n4477, B2 => 
                           n6582, ZN => n6559);
   U1030 : AOI211_X1 port map( C1 => n4489, C2 => n6561, A => n6560, B => n6559
                           , ZN => n6618);
   U1031 : OAI22_X1 port map( A1 => n4476, A2 => n6618, B1 => n4101, B2 => 
                           n6591, ZN => n6562);
   U1032 : AOI211_X1 port map( C1 => n7727, C2 => n6614, A => n6563, B => n6562
                           , ZN => n6596);
   U1033 : OAI222_X1 port map( A1 => n7730, A2 => n6595, B1 => n7720, B2 => 
                           n6564, C1 => n7758, C2 => n6596, ZN => n6620);
   U1034 : OAI22_X1 port map( A1 => n4234, A2 => n6626, B1 => n4235, B2 => 
                           n6670, ZN => n6567);
   U1035 : OAI22_X1 port map( A1 => n4463, A2 => n6599, B1 => n6565, B2 => 
                           n7738, ZN => n6566);
   U1036 : AOI211_X1 port map( C1 => n7794, C2 => n6620, A => n6567, B => n6566
                           , ZN => n6698);
   U1037 : OAI22_X1 port map( A1 => n4462, A2 => n6599, B1 => n4234, B2 => 
                           n6670, ZN => n6580);
   U1038 : INV_X1 port map( A => n6684, ZN => n6577);
   U1039 : AOI22_X1 port map( A1 => n4471, A2 => n6683, B1 => n4473, B2 => 
                           n6568, ZN => n6576);
   U1040 : AOI211_X1 port map( C1 => n4522, C2 => n4542, A => n4233, B => n7791
                           , ZN => n6569);
   U1041 : NAND2_X1 port map( A1 => n4540, A2 => n4501, ZN => n6855);
   U1042 : OAI211_X1 port map( C1 => n4511, C2 => n4490, A => n6569, B => n6855
                           , ZN => n6675);
   U1043 : AOI222_X1 port map( A1 => n6675, A2 => n4485, B1 => n4516, B2 => 
                           n3879, C1 => n6677, C2 => n4497, ZN => n6679);
   U1044 : AOI22_X1 port map( A1 => n4469, A2 => n6571, B1 => n4459, B2 => 
                           n6570, ZN => n6574);
   U1045 : INV_X1 port map( A => n6572, ZN => n6682);
   U1046 : AOI22_X1 port map( A1 => n7735, A2 => n6671, B1 => n7721, B2 => 
                           n6682, ZN => n6573);
   U1047 : OAI211_X1 port map( C1 => n4519, C2 => n6679, A => n6574, B => n6573
                           , ZN => n6686);
   U1048 : AOI22_X1 port map( A1 => n4466, A2 => n6686, B1 => n7765, B2 => 
                           n6685, ZN => n6575);
   U1049 : OAI211_X1 port map( C1 => n6577, C2 => n7719, A => n6576, B => n6575
                           , ZN => n6692);
   U1050 : AOI222_X1 port map( A1 => n6578, A2 => n4256, B1 => n6691, B2 => 
                           n4456, C1 => n6692, C2 => n4455, ZN => n6694);
   U1051 : OAI22_X1 port map( A1 => n4464, A2 => n6694, B1 => n6669, B2 => 
                           n7801, ZN => n6579);
   U1052 : AOI211_X1 port map( C1 => n7723, C2 => n6697, A => n6580, B => n6579
                           , ZN => n6701);
   U1053 : OAI22_X1 port map( A1 => n4460, A2 => n6698, B1 => n4507, B2 => 
                           n6701, ZN => n6581);
   U1054 : INV_X1 port map( A => n6581, ZN => n6604);
   U1055 : OAI22_X1 port map( A1 => n4478, A2 => n3807, B1 => n4291, B2 => 
                           n3804, ZN => n6584);
   U1056 : OAI22_X1 port map( A1 => n4477, A2 => n6590, B1 => n4519, B2 => 
                           n6582, ZN => n6583);
   U1057 : AOI211_X1 port map( C1 => n4474, C2 => n6012, A => n6584, B => n6583
                           , ZN => n6639);
   U1058 : OAI22_X1 port map( A1 => n4476, A2 => n6639, B1 => n4245, B2 => 
                           n6585, ZN => n6587);
   U1059 : OAI22_X1 port map( A1 => n4472, A2 => n6618, B1 => n6591, B2 => 
                           n7755, ZN => n6586);
   U1060 : AOI211_X1 port map( C1 => n7756, C2 => n6614, A => n6587, B => n6586
                           , ZN => n6621);
   U1061 : AOI22_X1 port map( A1 => n4480, A2 => n6012, B1 => n4289, B2 => 
                           n6011, ZN => n6589);
   U1062 : OAI222_X1 port map( A1 => n4521, A2 => n3877, B1 => n4483, B2 => 
                           n4426, C1 => n4495, C2 => n4425, ZN => n6654);
   U1063 : AOI22_X1 port map( A1 => n4469, A2 => n6013, B1 => n4459, B2 => 
                           n6654, ZN => n6588);
   U1064 : OAI211_X1 port map( C1 => n4519, C2 => n6590, A => n6589, B => n6588
                           , ZN => n6613);
   U1065 : OAI22_X1 port map( A1 => n6591, A2 => n7722, B1 => n6639, B2 => 
                           n7766, ZN => n6594);
   U1066 : INV_X1 port map( A => n6614, ZN => n6592);
   U1067 : OAI22_X1 port map( A1 => n4101, A2 => n6618, B1 => n6592, B2 => 
                           n7755, ZN => n6593);
   U1068 : AOI211_X1 port map( C1 => n4473, C2 => n6613, A => n6594, B => n6593
                           , ZN => n6622);
   U1069 : OAI222_X1 port map( A1 => n7730, A2 => n6621, B1 => n7720, B2 => 
                           n6596, C1 => n7758, C2 => n6622, ZN => n6662);
   U1070 : OAI22_X1 port map( A1 => n4464, A2 => n6599, B1 => n4235, B2 => 
                           n6626, ZN => n6598);
   U1071 : INV_X1 port map( A => n6620, ZN => n6625);
   U1072 : OAI222_X1 port map( A1 => n6621, A2 => n7758, B1 => n6596, B2 => 
                           n7730, C1 => n6595, C2 => n7720, ZN => n6643);
   U1073 : INV_X1 port map( A => n6643, ZN => n6627);
   U1074 : OAI22_X1 port map( A1 => n4463, A2 => n6625, B1 => n6627, B2 => 
                           n7749, ZN => n6597);
   U1075 : AOI211_X1 port map( C1 => n7794, C2 => n6662, A => n6598, B => n6597
                           , ZN => n6649);
   U1076 : OAI22_X1 port map( A1 => n4463, A2 => n6626, B1 => n6599, B2 => 
                           n7801, ZN => n6601);
   U1077 : OAI22_X1 port map( A1 => n4464, A2 => n6670, B1 => n4234, B2 => 
                           n6625, ZN => n6600);
   U1078 : AOI211_X1 port map( C1 => n7794, C2 => n6643, A => n6601, B => n6600
                           , ZN => n6699);
   U1079 : OAI22_X1 port map( A1 => n4250, A2 => n6649, B1 => n4094, B2 => 
                           n6699, ZN => n6602);
   U1080 : INV_X1 port map( A => n6602, ZN => n6603);
   U1081 : OAI211_X1 port map( C1 => n7805, C2 => n6702, A => n6604, B => n6603
                           , ZN => n6709);
   U1082 : INV_X1 port map( A => n6639, ZN => n6612);
   U1083 : AOI22_X1 port map( A1 => n4480, A2 => n6013, B1 => n4289, B2 => 
                           n6012, ZN => n6606);
   U1084 : OAI222_X1 port map( A1 => n4521, A2 => n3917, B1 => n4483, B2 => 
                           n4425, C1 => n4495, C2 => n3877, ZN => n6653);
   U1085 : AOI22_X1 port map( A1 => n4469, A2 => n6654, B1 => n4459, B2 => 
                           n6653, ZN => n6605);
   U1086 : OAI211_X1 port map( C1 => n4519, C2 => n3807, A => n6606, B => n6605
                           , ZN => n6615);
   U1087 : INV_X1 port map( A => n6615, ZN => n6710);
   U1088 : OAI22_X1 port map( A1 => n7759, A2 => n6710, B1 => n4245, B2 => 
                           n6618, ZN => n6611);
   U1089 : INV_X1 port map( A => n6653, ZN => n6712);
   U1090 : AOI22_X1 port map( A1 => n6013, A2 => n4289, B1 => n7760, B2 => 
                           n7792, ZN => n6608);
   U1091 : OAI222_X1 port map( A1 => n4521, A2 => n3916, B1 => n4483, B2 => 
                           n3877, C1 => n4495, C2 => n3917, ZN => n6711);
   U1092 : AOI22_X1 port map( A1 => n3927, A2 => n6654, B1 => n4459, B2 => 
                           n6711, ZN => n6607);
   U1093 : OAI211_X1 port map( C1 => n6712, C2 => n7767, A => n6608, B => n6607
                           , ZN => n6609);
   U1094 : INV_X1 port map( A => n6609, ZN => n6757);
   U1095 : INV_X1 port map( A => n6613, ZN => n6652);
   U1096 : OAI22_X1 port map( A1 => n7734, A2 => n6757, B1 => n7719, B2 => 
                           n6652, ZN => n6610);
   U1097 : AOI211_X1 port map( C1 => n6612, C2 => n4518, A => n6611, B => n6610
                           , ZN => n6660);
   U1098 : AOI22_X1 port map( A1 => n4471, A2 => n6613, B1 => n7756, B2 => 
                           n6612, ZN => n6617);
   U1099 : AOI22_X1 port map( A1 => n7761, A2 => n6615, B1 => n7739, B2 => 
                           n6614, ZN => n6616);
   U1100 : OAI211_X1 port map( C1 => n4244, C2 => n6618, A => n6617, B => n6616
                           , ZN => n6619);
   U1101 : INV_X1 port map( A => n6619, ZN => n6642);
   U1102 : OAI222_X1 port map( A1 => n6660, A2 => n7758, B1 => n6642, B2 => 
                           n7730, C1 => n6622, C2 => n7720, ZN => n6661);
   U1103 : INV_X1 port map( A => n6661, ZN => n6768);
   U1104 : AOI22_X1 port map( A1 => n7736, A2 => n6620, B1 => n7796, B2 => 
                           n6643, ZN => n6624);
   U1105 : OAI222_X1 port map( A1 => n7730, A2 => n6622, B1 => n7720, B2 => 
                           n6621, C1 => n7758, C2 => n6642, ZN => n6722);
   U1106 : AOI22_X1 port map( A1 => n4453, A2 => n6722, B1 => n7723, B2 => 
                           n6662, ZN => n6623);
   U1107 : OAI211_X1 port map( C1 => n4462, C2 => n6768, A => n6624, B => n6623
                           , ZN => n6755);
   U1108 : OAI22_X1 port map( A1 => n4464, A2 => n6626, B1 => n4235, B2 => 
                           n6625, ZN => n6629);
   U1109 : INV_X1 port map( A => n6662, ZN => n6646);
   U1110 : OAI22_X1 port map( A1 => n4463, A2 => n6627, B1 => n6646, B2 => 
                           n7749, ZN => n6628);
   U1111 : AOI211_X1 port map( C1 => n7794, C2 => n6722, A => n6629, B => n6628
                           , ZN => n6650);
   U1112 : OAI22_X1 port map( A1 => n4094, A2 => n6650, B1 => n6699, B2 => 
                           n7805, ZN => n6631);
   U1113 : OAI22_X1 port map( A1 => n4460, A2 => n6649, B1 => n4507, B2 => 
                           n6698, ZN => n6630);
   U1114 : AOI211_X1 port map( C1 => n7750, C2 => n6755, A => n6631, B => n6630
                           , ZN => n6632);
   U1115 : INV_X1 port map( A => n6632, ZN => n6668);
   U1116 : INV_X1 port map( A => n6649, ZN => n6651);
   U1117 : OAI22_X1 port map( A1 => n4098, A2 => n6698, B1 => n6699, B2 => 
                           n7799, ZN => n6634);
   U1118 : OAI22_X1 port map( A1 => n6702, A2 => n7751, B1 => n6650, B2 => 
                           n7808, ZN => n6633);
   U1119 : AOI211_X1 port map( C1 => n4436, C2 => n6651, A => n6634, B => n6633
                           , ZN => n6635);
   U1120 : INV_X1 port map( A => n6635, ZN => n6707);
   U1121 : AOI222_X1 port map( A1 => n7728, A2 => n6709, B1 => n7797, B2 => 
                           n6668, C1 => n7747, C2 => n6707, ZN => n6781);
   U1122 : INV_X1 port map( A => n6781, ZN => n6732);
   U1123 : OAI22_X1 port map( A1 => n4460, A2 => n6650, B1 => n4507, B2 => 
                           n6699, ZN => n6636);
   U1124 : INV_X1 port map( A => n6636, ZN => n6648);
   U1125 : AOI22_X1 port map( A1 => n4103, A2 => n6013, B1 => n4289, B2 => 
                           n6654, ZN => n6638);
   U1126 : AOI22_X1 port map( A1 => n4469, A2 => n6711, B1 => n4459, B2 => 
                           n6718, ZN => n6637);
   U1127 : OAI211_X1 port map( C1 => n4478, C2 => n6712, A => n6638, B => n6637
                           , ZN => n7097);
   U1128 : OAI22_X1 port map( A1 => n4472, A2 => n6757, B1 => n6652, B2 => 
                           n7755, ZN => n6641);
   U1129 : OAI22_X1 port map( A1 => n6639, A2 => n7722, B1 => n6710, B2 => 
                           n7719, ZN => n6640);
   U1130 : AOI211_X1 port map( C1 => n4473, C2 => n7097, A => n6641, B => n6640
                           , ZN => n6721);
   U1131 : OAI222_X1 port map( A1 => n7730, A2 => n6660, B1 => n7720, B2 => 
                           n6642, C1 => n7758, C2 => n6721, ZN => n7004);
   U1132 : AOI22_X1 port map( A1 => n7794, A2 => n7004, B1 => n7723, B2 => 
                           n6722, ZN => n6645);
   U1133 : AOI22_X1 port map( A1 => n4112, A2 => n6643, B1 => n7733, B2 => 
                           n6661, ZN => n6644);
   U1134 : OAI211_X1 port map( C1 => n4235, C2 => n6646, A => n6645, B => n6644
                           , ZN => n6776);
   U1135 : AOI22_X1 port map( A1 => n4436, A2 => n6755, B1 => n7750, B2 => 
                           n6776, ZN => n6647);
   U1136 : OAI211_X1 port map( C1 => n4098, C2 => n6649, A => n6648, B => n6647
                           , ZN => n6728);
   U1137 : AOI222_X1 port map( A1 => n7747, A2 => n6668, B1 => n6707, B2 => 
                           n7728, C1 => n6728, C2 => n7797, ZN => n6750);
   U1138 : INV_X1 port map( A => n6776, ZN => n6923);
   U1139 : INV_X1 port map( A => n6650, ZN => n6725);
   U1140 : AOI22_X1 port map( A1 => n4110, A2 => n6651, B1 => n4439, B2 => 
                           n6725, ZN => n6667);
   U1141 : INV_X1 port map( A => n6722, ZN => n6665);
   U1142 : OAI22_X1 port map( A1 => n6652, A2 => n7722, B1 => n6757, B2 => 
                           n7719, ZN => n6659);
   U1143 : AOI22_X1 port map( A1 => n4459, A2 => n6714, B1 => n7721, B2 => 
                           n6653, ZN => n6656);
   U1144 : AOI22_X1 port map( A1 => n4103, A2 => n6654, B1 => n3927, B2 => 
                           n6711, ZN => n6655);
   U1145 : NAND2_X1 port map( A1 => n6656, A2 => n6655, ZN => n6657);
   U1146 : AOI21_X1 port map( B1 => n4469, B2 => n6718, A => n6657, ZN => n7114
                           );
   U1147 : OAI22_X1 port map( A1 => n4244, A2 => n6710, B1 => n7114, B2 => 
                           n7734, ZN => n6658);
   U1148 : AOI211_X1 port map( C1 => n4243, C2 => n7097, A => n6659, B => n6658
                           , ZN => n6767);
   U1149 : OAI222_X1 port map( A1 => n7730, A2 => n6721, B1 => n7720, B2 => 
                           n6660, C1 => n7758, C2 => n6767, ZN => n7021);
   U1150 : AOI22_X1 port map( A1 => n7794, A2 => n7021, B1 => n7723, B2 => 
                           n6661, ZN => n6664);
   U1151 : AOI22_X1 port map( A1 => n4112, A2 => n6662, B1 => n7733, B2 => 
                           n7004, ZN => n6663);
   U1152 : OAI211_X1 port map( C1 => n4235, C2 => n6665, A => n6664, B => n6663
                           , ZN => n6773);
   U1153 : AOI22_X1 port map( A1 => n3921, A2 => n6755, B1 => n4461, B2 => 
                           n6773, ZN => n6666);
   U1154 : OAI211_X1 port map( C1 => n4094, C2 => n6923, A => n6667, B => n6666
                           , ZN => n6753);
   U1155 : AOI222_X1 port map( A1 => n7747, A2 => n6728, B1 => n6668, B2 => 
                           n7728, C1 => n6753, C2 => n7797, ZN => n6751);
   U1156 : OAI22_X1 port map( A1 => n6750, A2 => n7753, B1 => n6751, B2 => 
                           n4091, ZN => n6731);
   U1157 : OAI22_X1 port map( A1 => n4462, A2 => n6670, B1 => n6669, B2 => 
                           n7802, ZN => n6696);
   U1158 : INV_X1 port map( A => n6671, ZN => n6673);
   U1159 : OAI22_X1 port map( A1 => n4102, A2 => n6673, B1 => n6672, B2 => 
                           n7772, ZN => n6681);
   U1160 : NAND2_X1 port map( A1 => n4502, A2 => n7742, ZN => n6840);
   U1161 : NAND2_X1 port map( A1 => n4522, A2 => n7726, ZN => n6742);
   U1162 : NAND4_X1 port map( A1 => n3876, A2 => n6674, A3 => n6840, A4 => 
                           n6742, ZN => n6676);
   U1163 : AOI222_X1 port map( A1 => n6677, A2 => n4516, B1 => n6676, B2 => 
                           n4485, C1 => n6675, C2 => n4497, ZN => n6678);
   U1164 : OAI22_X1 port map( A1 => n4477, A2 => n6679, B1 => n4519, B2 => 
                           n6678, ZN => n6680);
   U1165 : AOI211_X1 port map( C1 => n7735, C2 => n6682, A => n6681, B => n6680
                           , ZN => n6689);
   U1166 : AOI22_X1 port map( A1 => n4471, A2 => n6684, B1 => n4473, B2 => 
                           n6683, ZN => n6688);
   U1167 : AOI22_X1 port map( A1 => n4518, A2 => n6686, B1 => n7756, B2 => 
                           n6685, ZN => n6687);
   U1168 : OAI211_X1 port map( C1 => n4245, C2 => n6689, A => n6688, B => n6687
                           , ZN => n6690);
   U1169 : AOI222_X1 port map( A1 => n7724, A2 => n6692, B1 => n6691, B2 => 
                           n7731, C1 => n6690, C2 => n7757, ZN => n6693);
   U1170 : OAI22_X1 port map( A1 => n4235, A2 => n6694, B1 => n6693, B2 => 
                           n7738, ZN => n6695);
   U1171 : AOI211_X1 port map( C1 => n7733, C2 => n6697, A => n6696, B => n6695
                           , ZN => n6706);
   U1172 : OAI22_X1 port map( A1 => n4250, A2 => n6699, B1 => n4094, B2 => 
                           n6698, ZN => n6700);
   U1173 : INV_X1 port map( A => n6700, ZN => n6705);
   U1174 : OAI22_X1 port map( A1 => n7799, A2 => n6702, B1 => n4098, B2 => 
                           n6701, ZN => n6703);
   U1175 : INV_X1 port map( A => n6703, ZN => n6704);
   U1176 : OAI211_X1 port map( C1 => n6706, C2 => n7751, A => n6705, B => n6704
                           , ZN => n6708);
   U1177 : AOI222_X1 port map( A1 => n6709, A2 => n4219, B1 => n6708, B2 => 
                           n4444, C1 => n6707, C2 => n3906, ZN => n6729);
   U1178 : OAI22_X1 port map( A1 => n6710, A2 => n7722, B1 => n6757, B2 => 
                           n7755, ZN => n6720);
   U1179 : INV_X1 port map( A => n6711, ZN => n6759);
   U1180 : OAI22_X1 port map( A1 => n4519, A2 => n6712, B1 => n6759, B2 => 
                           n7732, ZN => n6717);
   U1181 : AOI22_X1 port map( A1 => n6714, A2 => n4469, B1 => n6713, B2 => 
                           n4505, ZN => n6715);
   U1182 : INV_X1 port map( A => n6715, ZN => n6716);
   U1183 : AOI211_X1 port map( C1 => n3927, C2 => n6718, A => n6717, B => n6716
                           , ZN => n7134);
   U1184 : OAI22_X1 port map( A1 => n4472, A2 => n7114, B1 => n7134, B2 => 
                           n7734, ZN => n6719);
   U1185 : AOI211_X1 port map( C1 => n4468, C2 => n7097, A => n6720, B => n6719
                           , ZN => n7067);
   U1186 : OAI222_X1 port map( A1 => n7730, A2 => n6767, B1 => n7720, B2 => 
                           n6721, C1 => n7758, C2 => n7067, ZN => n7036);
   U1187 : AOI22_X1 port map( A1 => n7794, A2 => n7036, B1 => n7733, B2 => 
                           n7021, ZN => n6724);
   U1188 : AOI22_X1 port map( A1 => n4112, A2 => n6722, B1 => n7723, B2 => 
                           n7004, ZN => n6723);
   U1189 : OAI211_X1 port map( C1 => n4235, C2 => n6768, A => n6724, B => n6723
                           , ZN => n6754);
   U1190 : AOI22_X1 port map( A1 => n7750, A2 => n6754, B1 => n7804, B2 => 
                           n6725, ZN => n6727);
   U1191 : AOI22_X1 port map( A1 => n4436, A2 => n6773, B1 => n7800, B2 => 
                           n6755, ZN => n6726);
   U1192 : OAI211_X1 port map( C1 => n4460, C2 => n6923, A => n6727, B => n6726
                           , ZN => n6777);
   U1193 : AOI222_X1 port map( A1 => n7747, A2 => n6753, B1 => n6728, B2 => 
                           n7728, C1 => n6777, C2 => n7797, ZN => n6752);
   U1194 : OAI22_X1 port map( A1 => n4441, A2 => n6729, B1 => n6752, B2 => 
                           n7813, ZN => n6730);
   U1195 : AOI211_X1 port map( C1 => n4218, C2 => n6732, A => n6731, B => n6730
                           , ZN => n6784);
   U1196 : XNOR2_X1 port map( A => n4293, B => n7726, ZN => n6749);
   U1197 : AOI21_X1 port map( B1 => n4211, B2 => n4084, A => n4083, ZN => n6869
                           );
   U1198 : XNOR2_X1 port map( A => n4394, B => n4458, ZN => n6860);
   U1199 : OAI21_X1 port map( B1 => n4421, B2 => n6869, A => n6860, ZN => n6859
                           );
   U1200 : NAND2_X1 port map( A1 => n4395, A2 => n7762, ZN => n6736);
   U1201 : OAI21_X1 port map( B1 => n4395, B2 => n7762, A => n6736, ZN => n6850
                           );
   U1202 : AOI21_X1 port map( B1 => n4212, B2 => n6859, A => n6850, ZN => n6785
                           );
   U1203 : XOR2_X1 port map( A => n6022, B => n4397, Z => n6738);
   U1204 : INV_X1 port map( A => n6738, ZN => n6799);
   U1205 : NAND2_X1 port map( A1 => n4542, A2 => n4396, ZN => n6740);
   U1206 : OAI21_X1 port map( B1 => n6738, B2 => n6736, A => n6740, ZN => n6733
                           );
   U1207 : AOI21_X1 port map( B1 => n6785, B2 => n6799, A => n6733, ZN => n6735
                           );
   U1208 : AOI21_X1 port map( B1 => n4211, B2 => n7810, A => n4082, ZN => n6870
                           );
   U1209 : OAI21_X1 port map( B1 => n6870, B2 => n4421, A => n6860, ZN => n6858
                           );
   U1210 : AOI21_X1 port map( B1 => n4212, B2 => n6858, A => n6850, ZN => n6786
                           );
   U1211 : AOI21_X1 port map( B1 => n6786, B2 => n6799, A => n6733, ZN => n6734
                           );
   U1212 : OAI22_X1 port map( A1 => n4213, A2 => n6735, B1 => n4418, B2 => 
                           n6734, ZN => n6748);
   U1213 : INV_X1 port map( A => n6736, ZN => n6796);
   U1214 : OAI22_X1 port map( A1 => n7807, A2 => n6786, B1 => n7754, B2 => 
                           n6785, ZN => n6737);
   U1215 : INV_X1 port map( A => n6737, ZN => n6843);
   U1216 : OAI21_X1 port map( B1 => n4206, B2 => n4417, A => n6738, ZN => n6739
                           );
   U1217 : OAI21_X1 port map( B1 => n6796, B2 => n6843, A => n6739, ZN => n6795
                           );
   U1218 : NAND2_X1 port map( A1 => n6795, A2 => n6740, ZN => n6746);
   U1219 : OAI221_X1 port map( B1 => n5995, B2 => n4223, C1 => n7726, C2 => 
                           n4254, A => n4224, ZN => n6744);
   U1220 : NOR2_X1 port map( A1 => n5995, A2 => n4530, ZN => n7341);
   U1221 : AOI22_X1 port map( A1 => n7341, A2 => n4509, B1 => n4510, B2 => 
                           n3934, ZN => n6741);
   U1222 : OAI21_X1 port map( B1 => n4251, B2 => n6742, A => n6741, ZN => n6743
                           );
   U1223 : AOI21_X1 port map( B1 => n4530, B2 => n6744, A => n6743, ZN => n6745
                           );
   U1224 : OAI21_X1 port map( B1 => n6746, B2 => n6749, A => n6745, ZN => n6747
                           );
   U1225 : AOI21_X1 port map( B1 => n6749, B2 => n6748, A => n6747, ZN => n6783
                           );
   U1226 : INV_X1 port map( A => n6750, ZN => n6844);
   U1227 : INV_X1 port map( A => n6751, ZN => n6854);
   U1228 : AOI22_X1 port map( A1 => n4218, A2 => n6844, B1 => n4424, B2 => 
                           n6854, ZN => n6780);
   U1229 : INV_X1 port map( A => n6752, ZN => n6868);
   U1230 : INV_X1 port map( A => n6753, ZN => n6778);
   U1231 : INV_X1 port map( A => n6754, ZN => n6948);
   U1232 : INV_X1 port map( A => n6755, ZN => n6756);
   U1233 : OAI22_X1 port map( A1 => n4094, A2 => n6948, B1 => n6756, B2 => 
                           n7751, ZN => n6775);
   U1234 : OAI22_X1 port map( A1 => n4245, A2 => n6757, B1 => n7114, B2 => 
                           n7719, ZN => n6766);
   U1235 : OAI22_X1 port map( A1 => n6759, A2 => n7725, B1 => n6758, B2 => 
                           n7763, ZN => n6763);
   U1236 : OAI22_X1 port map( A1 => n4477, A2 => n6761, B1 => n6760, B2 => 
                           n7767, ZN => n6762);
   U1237 : AOI211_X1 port map( C1 => n4505, C2 => n6764, A => n6763, B => n6762
                           , ZN => n7152);
   U1238 : OAI22_X1 port map( A1 => n7134, A2 => n7759, B1 => n7152, B2 => 
                           n7734, ZN => n6765);
   U1239 : AOI211_X1 port map( C1 => n4518, C2 => n7097, A => n6766, B => n6765
                           , ZN => n7083);
   U1240 : OAI222_X1 port map( A1 => n7730, A2 => n7067, B1 => n7720, B2 => 
                           n6767, C1 => n7758, C2 => n7083, ZN => n7044);
   U1241 : INV_X1 port map( A => n7021, ZN => n6769);
   U1242 : OAI22_X1 port map( A1 => n4463, A2 => n6769, B1 => n6768, B2 => 
                           n7738, ZN => n6772);
   U1243 : AOI22_X1 port map( A1 => n7733, A2 => n7036, B1 => n7796, B2 => 
                           n7004, ZN => n6770);
   U1244 : INV_X1 port map( A => n6770, ZN => n6771);
   U1245 : AOI211_X1 port map( C1 => n7794, C2 => n7044, A => n6772, B => n6771
                           , ZN => n6955);
   U1246 : INV_X1 port map( A => n6773, ZN => n6934);
   U1247 : OAI22_X1 port map( A1 => n4250, A2 => n6955, B1 => n4460, B2 => 
                           n6934, ZN => n6774);
   U1248 : AOI211_X1 port map( C1 => n7800, C2 => n6776, A => n6775, B => n6774
                           , ZN => n6903);
   U1249 : INV_X1 port map( A => n6777, ZN => n6894);
   U1250 : OAI222_X1 port map( A1 => n4113, A2 => n6778, B1 => n4445, B2 => 
                           n6903, C1 => n4443, C2 => n6894, ZN => n6890);
   U1251 : AOI22_X1 port map( A1 => n4416, A2 => n6868, B1 => n4252, B2 => 
                           n6890, ZN => n6779);
   U1252 : OAI211_X1 port map( C1 => n4441, C2 => n6781, A => n6780, B => n6779
                           , ZN => n6794);
   U1253 : NAND3_X1 port map( A1 => n4513, A2 => n4205, A3 => n6794, ZN => 
                           n6782);
   U1254 : OAI211_X1 port map( C1 => n4222, C2 => n6784, A => n6783, B => n6782
                           , ZN => OUTALU(31));
   U1255 : AOI22_X1 port map( A1 => n4206, A2 => n6786, B1 => n4417, B2 => 
                           n6785, ZN => n6800);
   U1256 : NAND2_X1 port map( A1 => n4542, A2 => n4415, ZN => n6788);
   U1257 : NAND2_X1 port map( A1 => n6022, A2 => n4529, ZN => n6787);
   U1258 : NAND2_X1 port map( A1 => n6788, A2 => n6787, ZN => n7323);
   U1259 : INV_X1 port map( A => n7323, ZN => n7338);
   U1260 : AOI22_X1 port map( A1 => n3935, A2 => n4437, B1 => n4450, B2 => 
                           n7815, ZN => n6792);
   U1261 : NOR2_X1 port map( A1 => n5995, A2 => n4106, ZN => n6790);
   U1262 : OAI22_X1 port map( A1 => n4415, A2 => n7817, B1 => n4255, B2 => 
                           n7748, ZN => n6789);
   U1263 : AOI22_X1 port map( A1 => n6790, A2 => n4508, B1 => n7742, B2 => 
                           n6789, ZN => n6791);
   U1264 : OAI211_X1 port map( C1 => n7338, C2 => n4254, A => n6792, B => n6791
                           , ZN => n6793);
   U1265 : AOI21_X1 port map( B1 => n4447, B2 => n6794, A => n6793, ZN => n6798
                           );
   U1266 : OAI21_X1 port map( B1 => n6796, B2 => n6799, A => n6795, ZN => n6797
                           );
   U1267 : OAI211_X1 port map( C1 => n6800, C2 => n6799, A => n6798, B => n6797
                           , ZN => OUTALU(30));
   U1268 : NOR2_X1 port map( A1 => n7227, A2 => n7707, ZN => n6802);
   U1269 : NOR2_X1 port map( A1 => n1939, A2 => n7696, ZN => n7679);
   U1270 : AOI211_X1 port map( C1 => n7691, C2 => DATA1(0), A => n6802, B => 
                           n7679, ZN => n1979);
   U1271 : OAI22_X1 port map( A1 => n6809, A2 => n1896, B1 => n6807, B2 => 
                           n7162, ZN => n6801);
   U1272 : AOI22_X1 port map( A1 => n4257, A2 => n7823, B1 => n6810, B2 => 
                           n6801, ZN => n1978);
   U1273 : OAI21_X1 port map( B1 => n7158, B2 => n7227, A => n7143, ZN => n1976
                           );
   U1274 : AOI211_X1 port map( C1 => DATA1(6), C2 => n7709, A => n6803, B => 
                           n6802, ZN => n6805);
   U1275 : OAI211_X1 port map( C1 => n7711, C2 => n6806, A => n6805, B => n6804
                           , ZN => n2433);
   U1276 : AOI222_X1 port map( A1 => n1936, A2 => n1068, B1 => n6971, B2 => 
                           n6970, C1 => n2433, C2 => n6969, ZN => n2441);
   U1277 : AOI22_X1 port map( A1 => DATA1(2), A2 => DATA2(2), B1 => n1970, B2 
                           => n7227, ZN => n7222);
   U1278 : INV_X1 port map( A => n7222, ZN => n7177);
   U1279 : AOI22_X1 port map( A1 => n7166, A2 => n6809, B1 => n6808, B2 => 
                           n6807, ZN => n6811);
   U1280 : OAI22_X1 port map( A1 => n7177, A2 => n7161, B1 => n6811, B2 => 
                           n6810, ZN => n1974);
   U1281 : AOI211_X1 port map( C1 => n4524, C2 => n4079, A => n3872, B => n7820
                           , ZN => n6837);
   U1282 : OAI22_X1 port map( A1 => n6813, A2 => n7753, B1 => n6812, B2 => 
                           n7814, ZN => n6835);
   U1283 : AOI22_X1 port map( A1 => n4436, A2 => n6975, B1 => n6814, B2 => 
                           n7750, ZN => n6831);
   U1284 : INV_X1 port map( A => n7287, ZN => n6823);
   U1285 : OAI22_X1 port map( A1 => n4477, A2 => n3815, B1 => n4519, B2 => 
                           n3802, ZN => n6817);
   U1286 : OAI22_X1 port map( A1 => n4478, A2 => n6976, B1 => n4290, B2 => 
                           n6815, ZN => n6816);
   U1287 : AOI211_X1 port map( C1 => n4474, C2 => n6818, A => n6817, B => n6816
                           , ZN => n7284);
   U1288 : INV_X1 port map( A => n7290, ZN => n6819);
   U1289 : OAI22_X1 port map( A1 => n4245, A2 => n7284, B1 => n6819, B2 => 
                           n4101, ZN => n6822);
   U1290 : OAI22_X1 port map( A1 => n4472, A2 => n6980, B1 => n4476, B2 => 
                           n6820, ZN => n6821);
   U1291 : AOI211_X1 port map( C1 => n4518, C2 => n6823, A => n6822, B => n6821
                           , ZN => n7293);
   U1292 : OAI222_X1 port map( A1 => n4512, A2 => n6824, B1 => n4506, B2 => 
                           n7293, C1 => n4248, C2 => n6983, ZN => n7294);
   U1293 : OAI22_X1 port map( A1 => n6988, A2 => n7802, B1 => n6825, B2 => 
                           n4462, ZN => n6828);
   U1294 : OAI22_X1 port map( A1 => n7300, A2 => n7801, B1 => n6826, B2 => 
                           n7749, ZN => n6827);
   U1295 : AOI211_X1 port map( C1 => n4112, C2 => n7294, A => n6828, B => n6827
                           , ZN => n7305);
   U1296 : INV_X1 port map( A => n7305, ZN => n6829);
   U1297 : AOI22_X1 port map( A1 => n4110, A2 => n6829, B1 => n4439, B2 => 
                           n7279, ZN => n6830);
   U1298 : OAI211_X1 port map( C1 => n6832, C2 => n7799, A => n6831, B => n6830
                           , ZN => n7306);
   U1299 : AOI222_X1 port map( A1 => n7728, A2 => n7306, B1 => n7797, B2 => 
                           n6833, C1 => n6991, C2 => n7747, ZN => n7309);
   U1300 : OAI22_X1 port map( A1 => n7309, A2 => n7729, B1 => n7312, B2 => 
                           n7806, ZN => n6834);
   U1301 : OAI21_X1 port map( B1 => n6835, B2 => n6834, A => n7795, ZN => n6836
                           );
   U1302 : OAI211_X1 port map( C1 => n4222, C2 => n3875, A => n6837, B => n6836
                           , ZN => OUTALU(2));
   U1303 : AOI22_X1 port map( A1 => n6016, A2 => n4528, B1 => n4540, B2 => 
                           n4414, ZN => n7327);
   U1304 : INV_X1 port map( A => n7327, ZN => n6838);
   U1305 : AOI22_X1 port map( A1 => n3936, A2 => n4437, B1 => n4509, B2 => 
                           n6838, ZN => n6853);
   U1306 : OAI21_X1 port map( B1 => n6016, B2 => n4223, A => n4224, ZN => n6842
                           );
   U1307 : OAI211_X1 port map( C1 => n5995, C2 => n4107, A => n6840, B => n6839
                           , ZN => n6841);
   U1308 : AOI22_X1 port map( A1 => n4528, A2 => n6842, B1 => n4508, B2 => 
                           n6841, ZN => n6852);
   U1309 : OAI22_X1 port map( A1 => n7807, A2 => n6858, B1 => n7754, B2 => 
                           n6859, ZN => n6849);
   U1310 : AOI21_X1 port map( B1 => n4212, B2 => n6850, A => n6843, ZN => n6848
                           );
   U1311 : AOI22_X1 port map( A1 => n4218, A2 => n6854, B1 => n4092, B2 => 
                           n6844, ZN => n6846);
   U1312 : AOI22_X1 port map( A1 => n4416, A2 => n6890, B1 => n4424, B2 => 
                           n6868, ZN => n6845);
   U1313 : AOI21_X1 port map( B1 => n6846, B2 => n6845, A => n4222, ZN => n6847
                           );
   U1314 : AOI211_X1 port map( C1 => n6850, C2 => n6849, A => n6848, B => n6847
                           , ZN => n6851);
   U1315 : NAND3_X1 port map( A1 => n6853, A2 => n6852, A3 => n6851, ZN => 
                           OUTALU(29));
   U1316 : AOI22_X1 port map( A1 => DATA1(28), A2 => n1944, B1 => DATA2(28), B2
                           => n1906, ZN => n2670);
   U1317 : NAND3_X1 port map( A1 => DATA1(28), A2 => DATA2(28), A3 => n7105, ZN
                           => n2011);
   U1318 : AOI222_X1 port map( A1 => n6868, A2 => n4218, B1 => n6854, B2 => 
                           n4092, C1 => n6890, C2 => n4424, ZN => n6867);
   U1319 : OAI211_X1 port map( C1 => n6022, C2 => n7818, A => n4215, B => n6855
                           , ZN => n6856);
   U1320 : OAI221_X1 port map( B1 => n6856, B2 => n4500, C1 => n6856, C2 => 
                           n7726, A => n4508, ZN => n6857);
   U1321 : OAI211_X1 port map( C1 => n3871, C2 => n4254, A => n3870, B => n6857
                           , ZN => n6865);
   U1322 : AOI22_X1 port map( A1 => n4417, A2 => n6859, B1 => n6858, B2 => 
                           n7752, ZN => n6863);
   U1323 : NOR2_X1 port map( A1 => n4421, A2 => n6860, ZN => n6862);
   U1324 : AOI22_X1 port map( A1 => n6870, A2 => n7752, B1 => n4417, B2 => 
                           n6869, ZN => n6861);
   U1325 : OAI22_X1 port map( A1 => n6863, A2 => n6862, B1 => n6861, B2 => 
                           n6860, ZN => n6864);
   U1326 : AOI211_X1 port map( C1 => n4437, C2 => n3937, A => n6865, B => n6864
                           , ZN => n6866);
   U1327 : OAI21_X1 port map( B1 => n4222, B2 => n6867, A => n6866, ZN => 
                           OUTALU(28));
   U1328 : INV_X1 port map( A => DATA2(27), ZN => n7351);
   U1329 : OAI21_X1 port map( B1 => n7158, B2 => n7351, A => n7143, ZN => n2028
                           );
   U1330 : NAND2_X1 port map( A1 => DATA1(27), A2 => n7351, ZN => n2594);
   U1331 : NAND2_X1 port map( A1 => DATA2(27), A2 => n1907, ZN => n2669);
   U1332 : AOI21_X1 port map( B1 => n2669, B2 => n2594, A => n7161, ZN => n2026
                           );
   U1333 : AOI22_X1 port map( A1 => n4218, A2 => n6890, B1 => n4092, B2 => 
                           n6868, ZN => n6879);
   U1334 : NOR2_X1 port map( A1 => n6869, A2 => n4213, ZN => n6875);
   U1335 : NOR3_X1 port map( A1 => n4503, A2 => n6881, A3 => n4251, ZN => n6874
                           );
   U1336 : NOR2_X1 port map( A1 => n6870, A2 => n4418, ZN => n6876);
   U1337 : AOI22_X1 port map( A1 => n5993, A2 => n6876, B1 => n4078, B2 => 
                           n4538, ZN => n6872);
   U1338 : AOI21_X1 port map( B1 => n3938, B2 => n4437, A => n4077, ZN => n6871
                           );
   U1339 : NAND2_X1 port map( A1 => n6872, A2 => n6871, ZN => n6873);
   U1340 : AOI211_X1 port map( C1 => n4412, C2 => n6875, A => n6874, B => n6873
                           , ZN => n6878);
   U1341 : OAI22_X1 port map( A1 => n6876, A2 => n6875, B1 => n4411, B2 => 
                           n4410, ZN => n6877);
   U1342 : OAI211_X1 port map( C1 => n6879, C2 => n7803, A => n6878, B => n6877
                           , ZN => OUTALU(27));
   U1343 : NAND3_X1 port map( A1 => DATA2(26), A2 => DATA1(26), A3 => n7105, ZN
                           => n2052);
   U1344 : OAI22_X1 port map( A1 => n4482, A2 => n6881, B1 => n4503, B2 => 
                           n6880, ZN => n6882);
   U1345 : INV_X1 port map( A => n6882, ZN => n6893);
   U1346 : NOR2_X1 port map( A1 => n4213, A2 => n4412, ZN => n6885);
   U1347 : NAND2_X1 port map( A1 => n4208, A2 => n6885, ZN => n6883);
   U1348 : OAI211_X1 port map( C1 => n4254, C2 => n3869, A => n3868, B => n6883
                           , ZN => n6889);
   U1349 : NAND2_X1 port map( A1 => n7810, A2 => n7752, ZN => n6887);
   U1350 : INV_X1 port map( A => n6887, ZN => n6884);
   U1351 : OAI22_X1 port map( A1 => n6885, A2 => n6884, B1 => n4420, B2 => 
                           n4207, ZN => n6886);
   U1352 : OAI21_X1 port map( B1 => n4081, B2 => n6887, A => n6886, ZN => n6888
                           );
   U1353 : AOI211_X1 port map( C1 => n4437, C2 => n3941, A => n6889, B => n6888
                           , ZN => n6892);
   U1354 : NAND3_X1 port map( A1 => n4092, A2 => n4447, A3 => n6890, ZN => 
                           n6891);
   U1355 : OAI211_X1 port map( C1 => n6893, C2 => n7748, A => n6892, B => n6891
                           , ZN => OUTALU(26));
   U1356 : AOI22_X1 port map( A1 => n7821, A2 => n2521_port, B1 => n7823, B2 =>
                           n3943, ZN => n2078);
   U1357 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n7105, ZN
                           => n2075);
   U1358 : OAI22_X1 port map( A1 => n4113, A2 => n6894, B1 => n4443, B2 => 
                           n6903, ZN => n6897);
   U1359 : AOI211_X1 port map( C1 => n4085, C2 => n4210, A => n4213, B => n4208
                           , ZN => n6896);
   U1360 : INV_X1 port map( A => n6940, ZN => n6924);
   U1361 : NOR3_X1 port map( A1 => n6924, A2 => n7725, A3 => n7748, ZN => n6895
                           );
   U1362 : AOI211_X1 port map( C1 => n4447, C2 => n6897, A => n6896, B => n6895
                           , ZN => n6900);
   U1363 : AOI21_X1 port map( B1 => n4085, B2 => n4202, A => n4419, ZN => n6898
                           );
   U1364 : NAND2_X1 port map( A1 => n7752, A2 => n6898, ZN => n6899);
   U1365 : NAND4_X1 port map( A1 => n3867, A2 => n3866, A3 => n6900, A4 => 
                           n6899, ZN => OUTALU(25));
   U1366 : AOI22_X1 port map( A1 => DATA1(24), A2 => n1945, B1 => DATA2(24), B2
                           => n1912, ZN => n7272);
   U1367 : INV_X1 port map( A => n7272, ZN => n6901);
   U1368 : AOI22_X1 port map( A1 => n3944, A2 => n7823, B1 => n7821, B2 => 
                           n6901, ZN => n2085);
   U1369 : INV_X1 port map( A => n1846, ZN => n6902);
   U1370 : NAND3_X1 port map( A1 => n6902, A2 => n1845, A3 => n2082, ZN => 
                           n2084);
   U1371 : OAI22_X1 port map( A1 => n6926, A2 => n7725, B1 => n6924, B2 => 
                           n7732, ZN => n6907);
   U1372 : NOR3_X1 port map( A1 => n4113, A2 => n4222, A3 => n6903, ZN => n6906
                           );
   U1373 : AOI22_X1 port map( A1 => n4417, A2 => n4393, B1 => n4449, B2 => 
                           n4526, ZN => n6904);
   U1374 : AOI21_X1 port map( B1 => n4224, B2 => n6904, A => n4491, ZN => n6905
                           );
   U1375 : AOI211_X1 port map( C1 => n7795, C2 => n6907, A => n6906, B => n6905
                           , ZN => n6909);
   U1376 : NAND2_X1 port map( A1 => n4417, A2 => n4209, ZN => n6908);
   U1377 : NAND4_X1 port map( A1 => n3865, A2 => n4075, A3 => n6909, A4 => 
                           n6908, ZN => OUTALU(24));
   U1378 : INV_X1 port map( A => DATA2(23), ZN => n7354);
   U1379 : NAND2_X1 port map( A1 => DATA1(23), A2 => n7354, ZN => n7215);
   U1380 : NAND2_X1 port map( A1 => DATA2(23), A2 => n1914, ZN => n7271);
   U1381 : AOI21_X1 port map( B1 => n7215, B2 => n7271, A => n7161, ZN => n2097
                           );
   U1382 : AOI21_X1 port map( B1 => DATA2(23), B2 => n1901, A => n1900, ZN => 
                           n2094);
   U1383 : INV_X1 port map( A => n1855, ZN => n7716);
   U1384 : AND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n6910);
   U1385 : AOI21_X1 port map( B1 => n6954, B2 => n1850, A => n6910, ZN => n7715
                           );
   U1386 : INV_X1 port map( A => n7715, ZN => n6947);
   U1387 : AOI21_X1 port map( B1 => n1849, B2 => n6947, A => n6911, ZN => n6913
                           );
   U1388 : AOI22_X1 port map( A1 => n6912, A2 => n7716, B1 => n1856, B2 => 
                           n6913, ZN => n2134);
   U1389 : INV_X1 port map( A => n6913, ZN => n6915);
   U1390 : AOI22_X1 port map( A1 => n1856, A2 => n6915, B1 => n7716, B2 => 
                           n6914, ZN => n1848);
   U1391 : INV_X1 port map( A => n6919, ZN => n6922);
   U1392 : INV_X1 port map( A => n6917, ZN => n6916);
   U1393 : AOI211_X1 port map( C1 => n1847, C2 => n2134, A => n6916, B => n7829
                           , ZN => n6921);
   U1394 : INV_X1 port map( A => n1847, ZN => n6918);
   U1395 : OAI22_X1 port map( A1 => n1848, A2 => n6918, B1 => n7829, B2 => 
                           n6917, ZN => n6920);
   U1396 : AOI22_X1 port map( A1 => n6922, A2 => n6921, B1 => n6920, B2 => 
                           n6919, ZN => n2116);
   U1397 : OAI22_X1 port map( A1 => n4507, A2 => n6923, B1 => n4098, B2 => 
                           n6934, ZN => n6931);
   U1398 : OAI22_X1 port map( A1 => n4460, A2 => n6948, B1 => n4094, B2 => 
                           n6955, ZN => n6930);
   U1399 : OAI222_X1 port map( A1 => n7732, A2 => n6926, B1 => n7725, B2 => 
                           n6925, C1 => n7763, C2 => n6924, ZN => n6927);
   U1400 : AOI21_X1 port map( B1 => n7795, B2 => n6927, A => n4074, ZN => n6928
                           );
   U1401 : NAND2_X1 port map( A1 => n3863, A2 => n6928, ZN => n6929);
   U1402 : AOI221_X1 port map( B1 => n6931, B2 => n4447, C1 => n6930, C2 => 
                           n4447, A => n6929, ZN => n6933);
   U1403 : NAND2_X1 port map( A1 => n4510, A2 => n3945, ZN => n6932);
   U1404 : OAI211_X1 port map( C1 => n4073, C2 => n4494, A => n6933, B => n6932
                           , ZN => OUTALU(23));
   U1405 : INV_X1 port map( A => DATA2(22), ZN => n7355);
   U1406 : AOI22_X1 port map( A1 => DATA1(22), A2 => DATA2(22), B1 => n7355, B2
                           => n7168, ZN => n7267);
   U1407 : AOI22_X1 port map( A1 => n3947, A2 => n7823, B1 => n7821, B2 => 
                           n7267, ZN => n2127);
   U1408 : OAI222_X1 port map( A1 => n4460, A2 => n6955, B1 => n4507, B2 => 
                           n6934, C1 => n4098, C2 => n6948, ZN => n6936);
   U1409 : OAI22_X1 port map( A1 => n4422, A2 => n4407, B1 => n4214, B2 => 
                           n3864, ZN => n6935);
   U1410 : AOI21_X1 port map( B1 => n4447, B2 => n6936, A => n6935, ZN => n6945
                           );
   U1411 : AOI22_X1 port map( A1 => n4289, A2 => n6938, B1 => n4489, B2 => 
                           n6937, ZN => n6942);
   U1412 : AOI22_X1 port map( A1 => n4474, A2 => n6940, B1 => n4480, B2 => 
                           n6939, ZN => n6941);
   U1413 : AOI21_X1 port map( B1 => n6942, B2 => n6941, A => n4251, ZN => n6943
                           );
   U1414 : NOR2_X1 port map( A1 => n6943, A2 => n3862, ZN => n6944);
   U1415 : NAND3_X1 port map( A1 => n3861, A2 => n6945, A3 => n6944, ZN => 
                           OUTALU(22));
   U1416 : AOI22_X1 port map( A1 => n1856, A2 => n6947, B1 => n7716, B2 => 
                           n6946, ZN => n2150);
   U1417 : AOI21_X1 port map( B1 => DATA2(21), B2 => n1901, A => n1900, ZN => 
                           n2144);
   U1418 : NOR2_X1 port map( A1 => DATA2(21), A2 => n1921, ZN => n7264);
   U1419 : NAND2_X1 port map( A1 => DATA2(21), A2 => n1921, ZN => n7213);
   U1420 : INV_X1 port map( A => n7213, ZN => n7268);
   U1421 : OR2_X1 port map( A1 => n7264, A2 => n7268, ZN => n7172);
   U1422 : AOI22_X1 port map( A1 => n7821, A2 => n7172, B1 => n7823, B2 => 
                           n3948, ZN => n2143);
   U1423 : OAI22_X1 port map( A1 => n4507, A2 => n6948, B1 => n4098, B2 => 
                           n6955, ZN => n6951);
   U1424 : INV_X1 port map( A => n7019, ZN => n7003);
   U1425 : NOR3_X1 port map( A1 => n7003, A2 => n7722, A3 => n7748, ZN => n6950
                           );
   U1426 : OAI22_X1 port map( A1 => n4086, A2 => n4406, B1 => n4072, B2 => 
                           n4493, ZN => n6949);
   U1427 : AOI211_X1 port map( C1 => n4447, C2 => n6951, A => n6950, B => n6949
                           , ZN => n6952);
   U1428 : OAI211_X1 port map( C1 => n4409, C2 => n3860, A => n3859, B => n6952
                           , ZN => OUTALU(21));
   U1429 : AOI22_X1 port map( A1 => n1856, A2 => n6954, B1 => n7716, B2 => 
                           n6953, ZN => n2165);
   U1430 : INV_X1 port map( A => DATA2(20), ZN => n7357);
   U1431 : OAI21_X1 port map( B1 => n7158, B2 => n7357, A => n7143, ZN => n2161
                           );
   U1432 : AOI22_X1 port map( A1 => DATA1(20), A2 => DATA2(20), B1 => n7357, B2
                           => n1922, ZN => n7179);
   U1433 : AOI22_X1 port map( A1 => n3949, A2 => n7823, B1 => n7821, B2 => 
                           n7179, ZN => n2157);
   U1434 : OAI22_X1 port map( A1 => n7001, A2 => n7722, B1 => n7003, B2 => 
                           n7755, ZN => n6959);
   U1435 : NOR3_X1 port map( A1 => n4507, A2 => n4222, A3 => n6955, ZN => n6958
                           );
   U1436 : NAND2_X1 port map( A1 => n4071, A2 => n4535, ZN => n6956);
   U1437 : OAI21_X1 port map( B1 => n4087, B2 => n3857, A => n6956, ZN => n6957
                           );
   U1438 : AOI211_X1 port map( C1 => n7795, C2 => n6959, A => n6958, B => n6957
                           , ZN => n6960);
   U1439 : OAI211_X1 port map( C1 => n4405, C2 => n3858, A => n3856, B => n6960
                           , ZN => OUTALU(20));
   U1440 : NOR2_X1 port map( A1 => DATA1(1), A2 => n7374, ZN => n7223);
   U1441 : INV_X1 port map( A => n7223, ZN => n6961);
   U1442 : NAND2_X1 port map( A1 => DATA1(1), A2 => n7374, ZN => n7225);
   U1443 : NAND2_X1 port map( A1 => n6961, A2 => n7225, ZN => n2513);
   U1444 : AOI211_X1 port map( C1 => n7159, C2 => n6972, A => n6962, B => n7162
                           , ZN => n6964);
   U1445 : AND2_X1 port map( A1 => n7823, A2 => n3794, ZN => n6963);
   U1446 : AOI211_X1 port map( C1 => n7821, C2 => n2513, A => n6964, B => n6963
                           , ZN => n2212);
   U1447 : AOI21_X1 port map( B1 => n7827, B2 => n1902, A => n1900, ZN => n7157
                           );
   U1448 : OAI21_X1 port map( B1 => n7374, B2 => n7158, A => n7157, ZN => n2204
                           );
   U1449 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(1), A => n6966, B => 
                           n6965, ZN => n6968);
   U1450 : OAI211_X1 port map( C1 => n7711, C2 => n7183, A => n6968, B => n6967
                           , ZN => n2435);
   U1451 : AOI222_X1 port map( A1 => n6971, A2 => n1068, B1 => n2433, B2 => 
                           n6970, C1 => n2435, C2 => n6969, ZN => n2425);
   U1452 : NAND3_X1 port map( A1 => DATA1(0), A2 => n7825, A3 => n1902, ZN => 
                           n2210);
   U1453 : OAI221_X1 port map( B1 => n7160, B2 => n6974, C1 => n6973, C2 => 
                           n6972, A => n7166, ZN => n2209);
   U1454 : AOI22_X1 port map( A1 => n4461, A2 => n6975, B1 => n4436, B2 => 
                           n7278, ZN => n6990);
   U1455 : OAI22_X1 port map( A1 => n4478, A2 => n3815, B1 => n4477, B2 => 
                           n3802, ZN => n6979);
   U1456 : OAI22_X1 port map( A1 => n4290, A2 => n6977, B1 => n6976, B2 => 
                           n7767, ZN => n6978);
   U1457 : AOI211_X1 port map( C1 => n6010, C2 => n7790, A => n6979, B => n6978
                           , ZN => n7286);
   U1458 : OAI22_X1 port map( A1 => n4245, A2 => n7286, B1 => n7284, B2 => 
                           n7755, ZN => n6982);
   U1459 : OAI22_X1 port map( A1 => n4476, A2 => n6980, B1 => n4101, B2 => 
                           n7287, ZN => n6981);
   U1460 : AOI211_X1 port map( C1 => n7727, C2 => n7290, A => n6982, B => n6981
                           , ZN => n7291);
   U1461 : OAI222_X1 port map( A1 => n4512, A2 => n6983, B1 => n4506, B2 => 
                           n7291, C1 => n7293, C2 => n4248, ZN => n7297);
   U1462 : AOI22_X1 port map( A1 => n4112, A2 => n7297, B1 => n6984, B2 => 
                           n7723, ZN => n6987);
   U1463 : AOI22_X1 port map( A1 => n4249, A2 => n6985, B1 => n4454, B2 => 
                           n7294, ZN => n6986);
   U1464 : OAI211_X1 port map( C1 => n6988, C2 => n7749, A => n6987, B => n6986
                           , ZN => n7301);
   U1465 : AOI22_X1 port map( A1 => n4110, A2 => n7301, B1 => n3921, B2 => 
                           n7279, ZN => n6989);
   U1466 : OAI211_X1 port map( C1 => n7305, C2 => n4098, A => n6990, B => n6989
                           , ZN => n7307);
   U1467 : AOI222_X1 port map( A1 => n7307, A2 => n4444, B1 => n7306, B2 => 
                           n4219, C1 => n6991, C2 => n3906, ZN => n7317);
   U1468 : OAI22_X1 port map( A1 => n7729, A2 => n7317, B1 => n4217, B2 => 
                           n7312, ZN => n6992);
   U1469 : INV_X1 port map( A => n6992, ZN => n6995);
   U1470 : AOI22_X1 port map( A1 => n4252, A2 => n6993, B1 => n4416, B2 => 
                           n7313, ZN => n6994);
   U1471 : OAI211_X1 port map( C1 => n7309, C2 => n7806, A => n6995, B => n6994
                           , ZN => n7347);
   U1472 : AOI22_X1 port map( A1 => n4070, A2 => n4531, B1 => n4508, B2 => 
                           n7347, ZN => n6996);
   U1473 : NAND4_X1 port map( A1 => n4069, A2 => n3822, A3 => n3854, A4 => 
                           n6996, ZN => OUTALU(1));
   U1474 : AOI22_X1 port map( A1 => n6998, A2 => n7716, B1 => n1856, B2 => 
                           n6997, ZN => n2226);
   U1475 : INV_X1 port map( A => DATA2(19), ZN => n7358);
   U1476 : OAI21_X1 port map( B1 => n7158, B2 => n7358, A => n7143, ZN => n6999
                           );
   U1477 : AOI22_X1 port map( A1 => DATA1(19), A2 => n6999, B1 => n7823, B2 => 
                           n3950, ZN => n2220);
   U1478 : NOR2_X1 port map( A1 => DATA2(19), A2 => n7000, ZN => n7209);
   U1479 : NAND2_X1 port map( A1 => DATA2(19), A2 => n7000, ZN => n7210);
   U1480 : INV_X1 port map( A => n7210, ZN => n7180);
   U1481 : OAI21_X1 port map( B1 => n7209, B2 => n7180, A => n7821, ZN => n2219
                           );
   U1482 : OAI222_X1 port map( A1 => n7719, A2 => n7003, B1 => n7722, B2 => 
                           n7002, C1 => n7755, C2 => n7001, ZN => n7009);
   U1483 : AOI22_X1 port map( A1 => n7736, A2 => n7004, B1 => n7796, B2 => 
                           n7021, ZN => n7006);
   U1484 : AOI22_X1 port map( A1 => n7723, A2 => n7036, B1 => n7733, B2 => 
                           n7044, ZN => n7005);
   U1485 : AOI21_X1 port map( B1 => n7006, B2 => n7005, A => n7803, ZN => n7008
                           );
   U1486 : OAI22_X1 port map( A1 => n4404, A2 => n4403, B1 => n4090, B2 => 
                           n3852, ZN => n7007);
   U1487 : AOI211_X1 port map( C1 => n7795, C2 => n7009, A => n7008, B => n7007
                           , ZN => n7010);
   U1488 : NAND3_X1 port map( A1 => n3851, A2 => n4068, A3 => n7010, ZN => 
                           OUTALU(19));
   U1489 : INV_X1 port map( A => DATA2(18), ZN => n7359);
   U1490 : OAI21_X1 port map( B1 => n7158, B2 => n7359, A => n7143, ZN => n2245
                           );
   U1491 : NAND2_X1 port map( A1 => n7012, A2 => n7011, ZN => n7016);
   U1492 : INV_X1 port map( A => n7016, ZN => n7014);
   U1493 : AOI211_X1 port map( C1 => n7014, C2 => n7032, A => n7013, B => n1855
                           , ZN => n2244);
   U1494 : NAND2_X1 port map( A1 => DATA2(18), A2 => n1925, ZN => n7181);
   U1495 : OAI21_X1 port map( B1 => DATA2(18), B2 => n1925, A => n7181, ZN => 
                           n7263);
   U1496 : AOI22_X1 port map( A1 => n3951, A2 => n7823, B1 => n7821, B2 => 
                           n7263, ZN => n2240);
   U1497 : OAI211_X1 port map( C1 => n7030, C2 => n7016, A => n1856, B => n7015
                           , ZN => n2250);
   U1498 : AOI22_X1 port map( A1 => n4518, A2 => n7018, B1 => n4466, B2 => 
                           n7017, ZN => n7026);
   U1499 : AOI22_X1 port map( A1 => n4468, A2 => n7020, B1 => n4243, B2 => 
                           n7019, ZN => n7025);
   U1500 : AOI222_X1 port map( A1 => n7796, A2 => n7036, B1 => n7021, B2 => 
                           n7736, C1 => n7044, C2 => n7723, ZN => n7022);
   U1501 : OAI211_X1 port map( C1 => n4222, C2 => n7022, A => n3848, B => n3849
                           , ZN => n7023);
   U1502 : AOI211_X1 port map( C1 => n4067, C2 => n4534, A => n3850, B => n7023
                           , ZN => n7024);
   U1503 : OAI221_X1 port map( B1 => n4251, B2 => n7026, C1 => n4251, C2 => 
                           n7025, A => n7024, ZN => OUTALU(18));
   U1504 : NOR2_X1 port map( A1 => DATA2(17), A2 => n7027, ZN => n7260);
   U1505 : INV_X1 port map( A => n7260, ZN => n7028);
   U1506 : NAND2_X1 port map( A1 => DATA2(17), A2 => n7027, ZN => n7258);
   U1507 : NAND2_X1 port map( A1 => n7028, A2 => n7258, ZN => n7171);
   U1508 : AOI22_X1 port map( A1 => n7821, A2 => n7171, B1 => n7823, B2 => 
                           n3952, ZN => n2267);
   U1509 : AOI211_X1 port map( C1 => n7031, C2 => n7034, A => n7030, B => n7029
                           , ZN => n2262);
   U1510 : NAND2_X1 port map( A1 => DATA2_I_16_port, A2 => DATA1(16), ZN => 
                           n7035);
   U1511 : INV_X1 port map( A => n7032, ZN => n7033);
   U1512 : AOI211_X1 port map( C1 => n7035, C2 => n7034, A => n7033, B => n1855
                           , ZN => n2261);
   U1513 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n7105, ZN
                           => n2264);
   U1514 : AOI22_X1 port map( A1 => n7736, A2 => n7036, B1 => n7796, B2 => 
                           n7044, ZN => n7037);
   U1515 : INV_X1 port map( A => n7037, ZN => n7038);
   U1516 : AOI211_X1 port map( C1 => n4447, C2 => n7038, A => n3846, B => n3845
                           , ZN => n7040);
   U1517 : NAND3_X1 port map( A1 => n4455, A2 => n4508, A3 => n7043, ZN => 
                           n7039);
   U1518 : NAND4_X1 port map( A1 => n3847, A2 => n3844, A3 => n7040, A4 => 
                           n7039, ZN => OUTALU(17));
   U1519 : OAI21_X1 port map( B1 => n7158, B2 => n7361, A => n7143, ZN => n2275
                           );
   U1520 : AOI22_X1 port map( A1 => n3953, A2 => n7823, B1 => n7821, B2 => 
                           n7041, ZN => n2271);
   U1521 : AOI22_X1 port map( A1 => n4456, A2 => n7043, B1 => n4455, B2 => 
                           n7042, ZN => n7049);
   U1522 : NOR2_X1 port map( A1 => n4402, A2 => n4201, ZN => n7047);
   U1523 : NAND3_X1 port map( A1 => n7736, A2 => n7798, A3 => n7044, ZN => 
                           n7045);
   U1524 : OAI211_X1 port map( C1 => n4089, C2 => n4408, A => n3843, B => n7045
                           , ZN => n7046);
   U1525 : AOI211_X1 port map( C1 => n4066, C2 => n4533, A => n7047, B => n7046
                           , ZN => n7048);
   U1526 : OAI21_X1 port map( B1 => n4251, B2 => n7049, A => n7048, ZN => 
                           OUTALU(16));
   U1527 : NAND2_X1 port map( A1 => DATA1(11), A2 => DATA2_I_11_port, ZN => 
                           n7054);
   U1528 : OAI21_X1 port map( B1 => n7051, B2 => n7146, A => n7050, ZN => n7140
                           );
   U1529 : NAND2_X1 port map( A1 => n7052, A2 => n7140, ZN => n7128);
   U1530 : NAND2_X1 port map( A1 => n7133, A2 => n7128, ZN => n7053);
   U1531 : NAND2_X1 port map( A1 => n7054, A2 => n7053, ZN => n7107);
   U1532 : AOI21_X1 port map( B1 => n7056, B2 => n7107, A => n7055, ZN => n7075
                           );
   U1533 : OAI221_X1 port map( B1 => n2323, B2 => n7075, C1 => n2323, C2 => 
                           n7074, A => n7057, ZN => n7058);
   U1534 : XNOR2_X1 port map( A => n7063, B => n7058, ZN => n7062);
   U1535 : NAND3_X1 port map( A1 => DATA2(15), A2 => DATA1(15), A3 => n7105, ZN
                           => n7061);
   U1536 : NOR2_X1 port map( A1 => DATA2(15), A2 => n7695, ZN => n7203);
   U1537 : OAI21_X1 port map( B1 => n7203, B2 => n7059, A => n7821, ZN => n7060
                           );
   U1538 : OAI211_X1 port map( C1 => n7062, C2 => n1859, A => n7061, B => n7060
                           , ZN => n2294);
   U1539 : INV_X1 port map( A => n7064, ZN => n7066);
   U1540 : INV_X1 port map( A => n7063, ZN => n7065);
   U1541 : OAI221_X1 port map( B1 => n7066, B2 => n7065, C1 => n7064, C2 => 
                           n7063, A => n1860, ZN => n2300);
   U1542 : OAI22_X1 port map( A1 => n7067, A2 => n7720, B1 => n7083, B2 => 
                           n7730, ZN => n7068);
   U1543 : AOI22_X1 port map( A1 => n3954, A2 => n4510, B1 => n7798, B2 => 
                           n7068, ZN => n7071);
   U1544 : NOR3_X1 port map( A1 => n4464, A2 => n7082, A3 => n4251, ZN => n7069
                           );
   U1545 : NOR2_X1 port map( A1 => n7069, A2 => n3842, ZN => n7070);
   U1546 : NAND3_X1 port map( A1 => n3821, A2 => n7071, A3 => n7070, ZN => 
                           OUTALU(15));
   U1547 : AND2_X1 port map( A1 => n7075, A2 => n7074, ZN => n7072);
   U1548 : OAI22_X1 port map( A1 => n7073, A2 => n7129, B1 => n7072, B2 => 
                           n1859, ZN => n2322);
   U1549 : INV_X1 port map( A => n7074, ZN => n7077);
   U1550 : AOI22_X1 port map( A1 => n7076, A2 => n1860, B1 => n7147, B2 => 
                           n7075, ZN => n7093);
   U1551 : NOR3_X1 port map( A1 => n7077, A2 => n7093, A3 => n2323, ZN => n2321
                           );
   U1552 : NAND2_X1 port map( A1 => n4319, A2 => n4314, ZN => n7078);
   U1553 : OAI21_X1 port map( B1 => n4319, B2 => n4314, A => n7078, ZN => n7607
                           );
   U1554 : NOR3_X1 port map( A1 => n7607, A2 => n7746, A3 => n7777, ZN => n3020
                           );
   U1555 : INV_X1 port map( A => n7607, ZN => n7606);
   U1556 : NAND2_X1 port map( A1 => n7606, A2 => n4329, ZN => n7079);
   U1557 : AOI21_X1 port map( B1 => n7079, B2 => n7777, A => n3020, ZN => n2313
                           );
   U1558 : OAI21_X1 port map( B1 => n7158, B2 => n7080, A => n7143, ZN => n7081
                           );
   U1559 : AOI22_X1 port map( A1 => DATA2(14), A2 => n7081, B1 => n7823, B2 => 
                           n4200, ZN => n2319);
   U1560 : INV_X1 port map( A => n7082, ZN => n7119);
   U1561 : AOI22_X1 port map( A1 => n4112, A2 => n7118, B1 => n4454, B2 => 
                           n7119, ZN => n7089);
   U1562 : NOR3_X1 port map( A1 => n7083, A2 => n7720, A3 => n7803, ZN => n7087
                           );
   U1563 : NOR2_X1 port map( A1 => n4254, A2 => n3840, ZN => n7084);
   U1564 : AOI21_X1 port map( B1 => n3841, B2 => n4088, A => n7084, ZN => n7085
                           );
   U1565 : NAND2_X1 port map( A1 => n7085, A2 => n3839, ZN => n7086);
   U1566 : NOR3_X1 port map( A1 => n7087, A2 => n4065, A3 => n7086, ZN => n7088
                           );
   U1567 : OAI21_X1 port map( B1 => n4251, B2 => n7089, A => n7088, ZN => 
                           OUTALU(14));
   U1568 : INV_X1 port map( A => n7111, ZN => n7113);
   U1569 : AOI211_X1 port map( C1 => n7091, C2 => n7110, A => n7090, B => n7829
                           , ZN => n7092);
   U1570 : NAND3_X1 port map( A1 => n7113, A2 => n7092, A3 => n7107, ZN => 
                           n2340);
   U1571 : OAI21_X1 port map( B1 => n7158, B2 => n7364, A => n7143, ZN => n2338
                           );
   U1572 : AOI21_X1 port map( B1 => n7095, B2 => n7094, A => n7093, ZN => n2337
                           );
   U1573 : NOR2_X1 port map( A1 => DATA2(13), A2 => n1933, ZN => n7253);
   U1574 : INV_X1 port map( A => n7253, ZN => n7096);
   U1575 : NAND2_X1 port map( A1 => DATA2(13), A2 => n1933, ZN => n7251);
   U1576 : NAND2_X1 port map( A1 => n7096, A2 => n7251, ZN => n7170);
   U1577 : AOI22_X1 port map( A1 => n7821, A2 => n7170, B1 => n7823, B2 => 
                           n3970, ZN => n2333);
   U1578 : INV_X1 port map( A => n7114, ZN => n7098);
   U1579 : AOI22_X1 port map( A1 => n4518, A2 => n7098, B1 => n4466, B2 => 
                           n7097, ZN => n7104);
   U1580 : OAI22_X1 port map( A1 => n7719, A2 => n7134, B1 => n7759, B2 => 
                           n7152, ZN => n7099);
   U1581 : INV_X1 port map( A => n7099, ZN => n7103);
   U1582 : AOI222_X1 port map( A1 => n7116, A2 => n4112, B1 => n7118, B2 => 
                           n4454, C1 => n7119, C2 => n4114, ZN => n7100);
   U1583 : OAI211_X1 port map( C1 => n4251, C2 => n7100, A => n3838, B => n3837
                           , ZN => n7101);
   U1584 : AOI211_X1 port map( C1 => n4064, C2 => n4532, A => n4063, B => n7101
                           , ZN => n7102);
   U1585 : OAI221_X1 port map( B1 => n4222, B2 => n7104, C1 => n4222, C2 => 
                           n7103, A => n7102, ZN => OUTALU(13));
   U1586 : NAND3_X1 port map( A1 => DATA2(12), A2 => DATA1(12), A3 => n7105, ZN
                           => n7109);
   U1587 : INV_X1 port map( A => n7107, ZN => n7106);
   U1588 : OAI221_X1 port map( B1 => n7113, B2 => n7107, C1 => n7111, C2 => 
                           n7106, A => n7147, ZN => n7108);
   U1589 : OAI211_X1 port map( C1 => n7247, C2 => n7161, A => n7109, B => n7108
                           , ZN => n2355);
   U1590 : OAI221_X1 port map( B1 => n7113, B2 => n7112, C1 => n7111, C2 => 
                           n7110, A => n1860, ZN => n2361);
   U1591 : OAI222_X1 port map( A1 => n7719, A2 => n7152, B1 => n7722, B2 => 
                           n7114, C1 => n7755, C2 => n7134, ZN => n7115);
   U1592 : AOI22_X1 port map( A1 => n4263, A2 => n4510, B1 => n7798, B2 => 
                           n7115, ZN => n7124);
   U1593 : AOI22_X1 port map( A1 => n4112, A2 => n7117, B1 => n4454, B2 => 
                           n7116, ZN => n7121);
   U1594 : AOI22_X1 port map( A1 => n4453, A2 => n7119, B1 => n4114, B2 => 
                           n7118, ZN => n7120);
   U1595 : AOI21_X1 port map( B1 => n7121, B2 => n7120, A => n4251, ZN => n7122
                           );
   U1596 : NOR2_X1 port map( A1 => n7122, A2 => n3836, ZN => n7123);
   U1597 : NAND3_X1 port map( A1 => n3835, A2 => n7124, A3 => n7123, ZN => 
                           OUTALU(12));
   U1598 : AOI211_X1 port map( C1 => n7143, C2 => n7158, A => n7125, B => n7366
                           , ZN => n7127);
   U1599 : NAND2_X1 port map( A1 => DATA1(11), A2 => n7366, ZN => n7196);
   U1600 : AOI21_X1 port map( B1 => n7196, B2 => n7246, A => n7161, ZN => n7126
                           );
   U1601 : AOI211_X1 port map( C1 => n3986, C2 => n7823, A => n7127, B => n7126
                           , ZN => n2381);
   U1602 : INV_X1 port map( A => n7133, ZN => n7131);
   U1603 : XNOR2_X1 port map( A => n7131, B => n7128, ZN => n2379);
   U1604 : INV_X1 port map( A => n7132, ZN => n7130);
   U1605 : AOI221_X1 port map( B1 => n7133, B2 => n7132, C1 => n7131, C2 => 
                           n7130, A => n7129, ZN => n2378);
   U1606 : OAI22_X1 port map( A1 => n7134, A2 => n7722, B1 => n7152, B2 => 
                           n7755, ZN => n7135);
   U1607 : AOI22_X1 port map( A1 => n4199, A2 => n4226, B1 => n7798, B2 => 
                           n7135, ZN => n7138);
   U1608 : NOR3_X1 port map( A1 => n4507, A2 => n7148, A3 => n4251, ZN => n7136
                           );
   U1609 : NOR2_X1 port map( A1 => n7136, A2 => n3820, ZN => n7137);
   U1610 : NAND3_X1 port map( A1 => n4062, A2 => n7138, A3 => n7137, ZN => 
                           OUTALU(11));
   U1611 : NAND2_X1 port map( A1 => n1860, A2 => n7139, ZN => n2401);
   U1612 : NAND2_X1 port map( A1 => n7147, A2 => n7140, ZN => n7141);
   U1613 : AOI22_X1 port map( A1 => n7142, A2 => n7145, B1 => n7141, B2 => 
                           n2401, ZN => n2403);
   U1614 : OAI21_X1 port map( B1 => n7158, B2 => n7367, A => n7143, ZN => n7144
                           );
   U1615 : AOI22_X1 port map( A1 => DATA1(10), A2 => DATA2(10), B1 => n7367, B2
                           => n7167, ZN => n7243);
   U1616 : AOI22_X1 port map( A1 => DATA1(10), A2 => n7144, B1 => n7821, B2 => 
                           n7243, ZN => n2399);
   U1617 : NAND3_X1 port map( A1 => n7147, A2 => n7146, A3 => n7145, ZN => 
                           n2407);
   U1618 : OAI22_X1 port map( A1 => n7149, A2 => n7751, B1 => n7148, B2 => 
                           n7805, ZN => n7151);
   U1619 : OAI21_X1 port map( B1 => n4198, B2 => n4423, A => n3833, ZN => n7150
                           );
   U1620 : AOI211_X1 port map( C1 => n7795, C2 => n7151, A => n3834, B => n7150
                           , ZN => n7155);
   U1621 : OR3_X1 port map( A1 => n7722, A2 => n7803, A3 => n7152, ZN => n7154)
                           ;
   U1622 : NAND2_X1 port map( A1 => n4510, A2 => n4266, ZN => n7153);
   U1623 : NAND4_X1 port map( A1 => n4061, A2 => n7155, A3 => n7154, A4 => 
                           n7153, ZN => OUTALU(10));
   U1624 : NOR2_X1 port map( A1 => DATA1(0), A2 => n7658, ZN => n7184);
   U1625 : NAND2_X1 port map( A1 => DATA1(0), A2 => n7658, ZN => n7224);
   U1626 : INV_X1 port map( A => n7224, ZN => n7156);
   U1627 : NOR2_X1 port map( A1 => n7184, A2 => n7156, ZN => n1940);
   U1628 : OAI21_X1 port map( B1 => n7658, B2 => n7158, A => n7157, ZN => n7164
                           );
   U1629 : NOR2_X1 port map( A1 => n7160, A2 => n7159, ZN => n7165);
   U1630 : OAI22_X1 port map( A1 => n7165, A2 => n7162, B1 => n1940, B2 => 
                           n7161, ZN => n7163);
   U1631 : AOI21_X1 port map( B1 => DATA1(0), B2 => n7164, A => n7163, ZN => 
                           n2694);
   U1632 : AOI22_X1 port map( A1 => n7166, A2 => n7165, B1 => n7823, B2 => 
                           n4192, ZN => n2693);
   U1633 : OAI21_X1 port map( B1 => DATA2(26), B2 => n1910, A => n2594, ZN => 
                           n2671);
   U1634 : OAI21_X1 port map( B1 => DATA2(10), B2 => n7167, A => n7196, ZN => 
                           n7248);
   U1635 : OAI21_X1 port map( B1 => DATA2(22), B2 => n7168, A => n7215, ZN => 
                           n7273);
   U1636 : AOI21_X1 port map( B1 => DATA1(14), B2 => n7363, A => n7203, ZN => 
                           n7256);
   U1637 : AOI21_X1 port map( B1 => DATA1(18), B2 => n7359, A => n7209, ZN => 
                           n7261);
   U1638 : NAND2_X1 port map( A1 => n7256, A2 => n7261, ZN => n7169);
   U1639 : NOR3_X1 port map( A1 => n7248, A2 => n7273, A3 => n7169, ZN => 
                           n2529_port);
   U1640 : NOR4_X1 port map( A1 => n7173, A2 => n7172, A3 => n7171, A4 => n7170
                           , ZN => n2527_port);
   U1641 : INV_X1 port map( A => n7238, ZN => n7178);
   U1642 : AOI22_X1 port map( A1 => DATA2(6), A2 => n7175, B1 => DATA2(7), B2 
                           => n7174, ZN => n7190);
   U1643 : NAND4_X1 port map( A1 => n7178, A2 => n7177, A3 => n7176, A4 => 
                           n7190, ZN => n2541_port);
   U1644 : INV_X1 port map( A => DATA2(26), ZN => n7352);
   U1645 : OAI21_X1 port map( B1 => DATA1(26), B2 => n7352, A => n2669, ZN => 
                           n2595);
   U1646 : OAI21_X1 port map( B1 => DATA1(22), B2 => n7355, A => n7271, ZN => 
                           n7216);
   U1647 : INV_X1 port map( A => n7216, ZN => n7182);
   U1648 : NOR2_X1 port map( A1 => n7180, A2 => n7179, ZN => n7266);
   U1649 : NAND4_X1 port map( A1 => n7272, A2 => n7182, A3 => n7266, A4 => 
                           n7181, ZN => n2539_port);
   U1650 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2(26), B1 => n7352, B2
                           => n1910, ZN => n1909);
   U1651 : AOI21_X1 port map( B1 => DATA1(14), B2 => n7363, A => n7201, ZN => 
                           n2635);
   U1652 : AOI22_X1 port map( A1 => DATA2(25), A2 => n1911, B1 => DATA2(24), B2
                           => n1912, ZN => n7219);
   U1653 : AOI22_X1 port map( A1 => DATA2(12), A2 => n7687, B1 => DATA2(13), B2
                           => n1933, ZN => n7200);
   U1654 : NOR2_X1 port map( A1 => DATA2(4), A2 => n7183, ZN => n7237);
   U1655 : AOI22_X1 port map( A1 => n7184, A2 => n7225, B1 => DATA2(1), B2 => 
                           n1939, ZN => n7185);
   U1656 : OAI22_X1 port map( A1 => DATA1(2), A2 => n1970, B1 => n7185, B2 => 
                           n7222, ZN => n7186);
   U1657 : OAI21_X1 port map( B1 => n7233, B2 => n7186, A => n7226, ZN => n7187
                           );
   U1658 : OAI211_X1 port map( C1 => n7237, C2 => n7187, A => n7228, B => n7234
                           , ZN => n7188);
   U1659 : NAND3_X1 port map( A1 => n7235, A2 => n7231, A3 => n7188, ZN => 
                           n7189);
   U1660 : AOI21_X1 port map( B1 => n7190, B2 => n7189, A => n7238, ZN => n7193
                           );
   U1661 : AOI22_X1 port map( A1 => n7193, A2 => n7192, B1 => DATA2(8), B2 => 
                           n7191, ZN => n7195);
   U1662 : AOI211_X1 port map( C1 => n7195, C2 => n7194, A => n7242, B => n7243
                           , ZN => n7198);
   U1663 : OAI211_X1 port map( C1 => n7198, C2 => n7197, A => n7247, B => n7196
                           , ZN => n7199);
   U1664 : AOI21_X1 port map( B1 => n7200, B2 => n7199, A => n7253, ZN => n7202
                           );
   U1665 : AOI21_X1 port map( B1 => n2635, B2 => n7202, A => n7201, ZN => n7205
                           );
   U1666 : AOI21_X1 port map( B1 => n7205, B2 => n7204, A => n7203, ZN => n7206
                           );
   U1667 : NAND2_X1 port map( A1 => DATA1(16), A2 => n7361, ZN => n7254);
   U1668 : AOI22_X1 port map( A1 => n7206, A2 => n7254, B1 => DATA2(16), B2 => 
                           n1929, ZN => n7207);
   U1669 : AOI211_X1 port map( C1 => n7207, C2 => n7258, A => n7260, B => n7263
                           , ZN => n7208);
   U1670 : AOI21_X1 port map( B1 => DATA2(18), B2 => n1925, A => n7208, ZN => 
                           n7211);
   U1671 : AOI21_X1 port map( B1 => n7211, B2 => n7210, A => n7209, ZN => n7212
                           );
   U1672 : NAND2_X1 port map( A1 => DATA1(20), A2 => n7357, ZN => n7269);
   U1673 : AOI22_X1 port map( A1 => n7212, A2 => n7269, B1 => DATA2(20), B2 => 
                           n1922, ZN => n7214);
   U1674 : AOI211_X1 port map( C1 => n7214, C2 => n7213, A => n7264, B => n7267
                           , ZN => n7217);
   U1675 : OAI211_X1 port map( C1 => n7217, C2 => n7216, A => n7272, B => n7215
                           , ZN => n7218);
   U1676 : AOI211_X1 port map( C1 => n7219, C2 => n7218, A => n7221, B => n1909
                           , ZN => n2596);
   U1677 : AOI21_X1 port map( B1 => DATA1(6), B2 => n7372, A => n7220, ZN => 
                           n2622);
   U1678 : AOI21_X1 port map( B1 => DATA1(24), B2 => n1945, A => n7221, ZN => 
                           n7277);
   U1679 : AOI211_X1 port map( C1 => n7225, C2 => n7224, A => n7223, B => n7222
                           , ZN => n7230);
   U1680 : OAI21_X1 port map( B1 => DATA2(2), B2 => n7227, A => n7226, ZN => 
                           n7229);
   U1681 : OAI21_X1 port map( B1 => n7230, B2 => n7229, A => n7228, ZN => n7232
                           );
   U1682 : OAI21_X1 port map( B1 => n7233, B2 => n7232, A => n7231, ZN => n7236
                           );
   U1683 : OAI211_X1 port map( C1 => n7237, C2 => n7236, A => n7235, B => n7234
                           , ZN => n7240);
   U1684 : NOR2_X1 port map( A1 => DATA1(7), A2 => n1946, ZN => n7239);
   U1685 : AOI211_X1 port map( C1 => n2622, C2 => n7240, A => n7239, B => n7238
                           , ZN => n7241);
   U1686 : AOI211_X1 port map( C1 => DATA1(8), C2 => n7369, A => n7242, B => 
                           n7241, ZN => n7244);
   U1687 : NOR3_X1 port map( A1 => n7245, A2 => n7244, A3 => n7243, ZN => n7249
                           );
   U1688 : OAI211_X1 port map( C1 => n7249, C2 => n7248, A => n7247, B => n7246
                           , ZN => n7250);
   U1689 : OAI21_X1 port map( B1 => DATA2(12), B2 => n7687, A => n7250, ZN => 
                           n7252);
   U1690 : OAI211_X1 port map( C1 => n7253, C2 => n7252, A => n2635, B => n7251
                           , ZN => n7255);
   U1691 : OAI221_X1 port map( B1 => n7257, B2 => n7256, C1 => n7257, C2 => 
                           n7255, A => n7254, ZN => n7259);
   U1692 : OAI21_X1 port map( B1 => n7260, B2 => n7259, A => n7258, ZN => n7262
                           );
   U1693 : OAI21_X1 port map( B1 => n7263, B2 => n7262, A => n7261, ZN => n7265
                           );
   U1694 : AOI21_X1 port map( B1 => n7266, B2 => n7265, A => n7264, ZN => n7270
                           );
   U1695 : AOI211_X1 port map( C1 => n7270, C2 => n7269, A => n7268, B => n7267
                           , ZN => n7274);
   U1696 : OAI211_X1 port map( C1 => n7274, C2 => n7273, A => n7272, B => n7271
                           , ZN => n7276);
   U1697 : AOI211_X1 port map( C1 => n7277, C2 => n7276, A => n7275, B => n1909
                           , ZN => n2672);
   U1698 : AOI22_X1 port map( A1 => n4436, A2 => n7279, B1 => n4461, B2 => 
                           n7278, ZN => n7304);
   U1699 : OAI22_X1 port map( A1 => n4102, A2 => n3815, B1 => n7778, B2 => 
                           n7732, ZN => n7282);
   U1700 : AOI222_X1 port map( A1 => n4517, A2 => n3873, B1 => n4498, B2 => 
                           n3853, C1 => n4401, C2 => n4486, ZN => n7280);
   U1701 : OAI22_X1 port map( A1 => n4478, A2 => n3802, B1 => n4519, B2 => 
                           n7280, ZN => n7281);
   U1702 : AOI211_X1 port map( C1 => n7740, C2 => n7283, A => n7282, B => n7281
                           , ZN => n7285);
   U1703 : OAI22_X1 port map( A1 => n4245, A2 => n7285, B1 => n4101, B2 => 
                           n7284, ZN => n7289);
   U1704 : OAI22_X1 port map( A1 => n4472, A2 => n7287, B1 => n7286, B2 => 
                           n7755, ZN => n7288);
   U1705 : AOI211_X1 port map( C1 => n7761, C2 => n7290, A => n7289, B => n7288
                           , ZN => n7292);
   U1706 : OAI222_X1 port map( A1 => n4512, A2 => n7293, B1 => n4506, B2 => 
                           n7292, C1 => n4248, C2 => n7291, ZN => n7295);
   U1707 : AOI22_X1 port map( A1 => n4112, A2 => n7295, B1 => n4114, B2 => 
                           n7294, ZN => n7299);
   U1708 : AOI22_X1 port map( A1 => n4454, A2 => n7297, B1 => n4249, B2 => 
                           n7296, ZN => n7298);
   U1709 : OAI211_X1 port map( C1 => n7300, C2 => n4234, A => n7299, B => n7298
                           , ZN => n7302);
   U1710 : AOI22_X1 port map( A1 => n4110, A2 => n7302, B1 => n7800, B2 => 
                           n7301, ZN => n7303);
   U1711 : OAI211_X1 port map( C1 => n7305, C2 => n7799, A => n7304, B => n7303
                           , ZN => n7308);
   U1712 : AOI222_X1 port map( A1 => n7308, A2 => n4444, B1 => n7307, B2 => 
                           n4219, C1 => n7306, C2 => n3906, ZN => n7310);
   U1713 : OAI22_X1 port map( A1 => n7729, A2 => n7310, B1 => n7753, B2 => 
                           n7309, ZN => n7311);
   U1714 : INV_X1 port map( A => n7311, ZN => n7316);
   U1715 : INV_X1 port map( A => n7312, ZN => n7314);
   U1716 : AOI22_X1 port map( A1 => n4416, A2 => n7314, B1 => n4252, B2 => 
                           n7313, ZN => n7315);
   U1717 : OAI211_X1 port map( C1 => n7317, C2 => n4440, A => n7316, B => n7315
                           , ZN => n7346);
   U1718 : NOR4_X1 port map( A1 => n4076, A2 => n4253, A3 => n3901, A4 => n3832
                           , ZN => n7321);
   U1719 : NOR2_X1 port map( A1 => n4057, A2 => n3826, ZN => n7318);
   U1720 : NAND3_X1 port map( A1 => n3871, A2 => n3829, A3 => n7318, ZN => 
                           n7319);
   U1721 : NOR3_X1 port map( A1 => n3828, A2 => n3827, A3 => n7319, ZN => n7320
                           );
   U1722 : NAND4_X1 port map( A1 => n7321, A2 => n3830, A3 => n4056, A4 => 
                           n7320, ZN => n7322);
   U1723 : NOR4_X1 port map( A1 => n4058, A2 => n3855, A3 => n7323, A4 => n7322
                           , ZN => n7326);
   U1724 : NAND2_X1 port map( A1 => n5995, A2 => n4530, ZN => n7325);
   U1725 : INV_X1 port map( A => n7341, ZN => n7324);
   U1726 : NAND4_X1 port map( A1 => n7327, A2 => n7326, A3 => n7325, A4 => 
                           n7324, ZN => n7328);
   U1727 : NAND2_X1 port map( A1 => n4513, A2 => n7328, ZN => n7329);
   U1728 : AOI211_X1 port map( C1 => n4546, C2 => n7329, A => n4548, B => n4400
                           , ZN => n7345);
   U1729 : AOI21_X1 port map( B1 => n4529, B2 => n6022, A => n7341, ZN => n7333
                           );
   U1730 : NAND2_X1 port map( A1 => n4540, A2 => n4414, ZN => n7334);
   U1731 : NAND2_X1 port map( A1 => n6016, A2 => n4528, ZN => n7336);
   U1732 : OAI211_X1 port map( C1 => n3825, C2 => n4057, A => n3871, B => n4203
                           , ZN => n7330);
   U1733 : OAI211_X1 port map( C1 => n4539, C2 => n4413, A => n7336, B => n7330
                           , ZN => n7331);
   U1734 : NAND3_X1 port map( A1 => n7338, A2 => n7334, A3 => n7331, ZN => 
                           n7332);
   U1735 : AOI22_X1 port map( A1 => n5995, A2 => n4530, B1 => n7333, B2 => 
                           n7332, ZN => n7343);
   U1736 : AOI22_X1 port map( A1 => n5995, A2 => n4530, B1 => n4542, B2 => 
                           n4415, ZN => n7340);
   U1737 : OAI211_X1 port map( C1 => n3824, C2 => n4059, A => n3871, B => n4204
                           , ZN => n7335);
   U1738 : OAI211_X1 port map( C1 => n4527, C2 => n4457, A => n7335, B => n7334
                           , ZN => n7337);
   U1739 : NAND3_X1 port map( A1 => n7338, A2 => n7337, A3 => n7336, ZN => 
                           n7339);
   U1740 : OAI221_X1 port map( B1 => n7341, B2 => n7340, C1 => n7341, C2 => 
                           n7339, A => n7816, ZN => n7342);
   U1741 : OAI211_X1 port map( C1 => n4545, C2 => n7343, A => n4514, B => n7342
                           , ZN => n7344);
   U1742 : AOI22_X1 port map( A1 => n4508, A2 => n7346, B1 => n7345, B2 => 
                           n7344, ZN => n7349);
   U1743 : NAND3_X1 port map( A1 => n4545, A2 => n4205, A3 => n7347, ZN => 
                           n7348);
   U1744 : NAND4_X1 port map( A1 => n4060, A2 => n3831, A3 => n7349, A4 => 
                           n7348, ZN => OUTALU(0));
   U1745 : NAND2_X1 port map( A1 => n7350, A2 => n1905, ZN => n7376);
   U1746 : CLKBUF_X1 port map( A => n7376, Z => n7371);
   U1747 : NAND2_X1 port map( A1 => n7350, A2 => FUNC(3), ZN => n7375);
   U1748 : AOI22_X1 port map( A1 => DATA2(31), A2 => n7371, B1 => n7370, B2 => 
                           n1941, ZN => N2548);
   U1749 : AOI22_X1 port map( A1 => DATA2(30), A2 => n7376, B1 => n7375, B2 => 
                           n1942, ZN => N2547);
   U1750 : AOI22_X1 port map( A1 => DATA2(29), A2 => n7371, B1 => n7370, B2 => 
                           n1943, ZN => N2546);
   U1751 : AOI22_X1 port map( A1 => DATA2(28), A2 => n7376, B1 => n7375, B2 => 
                           n1944, ZN => N2545);
   U1752 : AOI22_X1 port map( A1 => DATA2(27), A2 => n7371, B1 => n7370, B2 => 
                           n7351, ZN => N2544);
   U1753 : AOI22_X1 port map( A1 => DATA2(26), A2 => n7376, B1 => n7375, B2 => 
                           n7352, ZN => N2543);
   U1754 : AOI22_X1 port map( A1 => DATA2(25), A2 => n7371, B1 => n7370, B2 => 
                           n7353, ZN => N2542);
   U1755 : AOI22_X1 port map( A1 => DATA2(24), A2 => n7376, B1 => n7375, B2 => 
                           n1945, ZN => N2541);
   U1756 : AOI22_X1 port map( A1 => DATA2(23), A2 => n7371, B1 => n7370, B2 => 
                           n7354, ZN => N2540);
   U1757 : AOI22_X1 port map( A1 => DATA2(22), A2 => n7376, B1 => n7375, B2 => 
                           n7355, ZN => N2539);
   U1758 : INV_X1 port map( A => DATA2(21), ZN => n7356);
   U1759 : AOI22_X1 port map( A1 => DATA2(21), A2 => n7376, B1 => n7375, B2 => 
                           n7356, ZN => N2538);
   U1760 : AOI22_X1 port map( A1 => DATA2(20), A2 => n7376, B1 => n7375, B2 => 
                           n7357, ZN => N2537);
   U1761 : AOI22_X1 port map( A1 => DATA2(19), A2 => n7371, B1 => n7370, B2 => 
                           n7358, ZN => N2536);
   U1762 : AOI22_X1 port map( A1 => DATA2(18), A2 => n7371, B1 => n7370, B2 => 
                           n7359, ZN => N2535);
   U1763 : INV_X1 port map( A => DATA2(17), ZN => n7360);
   U1764 : AOI22_X1 port map( A1 => DATA2(17), A2 => n7371, B1 => n7370, B2 => 
                           n7360, ZN => N2534);
   U1765 : AOI22_X1 port map( A1 => DATA2(16), A2 => n7371, B1 => n7370, B2 => 
                           n7361, ZN => N2533);
   U1766 : INV_X1 port map( A => DATA2(15), ZN => n7362);
   U1767 : AOI22_X1 port map( A1 => DATA2(15), A2 => n7371, B1 => n7370, B2 => 
                           n7362, ZN => N2532);
   U1768 : AOI22_X1 port map( A1 => DATA2(14), A2 => n7371, B1 => n7370, B2 => 
                           n7363, ZN => N2531);
   U1769 : AOI22_X1 port map( A1 => DATA2(13), A2 => n7371, B1 => n7370, B2 => 
                           n7364, ZN => N2530);
   U1770 : AOI22_X1 port map( A1 => DATA2(12), A2 => n7371, B1 => n7370, B2 => 
                           n7365, ZN => N2529);
   U1771 : AOI22_X1 port map( A1 => DATA2(11), A2 => n7371, B1 => n7370, B2 => 
                           n7366, ZN => N2528);
   U1772 : AOI22_X1 port map( A1 => DATA2(10), A2 => n7371, B1 => n7370, B2 => 
                           n7367, ZN => N2527);
   U1773 : INV_X1 port map( A => DATA2(9), ZN => n7368);
   U1774 : AOI22_X1 port map( A1 => DATA2(9), A2 => n7371, B1 => n7370, B2 => 
                           n7368, ZN => N2526);
   U1775 : AOI22_X1 port map( A1 => DATA2(8), A2 => n7371, B1 => n7370, B2 => 
                           n7369, ZN => N2525);
   U1776 : AOI22_X1 port map( A1 => DATA2(7), A2 => n7376, B1 => n7375, B2 => 
                           n1946, ZN => N2524);
   U1777 : AOI22_X1 port map( A1 => DATA2(6), A2 => n7376, B1 => n7375, B2 => 
                           n7372, ZN => N2523);
   U1778 : AOI22_X1 port map( A1 => DATA2(5), A2 => n7376, B1 => n7375, B2 => 
                           n7373, ZN => N2522);
   U1779 : AOI22_X1 port map( A1 => DATA2(4), A2 => n7376, B1 => n7375, B2 => 
                           n7675, ZN => N2521);
   U1780 : AOI22_X1 port map( A1 => DATA2(3), A2 => n7376, B1 => n7375, B2 => 
                           n7661, ZN => N2520);
   U1781 : AOI22_X1 port map( A1 => DATA2(2), A2 => n7376, B1 => n7375, B2 => 
                           n1970, ZN => N2519);
   U1782 : AOI22_X1 port map( A1 => DATA2(1), A2 => n7376, B1 => n7375, B2 => 
                           n7374, ZN => N2518);
   U1783 : AOI22_X1 port map( A1 => DATA2(0), A2 => n7376, B1 => n7375, B2 => 
                           n7658, ZN => N2517);
   U1784 : NOR2_X1 port map( A1 => n7377, A2 => n1894, ZN => dataout_mul_0_port
                           );
   U1785 : INV_X1 port map( A => boothmul_pipelined_i_multiplicand_pip_2_3_port
                           , ZN => n7378);
   U1786 : NAND2_X1 port map( A1 => n7380, A2 => n7378, ZN => n7412);
   U1787 : NAND2_X1 port map( A1 => n7413, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, ZN 
                           => n7408);
   U1788 : INV_X1 port map( A => n7408, ZN => n7415);
   U1789 : NAND2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, 
                           ZN => n7379);
   U1790 : NOR2_X1 port map( A1 => n7415, A2 => n7410, ZN => n7381);
   U1791 : NAND2_X1 port map( A1 => n7380, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, ZN 
                           => n7417);
   U1792 : OAI222_X1 port map( A1 => n1893, A2 => n7412, B1 => n1894, B2 => 
                           n7381, C1 => n1892, C2 => n7417, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1793 : OAI22_X1 port map( A1 => n1890, A2 => n7417, B1 => n1892, B2 => 
                           n7408, ZN => n7382);
   U1794 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, A => n7382,
                           ZN => n7383);
   U1795 : OAI21_X1 port map( B1 => n1891, B2 => n7412, A => n7383, ZN => 
                           boothmul_pipelined_i_mux_out_1_4_port);
   U1796 : OAI22_X1 port map( A1 => n1890, A2 => n7408, B1 => n7417, B2 => 
                           n1888, ZN => n7384);
   U1797 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_4_63_port, B2
                           => n7410, A => n7384, ZN => n7385);
   U1798 : OAI21_X1 port map( B1 => n7412, B2 => n1889, A => n7385, ZN => 
                           boothmul_pipelined_i_mux_out_1_5_port);
   U1799 : OAI22_X1 port map( A1 => n7417, A2 => n1886, B1 => n7408, B2 => 
                           n1888, ZN => n7386);
   U1800 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, A => n7386,
                           ZN => n7387);
   U1801 : OAI21_X1 port map( B1 => n7412, B2 => n1887, A => n7387, ZN => 
                           boothmul_pipelined_i_mux_out_1_6_port);
   U1802 : OAI22_X1 port map( A1 => n7417, A2 => n1884, B1 => n7408, B2 => 
                           n1886, ZN => n7388);
   U1803 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, A => n7388,
                           ZN => n7389);
   U1804 : OAI21_X1 port map( B1 => n7412, B2 => n1885, A => n7389, ZN => 
                           boothmul_pipelined_i_mux_out_1_7_port);
   U1805 : OAI22_X1 port map( A1 => n7417, A2 => n1882, B1 => n7408, B2 => 
                           n1884, ZN => n7390);
   U1806 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, A => n7390,
                           ZN => n7391);
   U1807 : OAI21_X1 port map( B1 => n7412, B2 => n1883, A => n7391, ZN => 
                           boothmul_pipelined_i_mux_out_1_8_port);
   U1808 : OAI22_X1 port map( A1 => n7417, A2 => n1880, B1 => n7408, B2 => 
                           n1882, ZN => n7392);
   U1809 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, A => n7392,
                           ZN => n7393);
   U1810 : OAI21_X1 port map( B1 => n7412, B2 => n1881, A => n7393, ZN => 
                           boothmul_pipelined_i_mux_out_1_9_port);
   U1811 : OAI22_X1 port map( A1 => n7417, A2 => n1878, B1 => n7408, B2 => 
                           n1880, ZN => n7394);
   U1812 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_34_port, A => n7394,
                           ZN => n7395);
   U1813 : OAI21_X1 port map( B1 => n7412, B2 => n1879, A => n7395, ZN => 
                           boothmul_pipelined_i_mux_out_1_10_port);
   U1814 : OAI22_X1 port map( A1 => n7417, A2 => n1876, B1 => n7408, B2 => 
                           n1878, ZN => n7396);
   U1815 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_33_port, A => n7396,
                           ZN => n7397);
   U1816 : OAI21_X1 port map( B1 => n7412, B2 => n1877, A => n7397, ZN => 
                           boothmul_pipelined_i_mux_out_1_11_port);
   U1817 : OAI22_X1 port map( A1 => n7417, A2 => n1874, B1 => n7408, B2 => 
                           n1876, ZN => n7398);
   U1818 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_32_port, A => n7398,
                           ZN => n7399);
   U1819 : OAI21_X1 port map( B1 => n7412, B2 => n1875, A => n7399, ZN => 
                           boothmul_pipelined_i_mux_out_1_12_port);
   U1820 : OAI22_X1 port map( A1 => n7417, A2 => n1872, B1 => n7408, B2 => 
                           n1874, ZN => n7400);
   U1821 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_31_port, A => n7400,
                           ZN => n7401);
   U1822 : OAI21_X1 port map( B1 => n7412, B2 => n1873, A => n7401, ZN => 
                           boothmul_pipelined_i_mux_out_1_13_port);
   U1823 : OAI22_X1 port map( A1 => n7417, A2 => n1870, B1 => n7408, B2 => 
                           n1872, ZN => n7402);
   U1824 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_30_port, A => n7402,
                           ZN => n7403);
   U1825 : OAI21_X1 port map( B1 => n7412, B2 => n1871, A => n7403, ZN => 
                           boothmul_pipelined_i_mux_out_1_14_port);
   U1826 : OAI22_X1 port map( A1 => n7417, A2 => n1868, B1 => n7408, B2 => 
                           n1870, ZN => n7404);
   U1827 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_29_port, A => n7404,
                           ZN => n7405);
   U1828 : OAI21_X1 port map( B1 => n7412, B2 => n1869, A => n7405, ZN => 
                           boothmul_pipelined_i_mux_out_1_15_port);
   U1829 : OAI22_X1 port map( A1 => n7417, A2 => n1866, B1 => n7408, B2 => 
                           n1868, ZN => n7406);
   U1830 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_28_port, A => n7406,
                           ZN => n7407);
   U1831 : OAI21_X1 port map( B1 => n7412, B2 => n1867, A => n7407, ZN => 
                           boothmul_pipelined_i_mux_out_1_16_port);
   U1832 : OAI22_X1 port map( A1 => n7417, A2 => n1864, B1 => n7408, B2 => 
                           n1866, ZN => n7409);
   U1833 : AOI21_X1 port map( B1 => n7410, B2 => 
                           boothmul_pipelined_i_muxes_in_4_27_port, A => n7409,
                           ZN => n7411);
   U1834 : OAI21_X1 port map( B1 => n7412, B2 => n1865, A => n7411, ZN => 
                           boothmul_pipelined_i_mux_out_1_17_port);
   U1835 : XNOR2_X1 port map( A => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, B 
                           => n1865, ZN => n1863);
   U1836 : NOR3_X1 port map( A1 => n7413, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A3 
                           => n1865, ZN => n7414);
   U1837 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           B2 => n7415, A => n7414, ZN => n7416);
   U1838 : OAI21_X1 port map( B1 => n1863, B2 => n7417, A => n7416, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1839 : OR2_X1 port map( A1 => n7418, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n2806);
   U1840 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n4292, B1 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B2 => n3933
                           , ZN => n7419);
   U1841 : OAI221_X1 port map( B1 => n1894, B2 => n4191, C1 => n1894, C2 => 
                           n4055, A => n7419, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1842 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B2 => n3933
                           , ZN => n7421);
   U1843 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n4292, ZN => n7420);
   U1844 : OAI211_X1 port map( C1 => n4055, C2 => n1893, A => n7421, B => n7420
                           , ZN => boothmul_pipelined_i_mux_out_2_6_port);
   U1845 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_62_port, A2
                           => n3933, B1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B2 => 
                           n4292, ZN => n7423);
   U1846 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n4399, ZN => n7422);
   U1847 : OAI211_X1 port map( C1 => n4055, C2 => n1891, A => n7423, B => n7422
                           , ZN => boothmul_pipelined_i_mux_out_2_7_port);
   U1848 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B2 => 
                           n4292, ZN => n7425);
   U1849 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_61_port, A2
                           => n3933, ZN => n7424);
   U1850 : OAI211_X1 port map( C1 => n4055, C2 => n1889, A => n7425, B => n7424
                           , ZN => boothmul_pipelined_i_mux_out_2_8_port);
   U1851 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B2 => 
                           n4292, ZN => n7427);
   U1852 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_60_port, A2
                           => n3933, ZN => n7426);
   U1853 : OAI211_X1 port map( C1 => n4055, C2 => n1887, A => n7427, B => n7426
                           , ZN => boothmul_pipelined_i_mux_out_2_9_port);
   U1854 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B2 => 
                           n4292, ZN => n7429);
   U1855 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_59_port, A2
                           => n3933, ZN => n7428);
   U1856 : OAI211_X1 port map( C1 => n4055, C2 => n1885, A => n7429, B => n7428
                           , ZN => boothmul_pipelined_i_mux_out_2_10_port);
   U1857 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B2 => 
                           n4292, ZN => n7431);
   U1858 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_34_port, A2
                           => n3933, ZN => n7430);
   U1859 : OAI211_X1 port map( C1 => n4055, C2 => n1883, A => n7431, B => n7430
                           , ZN => boothmul_pipelined_i_mux_out_2_11_port);
   U1860 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B2 => 
                           n4292, ZN => n7433);
   U1861 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_33_port, A2
                           => n3933, ZN => n7432);
   U1862 : OAI211_X1 port map( C1 => n4055, C2 => n1881, A => n7433, B => n7432
                           , ZN => boothmul_pipelined_i_mux_out_2_12_port);
   U1863 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B2 => 
                           n4292, ZN => n7435);
   U1864 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_32_port, A2
                           => n3933, ZN => n7434);
   U1865 : OAI211_X1 port map( C1 => n4055, C2 => n1879, A => n7435, B => n7434
                           , ZN => boothmul_pipelined_i_mux_out_2_13_port);
   U1866 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B2 => 
                           n4292, ZN => n7437);
   U1867 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_31_port, A2
                           => n3933, ZN => n7436);
   U1868 : OAI211_X1 port map( C1 => n4055, C2 => n1877, A => n7437, B => n7436
                           , ZN => boothmul_pipelined_i_mux_out_2_14_port);
   U1869 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B2 => 
                           n4292, ZN => n7439);
   U1870 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_30_port, A2
                           => n3933, ZN => n7438);
   U1871 : OAI211_X1 port map( C1 => n4055, C2 => n1875, A => n7439, B => n7438
                           , ZN => boothmul_pipelined_i_mux_out_2_15_port);
   U1872 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B2 => 
                           n4292, ZN => n7441);
   U1873 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_29_port, A2
                           => n3933, ZN => n7440);
   U1874 : OAI211_X1 port map( C1 => n4055, C2 => n1873, A => n7441, B => n7440
                           , ZN => boothmul_pipelined_i_mux_out_2_16_port);
   U1875 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B2 => 
                           n4292, ZN => n7443);
   U1876 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_28_port, A2
                           => n3933, ZN => n7442);
   U1877 : OAI211_X1 port map( C1 => n4055, C2 => n1871, A => n7443, B => n7442
                           , ZN => boothmul_pipelined_i_mux_out_2_17_port);
   U1878 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B2 => 
                           n4292, ZN => n7445);
   U1879 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_27_port, A2
                           => n3933, ZN => n7444);
   U1880 : OAI211_X1 port map( C1 => n4055, C2 => n1869, A => n7445, B => n7444
                           , ZN => boothmul_pipelined_i_mux_out_2_18_port);
   U1881 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n4399, B1 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B2 => 
                           n4292, ZN => n7447);
   U1882 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n3933, ZN => n7446
                           );
   U1883 : OAI211_X1 port map( C1 => n4055, C2 => n1867, A => n7447, B => n7446
                           , ZN => boothmul_pipelined_i_mux_out_2_19_port);
   U1884 : OAI222_X1 port map( A1 => n1864, A2 => n4191, B1 => n1865, B2 => 
                           n4054, C1 => n4398, C2 => n1863, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U1885 : NAND3_X1 port map( A1 => n6005, A2 => n4294, A3 => n4295, ZN => 
                           n7481);
   U1886 : NOR2_X1 port map( A1 => n4294, A2 => n4295, ZN => n7448);
   U1887 : NAND2_X1 port map( A1 => n7448, A2 => n7769, ZN => n7485);
   U1888 : NOR2_X1 port map( A1 => n7769, A2 => n7449, ZN => n7451);
   U1889 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n7480, B1 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B2 => n7451
                           , ZN => n7450);
   U1890 : OAI221_X1 port map( B1 => n1894, B2 => n7481, C1 => n1894, C2 => 
                           n7485, A => n7450, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1891 : INV_X1 port map( A => n7451, ZN => n7482);
   U1892 : OAI22_X1 port map( A1 => n1892, A2 => n7485, B1 => n1893, B2 => 
                           n7481, ZN => n7452);
   U1893 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           B2 => n7480, A => n7452, ZN => n7453);
   U1894 : OAI21_X1 port map( B1 => n1891, B2 => n7482, A => n7453, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1895 : OAI22_X1 port map( A1 => n1890, A2 => n7485, B1 => n1891, B2 => 
                           n7481, ZN => n7454);
   U1896 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           B2 => n7480, A => n7454, ZN => n7455);
   U1897 : OAI21_X1 port map( B1 => n1889, B2 => n7482, A => n7455, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1898 : OAI22_X1 port map( A1 => n1889, A2 => n7481, B1 => n1888, B2 => 
                           n7485, ZN => n7456);
   U1899 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           B2 => n7480, A => n7456, ZN => n7457);
   U1900 : OAI21_X1 port map( B1 => n1887, B2 => n7482, A => n7457, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1901 : OAI22_X1 port map( A1 => n1887, A2 => n7481, B1 => n1886, B2 => 
                           n7485, ZN => n7458);
   U1902 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           B2 => n7480, A => n7458, ZN => n7459);
   U1903 : OAI21_X1 port map( B1 => n1885, B2 => n7482, A => n7459, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1904 : OAI22_X1 port map( A1 => n1885, A2 => n7481, B1 => n1884, B2 => 
                           n7485, ZN => n7460);
   U1905 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           B2 => n7480, A => n7460, ZN => n7461);
   U1906 : OAI21_X1 port map( B1 => n1883, B2 => n7482, A => n7461, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1907 : OAI22_X1 port map( A1 => n1883, A2 => n7481, B1 => n1882, B2 => 
                           n7485, ZN => n7462);
   U1908 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           B2 => n7480, A => n7462, ZN => n7463);
   U1909 : OAI21_X1 port map( B1 => n1881, B2 => n7482, A => n7463, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U1910 : OAI22_X1 port map( A1 => n1881, A2 => n7481, B1 => n1880, B2 => 
                           n7485, ZN => n7464);
   U1911 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           B2 => n7480, A => n7464, ZN => n7465);
   U1912 : OAI21_X1 port map( B1 => n1879, B2 => n7482, A => n7465, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U1913 : OAI22_X1 port map( A1 => n1879, A2 => n7481, B1 => n1878, B2 => 
                           n7485, ZN => n7466);
   U1914 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           B2 => n7480, A => n7466, ZN => n7467);
   U1915 : OAI21_X1 port map( B1 => n1877, B2 => n7482, A => n7467, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U1916 : OAI22_X1 port map( A1 => n1877, A2 => n7481, B1 => n1876, B2 => 
                           n7485, ZN => n7468);
   U1917 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           B2 => n7480, A => n7468, ZN => n7469);
   U1918 : OAI21_X1 port map( B1 => n1875, B2 => n7482, A => n7469, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U1919 : OAI22_X1 port map( A1 => n1875, A2 => n7481, B1 => n1874, B2 => 
                           n7485, ZN => n7470);
   U1920 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           B2 => n7480, A => n7470, ZN => n7471);
   U1921 : OAI21_X1 port map( B1 => n1873, B2 => n7482, A => n7471, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U1922 : OAI22_X1 port map( A1 => n1873, A2 => n7481, B1 => n1872, B2 => 
                           n7485, ZN => n7472);
   U1923 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           B2 => n7480, A => n7472, ZN => n7473);
   U1924 : OAI21_X1 port map( B1 => n1871, B2 => n7482, A => n7473, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U1925 : OAI22_X1 port map( A1 => n1871, A2 => n7481, B1 => n1870, B2 => 
                           n7485, ZN => n7474);
   U1926 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           B2 => n7480, A => n7474, ZN => n7475);
   U1927 : OAI21_X1 port map( B1 => n1869, B2 => n7482, A => n7475, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U1928 : OAI22_X1 port map( A1 => n1869, A2 => n7481, B1 => n1868, B2 => 
                           n7485, ZN => n7476);
   U1929 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           B2 => n7480, A => n7476, ZN => n7477);
   U1930 : OAI21_X1 port map( B1 => n1867, B2 => n7482, A => n7477, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U1931 : OAI22_X1 port map( A1 => n1867, A2 => n7481, B1 => n1866, B2 => 
                           n7485, ZN => n7478);
   U1932 : AOI21_X1 port map( B1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           B2 => n7480, A => n7478, ZN => n7479);
   U1933 : OAI21_X1 port map( B1 => n1865, B2 => n7482, A => n7479, ZN => 
                           boothmul_pipelined_i_mux_out_3_21_port);
   U1934 : INV_X1 port map( A => n7480, ZN => n7484);
   U1935 : AND2_X1 port map( A1 => n7482, A2 => n7481, ZN => n7483);
   U1936 : OAI222_X1 port map( A1 => n7485, A2 => n1864, B1 => n7484, B2 => 
                           n1863, C1 => n1865, C2 => n7483, ZN => 
                           boothmul_pipelined_i_mux_out_3_22_port);
   U1937 : NAND3_X1 port map( A1 => n6009, A2 => n4296, A3 => n4298, ZN => 
                           n7524);
   U1938 : OR2_X1 port map( A1 => n4296, A2 => n4298, ZN => n7486);
   U1939 : INV_X1 port map( A => n7522, ZN => n7490);
   U1940 : NAND2_X1 port map( A1 => n6009, A2 => n7487, ZN => n7525);
   U1941 : INV_X1 port map( A => n7525, ZN => n7518);
   U1942 : AOI22_X1 port map( A1 => n7518, A2 => n4336, B1 => n7521, B2 => 
                           n4174, ZN => n7489);
   U1943 : OAI221_X1 port map( B1 => n7743, B2 => n7524, C1 => n7743, C2 => 
                           n7490, A => n7489, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U1944 : INV_X1 port map( A => n7524, ZN => n7517);
   U1945 : AOI22_X1 port map( A1 => n4336, A2 => n7517, B1 => n7522, B2 => 
                           n4174, ZN => n7492);
   U1946 : AOI22_X1 port map( A1 => n7518, A2 => n4340, B1 => n7521, B2 => 
                           n4170, ZN => n7491);
   U1947 : NAND2_X1 port map( A1 => n7492, A2 => n7491, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U1948 : AOI22_X1 port map( A1 => n7517, A2 => n4340, B1 => n7522, B2 => 
                           n4170, ZN => n7494);
   U1949 : AOI22_X1 port map( A1 => n7518, A2 => n4344, B1 => n7521, B2 => 
                           n4166, ZN => n7493);
   U1950 : NAND2_X1 port map( A1 => n7494, A2 => n7493, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U1951 : AOI22_X1 port map( A1 => n7517, A2 => n4344, B1 => n7522, B2 => 
                           n4166, ZN => n7496);
   U1952 : AOI22_X1 port map( A1 => n7518, A2 => n4348, B1 => n7521, B2 => 
                           n4162, ZN => n7495);
   U1953 : NAND2_X1 port map( A1 => n7496, A2 => n7495, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U1954 : AOI22_X1 port map( A1 => n7517, A2 => n4348, B1 => n7522, B2 => 
                           n4162, ZN => n7498);
   U1955 : AOI22_X1 port map( A1 => n7518, A2 => n4352, B1 => n7521, B2 => 
                           n4158, ZN => n7497);
   U1956 : NAND2_X1 port map( A1 => n7498, A2 => n7497, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U1957 : AOI22_X1 port map( A1 => n7517, A2 => n4352, B1 => n7522, B2 => 
                           n4158, ZN => n7500);
   U1958 : AOI22_X1 port map( A1 => n7518, A2 => n4356, B1 => n7521, B2 => 
                           n4154, ZN => n7499);
   U1959 : NAND2_X1 port map( A1 => n7500, A2 => n7499, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U1960 : AOI22_X1 port map( A1 => n7517, A2 => n4356, B1 => n7522, B2 => 
                           n4154, ZN => n7502);
   U1961 : AOI22_X1 port map( A1 => n7518, A2 => n4360, B1 => n7521, B2 => 
                           n4150, ZN => n7501);
   U1962 : NAND2_X1 port map( A1 => n7502, A2 => n7501, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U1963 : AOI22_X1 port map( A1 => n7517, A2 => n4360, B1 => n7522, B2 => 
                           n4150, ZN => n7504);
   U1964 : AOI22_X1 port map( A1 => n7518, A2 => n4364, B1 => n7521, B2 => 
                           n4146, ZN => n7503);
   U1965 : NAND2_X1 port map( A1 => n7504, A2 => n7503, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U1966 : AOI22_X1 port map( A1 => n7517, A2 => n4364, B1 => n7522, B2 => 
                           n4146, ZN => n7506);
   U1967 : AOI22_X1 port map( A1 => n7518, A2 => n4368, B1 => n7521, B2 => 
                           n4142, ZN => n7505);
   U1968 : NAND2_X1 port map( A1 => n7506, A2 => n7505, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U1969 : AOI22_X1 port map( A1 => n7517, A2 => n4368, B1 => n7522, B2 => 
                           n4142, ZN => n7508);
   U1970 : AOI22_X1 port map( A1 => n7518, A2 => n4372, B1 => n7521, B2 => 
                           n4138, ZN => n7507);
   U1971 : NAND2_X1 port map( A1 => n7508, A2 => n7507, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U1972 : AOI22_X1 port map( A1 => n7517, A2 => n4372, B1 => n7522, B2 => 
                           n4138, ZN => n7510);
   U1973 : AOI22_X1 port map( A1 => n7518, A2 => n4376, B1 => n7521, B2 => 
                           n4134, ZN => n7509);
   U1974 : NAND2_X1 port map( A1 => n7510, A2 => n7509, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U1975 : AOI22_X1 port map( A1 => n7517, A2 => n4376, B1 => n7522, B2 => 
                           n4134, ZN => n7512);
   U1976 : AOI22_X1 port map( A1 => n7518, A2 => n4380, B1 => n7521, B2 => 
                           n4130, ZN => n7511);
   U1977 : NAND2_X1 port map( A1 => n7512, A2 => n7511, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U1978 : AOI22_X1 port map( A1 => n7517, A2 => n4380, B1 => n7522, B2 => 
                           n4130, ZN => n7514);
   U1979 : AOI22_X1 port map( A1 => n7518, A2 => n4384, B1 => n7521, B2 => 
                           n4126, ZN => n7513);
   U1980 : NAND2_X1 port map( A1 => n7514, A2 => n7513, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U1981 : AOI22_X1 port map( A1 => n7517, A2 => n4384, B1 => n7522, B2 => 
                           n4126, ZN => n7516);
   U1982 : AOI22_X1 port map( A1 => n7518, A2 => n4388, B1 => n7521, B2 => 
                           n4122, ZN => n7515);
   U1983 : NAND2_X1 port map( A1 => n7516, A2 => n7515, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U1984 : AOI22_X1 port map( A1 => n7517, A2 => n4388, B1 => n7522, B2 => 
                           n4122, ZN => n7520);
   U1985 : AOI22_X1 port map( A1 => n7518, A2 => n4392, B1 => n7521, B2 => 
                           n4118, ZN => n7519);
   U1986 : NAND2_X1 port map( A1 => n7520, A2 => n7519, ZN => 
                           boothmul_pipelined_i_mux_out_4_23_port);
   U1987 : AOI22_X1 port map( A1 => n7522, A2 => n4118, B1 => n7521, B2 => 
                           n4288, ZN => n7523);
   U1988 : OAI221_X1 port map( B1 => n7809, B2 => n7525, C1 => n7809, C2 => 
                           n7524, A => n7523, ZN => 
                           boothmul_pipelined_i_mux_out_4_24_port);
   U1989 : NAND3_X1 port map( A1 => n6008, A2 => n4300, A3 => n4303, ZN => 
                           n7564);
   U1990 : OR2_X1 port map( A1 => n4300, A2 => n4303, ZN => n7526);
   U1991 : INV_X1 port map( A => n7562, ZN => n7530);
   U1992 : NAND2_X1 port map( A1 => n6008, A2 => n7527, ZN => n7565);
   U1993 : INV_X1 port map( A => n7565, ZN => n7558);
   U1994 : AOI22_X1 port map( A1 => n7558, A2 => n4335, B1 => n7561, B2 => 
                           n4173, ZN => n7529);
   U1995 : OAI221_X1 port map( B1 => n7744, B2 => n7564, C1 => n7744, C2 => 
                           n7530, A => n7529, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U1996 : INV_X1 port map( A => n7564, ZN => n7557);
   U1997 : AOI22_X1 port map( A1 => n4335, A2 => n7557, B1 => n7562, B2 => 
                           n4173, ZN => n7532);
   U1998 : AOI22_X1 port map( A1 => n7558, A2 => n4339, B1 => n7561, B2 => 
                           n4169, ZN => n7531);
   U1999 : NAND2_X1 port map( A1 => n7532, A2 => n7531, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2000 : AOI22_X1 port map( A1 => n7557, A2 => n4339, B1 => n7562, B2 => 
                           n4169, ZN => n7534);
   U2001 : AOI22_X1 port map( A1 => n7558, A2 => n4343, B1 => n7561, B2 => 
                           n4165, ZN => n7533);
   U2002 : NAND2_X1 port map( A1 => n7534, A2 => n7533, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2003 : AOI22_X1 port map( A1 => n7557, A2 => n4343, B1 => n7562, B2 => 
                           n4165, ZN => n7536);
   U2004 : AOI22_X1 port map( A1 => n7558, A2 => n4347, B1 => n7561, B2 => 
                           n4161, ZN => n7535);
   U2005 : NAND2_X1 port map( A1 => n7536, A2 => n7535, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2006 : AOI22_X1 port map( A1 => n7557, A2 => n4347, B1 => n7562, B2 => 
                           n4161, ZN => n7538);
   U2007 : AOI22_X1 port map( A1 => n7558, A2 => n4351, B1 => n7561, B2 => 
                           n4157, ZN => n7537);
   U2008 : NAND2_X1 port map( A1 => n7538, A2 => n7537, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2009 : AOI22_X1 port map( A1 => n7557, A2 => n4351, B1 => n7562, B2 => 
                           n4157, ZN => n7540);
   U2010 : AOI22_X1 port map( A1 => n7558, A2 => n4355, B1 => n7561, B2 => 
                           n4153, ZN => n7539);
   U2011 : NAND2_X1 port map( A1 => n7540, A2 => n7539, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2012 : AOI22_X1 port map( A1 => n7557, A2 => n4355, B1 => n7562, B2 => 
                           n4153, ZN => n7542);
   U2013 : AOI22_X1 port map( A1 => n7558, A2 => n4359, B1 => n7561, B2 => 
                           n4149, ZN => n7541);
   U2014 : NAND2_X1 port map( A1 => n7542, A2 => n7541, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2015 : AOI22_X1 port map( A1 => n7557, A2 => n4359, B1 => n7562, B2 => 
                           n4149, ZN => n7544);
   U2016 : AOI22_X1 port map( A1 => n7558, A2 => n4363, B1 => n7561, B2 => 
                           n4145, ZN => n7543);
   U2017 : NAND2_X1 port map( A1 => n7544, A2 => n7543, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2018 : AOI22_X1 port map( A1 => n7557, A2 => n4363, B1 => n7562, B2 => 
                           n4145, ZN => n7546);
   U2019 : AOI22_X1 port map( A1 => n7558, A2 => n4367, B1 => n7561, B2 => 
                           n4141, ZN => n7545);
   U2020 : NAND2_X1 port map( A1 => n7546, A2 => n7545, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2021 : AOI22_X1 port map( A1 => n7557, A2 => n4367, B1 => n7562, B2 => 
                           n4141, ZN => n7548);
   U2022 : AOI22_X1 port map( A1 => n7558, A2 => n4371, B1 => n7561, B2 => 
                           n4137, ZN => n7547);
   U2023 : NAND2_X1 port map( A1 => n7548, A2 => n7547, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2024 : AOI22_X1 port map( A1 => n7557, A2 => n4371, B1 => n7562, B2 => 
                           n4137, ZN => n7550);
   U2025 : AOI22_X1 port map( A1 => n7558, A2 => n4375, B1 => n7561, B2 => 
                           n4133, ZN => n7549);
   U2026 : NAND2_X1 port map( A1 => n7550, A2 => n7549, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2027 : AOI22_X1 port map( A1 => n7557, A2 => n4375, B1 => n7562, B2 => 
                           n4133, ZN => n7552);
   U2028 : AOI22_X1 port map( A1 => n7558, A2 => n4379, B1 => n7561, B2 => 
                           n4129, ZN => n7551);
   U2029 : NAND2_X1 port map( A1 => n7552, A2 => n7551, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2030 : AOI22_X1 port map( A1 => n7557, A2 => n4379, B1 => n7562, B2 => 
                           n4129, ZN => n7554);
   U2031 : AOI22_X1 port map( A1 => n7558, A2 => n4383, B1 => n7561, B2 => 
                           n4125, ZN => n7553);
   U2032 : NAND2_X1 port map( A1 => n7554, A2 => n7553, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2033 : AOI22_X1 port map( A1 => n7557, A2 => n4383, B1 => n7562, B2 => 
                           n4125, ZN => n7556);
   U2034 : AOI22_X1 port map( A1 => n7558, A2 => n4387, B1 => n7561, B2 => 
                           n4121, ZN => n7555);
   U2035 : NAND2_X1 port map( A1 => n7556, A2 => n7555, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2036 : AOI22_X1 port map( A1 => n7557, A2 => n4387, B1 => n7562, B2 => 
                           n4121, ZN => n7560);
   U2037 : AOI22_X1 port map( A1 => n7558, A2 => n4391, B1 => n7561, B2 => 
                           n4117, ZN => n7559);
   U2038 : NAND2_X1 port map( A1 => n7560, A2 => n7559, ZN => 
                           boothmul_pipelined_i_mux_out_5_25_port);
   U2039 : AOI22_X1 port map( A1 => n7562, A2 => n4117, B1 => n7561, B2 => 
                           n4287, ZN => n7563);
   U2040 : OAI221_X1 port map( B1 => n7811, B2 => n7565, C1 => n7811, C2 => 
                           n7564, A => n7563, ZN => 
                           boothmul_pipelined_i_mux_out_5_26_port);
   U2041 : NAND3_X1 port map( A1 => n6006, A2 => n4306, A3 => n4310, ZN => 
                           n7604);
   U2042 : OR2_X1 port map( A1 => n4306, A2 => n4310, ZN => n7566);
   U2043 : INV_X1 port map( A => n7602, ZN => n7570);
   U2044 : NAND2_X1 port map( A1 => n6006, A2 => n7567, ZN => n7605);
   U2045 : INV_X1 port map( A => n7605, ZN => n7598);
   U2046 : AOI22_X1 port map( A1 => n7598, A2 => n4334, B1 => n7601, B2 => 
                           n4172, ZN => n7569);
   U2047 : OAI221_X1 port map( B1 => n7745, B2 => n7604, C1 => n7745, C2 => 
                           n7570, A => n7569, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2048 : INV_X1 port map( A => n7604, ZN => n7597);
   U2049 : AOI22_X1 port map( A1 => n4334, A2 => n7597, B1 => n7602, B2 => 
                           n4172, ZN => n7572);
   U2050 : AOI22_X1 port map( A1 => n7598, A2 => n4338, B1 => n7601, B2 => 
                           n4168, ZN => n7571);
   U2051 : NAND2_X1 port map( A1 => n7572, A2 => n7571, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2052 : AOI22_X1 port map( A1 => n7597, A2 => n4338, B1 => n7602, B2 => 
                           n4168, ZN => n7574);
   U2053 : AOI22_X1 port map( A1 => n7598, A2 => n4342, B1 => n7601, B2 => 
                           n4164, ZN => n7573);
   U2054 : NAND2_X1 port map( A1 => n7574, A2 => n7573, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2055 : AOI22_X1 port map( A1 => n7597, A2 => n4342, B1 => n7602, B2 => 
                           n4164, ZN => n7576);
   U2056 : AOI22_X1 port map( A1 => n7598, A2 => n4346, B1 => n7601, B2 => 
                           n4160, ZN => n7575);
   U2057 : NAND2_X1 port map( A1 => n7576, A2 => n7575, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2058 : AOI22_X1 port map( A1 => n7597, A2 => n4346, B1 => n7602, B2 => 
                           n4160, ZN => n7578);
   U2059 : AOI22_X1 port map( A1 => n7598, A2 => n4350, B1 => n7601, B2 => 
                           n4156, ZN => n7577);
   U2060 : NAND2_X1 port map( A1 => n7578, A2 => n7577, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2061 : AOI22_X1 port map( A1 => n7597, A2 => n4350, B1 => n7602, B2 => 
                           n4156, ZN => n7580);
   U2062 : AOI22_X1 port map( A1 => n7598, A2 => n4354, B1 => n7601, B2 => 
                           n4152, ZN => n7579);
   U2063 : NAND2_X1 port map( A1 => n7580, A2 => n7579, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2064 : AOI22_X1 port map( A1 => n7597, A2 => n4354, B1 => n7602, B2 => 
                           n4152, ZN => n7582);
   U2065 : AOI22_X1 port map( A1 => n7598, A2 => n4358, B1 => n7601, B2 => 
                           n4148, ZN => n7581);
   U2066 : NAND2_X1 port map( A1 => n7582, A2 => n7581, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2067 : AOI22_X1 port map( A1 => n7597, A2 => n4358, B1 => n7602, B2 => 
                           n4148, ZN => n7584);
   U2068 : AOI22_X1 port map( A1 => n7598, A2 => n4362, B1 => n7601, B2 => 
                           n4144, ZN => n7583);
   U2069 : NAND2_X1 port map( A1 => n7584, A2 => n7583, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2070 : AOI22_X1 port map( A1 => n7597, A2 => n4362, B1 => n7602, B2 => 
                           n4144, ZN => n7586);
   U2071 : AOI22_X1 port map( A1 => n7598, A2 => n4366, B1 => n7601, B2 => 
                           n4140, ZN => n7585);
   U2072 : NAND2_X1 port map( A1 => n7586, A2 => n7585, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2073 : AOI22_X1 port map( A1 => n7597, A2 => n4366, B1 => n7602, B2 => 
                           n4140, ZN => n7588);
   U2074 : AOI22_X1 port map( A1 => n7598, A2 => n4370, B1 => n7601, B2 => 
                           n4136, ZN => n7587);
   U2075 : NAND2_X1 port map( A1 => n7588, A2 => n7587, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2076 : AOI22_X1 port map( A1 => n7597, A2 => n4370, B1 => n7602, B2 => 
                           n4136, ZN => n7590);
   U2077 : AOI22_X1 port map( A1 => n7598, A2 => n4374, B1 => n7601, B2 => 
                           n4132, ZN => n7589);
   U2078 : NAND2_X1 port map( A1 => n7590, A2 => n7589, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2079 : AOI22_X1 port map( A1 => n7597, A2 => n4374, B1 => n7602, B2 => 
                           n4132, ZN => n7592);
   U2080 : AOI22_X1 port map( A1 => n7598, A2 => n4378, B1 => n7601, B2 => 
                           n4128, ZN => n7591);
   U2081 : NAND2_X1 port map( A1 => n7592, A2 => n7591, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2082 : AOI22_X1 port map( A1 => n7597, A2 => n4378, B1 => n7602, B2 => 
                           n4128, ZN => n7594);
   U2083 : AOI22_X1 port map( A1 => n7598, A2 => n4382, B1 => n7601, B2 => 
                           n4124, ZN => n7593);
   U2084 : NAND2_X1 port map( A1 => n7594, A2 => n7593, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2085 : AOI22_X1 port map( A1 => n7597, A2 => n4382, B1 => n7602, B2 => 
                           n4124, ZN => n7596);
   U2086 : AOI22_X1 port map( A1 => n7598, A2 => n4386, B1 => n7601, B2 => 
                           n4120, ZN => n7595);
   U2087 : NAND2_X1 port map( A1 => n7596, A2 => n7595, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2088 : AOI22_X1 port map( A1 => n7597, A2 => n4386, B1 => n7602, B2 => 
                           n4120, ZN => n7600);
   U2089 : AOI22_X1 port map( A1 => n7598, A2 => n4390, B1 => n7601, B2 => 
                           n4116, ZN => n7599);
   U2090 : NAND2_X1 port map( A1 => n7600, A2 => n7599, ZN => 
                           boothmul_pipelined_i_mux_out_6_27_port);
   U2091 : AOI22_X1 port map( A1 => n7602, A2 => n4116, B1 => n7601, B2 => 
                           n4286, ZN => n7603);
   U2092 : OAI221_X1 port map( B1 => n7812, B2 => n7605, C1 => n7812, C2 => 
                           n7604, A => n7603, ZN => 
                           boothmul_pipelined_i_mux_out_6_28_port);
   U2093 : NAND3_X1 port map( A1 => n6007, A2 => n4319, A3 => n4314, ZN => 
                           n7610);
   U2094 : INV_X1 port map( A => n7642, ZN => n7609);
   U2095 : AND2_X1 port map( A1 => n6007, A2 => n7606, ZN => n7640);
   U2096 : AOI22_X1 port map( A1 => n7640, A2 => n4333, B1 => n7641, B2 => 
                           n4171, ZN => n7608);
   U2097 : OAI221_X1 port map( B1 => n7746, B2 => n7610, C1 => n7746, C2 => 
                           n7609, A => n7608, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2098 : INV_X1 port map( A => n7610, ZN => n7639);
   U2099 : AOI22_X1 port map( A1 => n4333, A2 => n7639, B1 => n7642, B2 => 
                           n4171, ZN => n7612);
   U2100 : AOI22_X1 port map( A1 => n7640, A2 => n4337, B1 => n7641, B2 => 
                           n4167, ZN => n7611);
   U2101 : NAND2_X1 port map( A1 => n7612, A2 => n7611, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2102 : AOI22_X1 port map( A1 => n7639, A2 => n4337, B1 => n7642, B2 => 
                           n4167, ZN => n7614);
   U2103 : AOI22_X1 port map( A1 => n7640, A2 => n4341, B1 => n7641, B2 => 
                           n4163, ZN => n7613);
   U2104 : NAND2_X1 port map( A1 => n7614, A2 => n7613, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2105 : AOI22_X1 port map( A1 => n7639, A2 => n4341, B1 => n7642, B2 => 
                           n4163, ZN => n7616);
   U2106 : AOI22_X1 port map( A1 => n7640, A2 => n4345, B1 => n7641, B2 => 
                           n4159, ZN => n7615);
   U2107 : NAND2_X1 port map( A1 => n7616, A2 => n7615, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2108 : AOI22_X1 port map( A1 => n7639, A2 => n4345, B1 => n7642, B2 => 
                           n4159, ZN => n7618);
   U2109 : AOI22_X1 port map( A1 => n7640, A2 => n4349, B1 => n7641, B2 => 
                           n4155, ZN => n7617);
   U2110 : NAND2_X1 port map( A1 => n7618, A2 => n7617, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2111 : AOI22_X1 port map( A1 => n7639, A2 => n4349, B1 => n7642, B2 => 
                           n4155, ZN => n7620);
   U2112 : AOI22_X1 port map( A1 => n7640, A2 => n4353, B1 => n7641, B2 => 
                           n4151, ZN => n7619);
   U2113 : NAND2_X1 port map( A1 => n7620, A2 => n7619, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2114 : AOI22_X1 port map( A1 => n7639, A2 => n4353, B1 => n7642, B2 => 
                           n4151, ZN => n7622);
   U2115 : AOI22_X1 port map( A1 => n7640, A2 => n4357, B1 => n7641, B2 => 
                           n4147, ZN => n7621);
   U2116 : NAND2_X1 port map( A1 => n7622, A2 => n7621, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2117 : AOI22_X1 port map( A1 => n7639, A2 => n4357, B1 => n7642, B2 => 
                           n4147, ZN => n7624);
   U2118 : AOI22_X1 port map( A1 => n7640, A2 => n4361, B1 => n7641, B2 => 
                           n4143, ZN => n7623);
   U2119 : NAND2_X1 port map( A1 => n7624, A2 => n7623, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2120 : AOI22_X1 port map( A1 => n7639, A2 => n4361, B1 => n7642, B2 => 
                           n4143, ZN => n7626);
   U2121 : AOI22_X1 port map( A1 => n7640, A2 => n4365, B1 => n7641, B2 => 
                           n4139, ZN => n7625);
   U2122 : NAND2_X1 port map( A1 => n7626, A2 => n7625, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2123 : AOI22_X1 port map( A1 => n7639, A2 => n4365, B1 => n7642, B2 => 
                           n4139, ZN => n7628);
   U2124 : AOI22_X1 port map( A1 => n7640, A2 => n4369, B1 => n7641, B2 => 
                           n4135, ZN => n7627);
   U2125 : NAND2_X1 port map( A1 => n7628, A2 => n7627, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2126 : AOI22_X1 port map( A1 => n7639, A2 => n4369, B1 => n7642, B2 => 
                           n4135, ZN => n7630);
   U2127 : AOI22_X1 port map( A1 => n7640, A2 => n4373, B1 => n7641, B2 => 
                           n4131, ZN => n7629);
   U2128 : NAND2_X1 port map( A1 => n7630, A2 => n7629, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2129 : AOI22_X1 port map( A1 => n7639, A2 => n4373, B1 => n7642, B2 => 
                           n4131, ZN => n7632);
   U2130 : AOI22_X1 port map( A1 => n7640, A2 => n4377, B1 => n7641, B2 => 
                           n4127, ZN => n7631);
   U2131 : NAND2_X1 port map( A1 => n7632, A2 => n7631, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2132 : AOI22_X1 port map( A1 => n7639, A2 => n4377, B1 => n7642, B2 => 
                           n4127, ZN => n7634);
   U2133 : AOI22_X1 port map( A1 => n7640, A2 => n4381, B1 => n7641, B2 => 
                           n4123, ZN => n7633);
   U2134 : NAND2_X1 port map( A1 => n7634, A2 => n7633, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2135 : AOI22_X1 port map( A1 => n7639, A2 => n4381, B1 => n7642, B2 => 
                           n4123, ZN => n7636);
   U2136 : AOI22_X1 port map( A1 => n7640, A2 => n4385, B1 => n7641, B2 => 
                           n4119, ZN => n7635);
   U2137 : NAND2_X1 port map( A1 => n7636, A2 => n7635, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2138 : AOI22_X1 port map( A1 => n7639, A2 => n4385, B1 => n7642, B2 => 
                           n4119, ZN => n7638);
   U2139 : AOI22_X1 port map( A1 => n7640, A2 => n4389, B1 => n7641, B2 => 
                           n4115, ZN => n7637);
   U2140 : NAND2_X1 port map( A1 => n7638, A2 => n7637, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2141 : OAI21_X1 port map( B1 => n7640, B2 => n7639, A => n4389, ZN => n7644
                           );
   U2142 : AOI22_X1 port map( A1 => n7642, A2 => n4115, B1 => n7641, B2 => 
                           n4285, ZN => n7643);
   U2143 : NAND2_X1 port map( A1 => n7644, A2 => n7643, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2144 : INV_X1 port map( A => n7649, ZN => n7648);
   U2145 : OAI222_X1 port map( A1 => n1894, A2 => n7645, B1 => n1892, B2 => 
                           n7652, C1 => n7648, C2 => n1893, ZN => 
                           dataout_mul_1_port);
   U2146 : OAI222_X1 port map( A1 => n1890, A2 => n7645, B1 => n1888, B2 => 
                           n7652, C1 => n1889, C2 => n7648, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_3_port);
   U2147 : OAI222_X1 port map( A1 => n1887, A2 => n7648, B1 => n1886, B2 => 
                           n7652, C1 => n1888, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_4_port);
   U2148 : OAI222_X1 port map( A1 => n1885, A2 => n7648, B1 => n1884, B2 => 
                           n7652, C1 => n1886, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_5_port);
   U2149 : OAI222_X1 port map( A1 => n1883, A2 => n7648, B1 => n1882, B2 => 
                           n7652, C1 => n1884, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_6_port);
   U2150 : OAI222_X1 port map( A1 => n1881, A2 => n7648, B1 => n1880, B2 => 
                           n7652, C1 => n1882, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_7_port);
   U2151 : OAI222_X1 port map( A1 => n1879, A2 => n7648, B1 => n1878, B2 => 
                           n7652, C1 => n1880, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_8_port);
   U2152 : OAI222_X1 port map( A1 => n1877, A2 => n7648, B1 => n1876, B2 => 
                           n7652, C1 => n1878, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_9_port);
   U2153 : OAI222_X1 port map( A1 => n1875, A2 => n7648, B1 => n1874, B2 => 
                           n7652, C1 => n1876, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_10_port);
   U2154 : OAI222_X1 port map( A1 => n1873, A2 => n7648, B1 => n1872, B2 => 
                           n7652, C1 => n1874, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_11_port);
   U2155 : OAI222_X1 port map( A1 => n1871, A2 => n7648, B1 => n1870, B2 => 
                           n7652, C1 => n1872, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_12_port);
   U2156 : OAI222_X1 port map( A1 => n1869, A2 => n7648, B1 => n1868, B2 => 
                           n7652, C1 => n1870, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_13_port);
   U2157 : OAI222_X1 port map( A1 => n1867, A2 => n7648, B1 => n1866, B2 => 
                           n7652, C1 => n1868, C2 => n7645, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_14_port);
   U2158 : AOI22_X1 port map( A1 => n7646, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n7650, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n7647);
   U2159 : OAI21_X1 port map( B1 => n7648, B2 => n1865, A => n7647, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2160 : AOI22_X1 port map( A1 => n7650, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n7649, B2 => data1_mul_15_port, ZN => n7651);
   U2161 : OAI21_X1 port map( B1 => n1863, B2 => n7652, A => n7651, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U2162 : NOR3_X1 port map( A1 => DATA2(2), A2 => n7656, A3 => n7674, ZN => 
                           n5985);
   U2163 : NOR2_X1 port map( A1 => n7658, A2 => n7653, ZN => n7655);
   U2164 : NOR2_X1 port map( A1 => n7654, A2 => n7655, ZN => n1966);
   U2165 : NAND2_X1 port map( A1 => n7655, A2 => n1967, ZN => n5986);
   U2166 : NOR2_X1 port map( A1 => n1219, A2 => n7656, ZN => n5987);
   U2167 : INV_X1 port map( A => n7657, ZN => n7673);
   U2168 : NOR3_X1 port map( A1 => DATA2(1), A2 => n7658, A3 => n7673, ZN => 
                           n5988);
   U2169 : NOR3_X1 port map( A1 => n7675, A2 => n7669, A3 => n7659, ZN => n5991
                           );
   U2170 : NOR2_X1 port map( A1 => n7660, A2 => n7667, ZN => n5994);
   U2171 : AOI21_X1 port map( B1 => n7662, B2 => n7661, A => n1959, ZN => n7668
                           );
   U2172 : INV_X1 port map( A => n1960, ZN => n7663);
   U2173 : NOR2_X1 port map( A1 => n7668, A2 => n7663, ZN => n5996);
   U2174 : NOR3_X1 port map( A1 => n1102, A2 => n7665, A3 => n7664, ZN => n5997
                           );
   U2175 : NOR2_X1 port map( A1 => n7666, A2 => n7673, ZN => n5998);
   U2176 : NAND3_X1 port map( A1 => DATA2(4), A2 => n7667, A3 => n7673, ZN => 
                           n5999);
   U2177 : NOR3_X1 port map( A1 => n1961, A2 => n7669, A3 => n7677, ZN => n6001
                           );
   U2178 : OAI211_X1 port map( C1 => n7675, C2 => n7669, A => n7668, B => n1963
                           , ZN => n6003);
   U2179 : NOR3_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_4_port, 
                           A3 => n1895, ZN => n6004);
   U2180 : NOR2_X1 port map( A1 => n7670, A2 => n7829, ZN => n6018);
   U2181 : NOR2_X1 port map( A1 => n7672, A2 => n7671, ZN => n6023);
   U2182 : OAI21_X1 port map( B1 => n7675, B2 => n7674, A => n7673, ZN => n1969
                           );
   U2183 : OAI21_X1 port map( B1 => n7678, B2 => n7677, A => n7676, ZN => n1962
                           );
   U2184 : AOI211_X1 port map( C1 => n7827, C2 => DATA1(0), A => n7680, B => 
                           n7679, ZN => n7683);
   U2185 : NAND3_X1 port map( A1 => n7683, A2 => n7682, A3 => n7681, ZN => 
                           n1938);
   U2186 : NOR2_X1 port map( A1 => n1933, A2 => n7711, ZN => n7689);
   U2187 : AOI211_X1 port map( C1 => DATA1(14), C2 => n7709, A => n7684, B => 
                           n7689, ZN => n7686);
   U2188 : OAI211_X1 port map( C1 => n7708, C2 => n7687, A => n7686, B => n7685
                           , ZN => n1932);
   U2189 : NOR2_X1 port map( A1 => n7688, A2 => n7687, ZN => n7690);
   U2190 : AOI211_X1 port map( C1 => n7691, C2 => DATA1(14), A => n7690, B => 
                           n7689, ZN => n7694);
   U2191 : NAND2_X1 port map( A1 => DATA1(16), A2 => n7692, ZN => n7693);
   U2192 : OAI211_X1 port map( C1 => n7696, C2 => n7695, A => n7694, B => n7693
                           , ZN => n1931);
   U2193 : OAI211_X1 port map( C1 => n7707, C2 => n1925, A => n7698, B => n7697
                           , ZN => n7699);
   U2194 : AOI211_X1 port map( C1 => DATA1(22), C2 => n7709, A => n7700, B => 
                           n7699, ZN => n1917);
   U2195 : INV_X1 port map( A => n7701, ZN => n7706);
   U2196 : NAND3_X1 port map( A1 => n7704, A2 => n7703, A3 => n7702, ZN => 
                           n7705);
   U2197 : AOI211_X1 port map( C1 => DATA1(23), C2 => n7709, A => n7706, B => 
                           n7705, ZN => n1913);
   U2198 : NAND2_X1 port map( A1 => DATA1(26), A2 => n7825, ZN => n1556);
   U2199 : NOR2_X1 port map( A1 => n7707, A2 => n1907, ZN => n1203);
   U2200 : NOR2_X1 port map( A1 => n1911, A2 => n7708, ZN => n1559);
   U2201 : AOI211_X1 port map( C1 => DATA1(23), C2 => n7709, A => n1203, B => 
                           n1559, ZN => n7710);
   U2202 : OAI211_X1 port map( C1 => n7711, C2 => n1912, A => n7710, B => n1556
                           , ZN => n1908);
   U2203 : AOI21_X1 port map( B1 => n7714, B2 => n7713, A => n7712, ZN => n1862
                           );
   U2204 : AOI22_X1 port map( A1 => n7717, A2 => n7716, B1 => n1856, B2 => 
                           n7715, ZN => n1851);
   U2205 : INV_X1 port map( A => DATA2_I_27_port, ZN => n7718);
   U2206 : NOR2_X1 port map( A1 => n1907, A2 => n7718, ZN => n1840);
   U2207 : AOI21_X1 port map( B1 => n1907, B2 => n7718, A => n1840, ZN => n1841
                           );

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3987, n3991, n3994, n3997, n4000, n4005, n4009, n4034, n4039, n4043,
      n4046, n4049, n4052, n4055, n4059, n4063, n4067, n4071, n4075, n4079, 
      n4090, n4094, n4097, n4102, n4110, n4115, n4120, n4125, n4130, n4135, 
      n4140, n4177, n4442, n4621, n4710, n4754, n4803, n4804, n4825, n4855, 
      n4856, n4876, n4881, n4882, n4883, n4905, n4906, n4920, n5570, n5594, 
      n5599, n5624, n5625, n5645, n5648, n5654, n5655, n5686, n5688, n5694, 
      n5696, n5697, n5699, n5700, n9015, n9016, n9017, n9018, n9019, n9020, 
      n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, 
      n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, 
      n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, 
      n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, 
      n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, 
      n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, 
      n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, 
      n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, 
      n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, 
      n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, 
      n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, 
      n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, 
      n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, 
      n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, 
      n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, 
      n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, 
      n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, 
      n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, 
      n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, 
      n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, 
      n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, 
      n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, 
      n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, 
      n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, 
      n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, 
      n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, 
      n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, 
      n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, 
      n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, 
      n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, 
      n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, 
      n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, 
      n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, 
      n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, 
      n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, 
      n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, 
      n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, 
      n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, 
      n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, 
      n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, 
      n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, 
      n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, 
      n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, 
      n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, 
      n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, 
      n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, 
      n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, 
      n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, 
      n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, 
      n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, 
      n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, 
      n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, 
      n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, 
      n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, 
      n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, 
      n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, 
      n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, 
      n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, 
      n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, 
      n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, 
      n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, 
      n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, 
      n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, 
      n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, 
      n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, 
      n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, 
      n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, 
      n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, 
      n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, 
      n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, 
      n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, 
      n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, 
      n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, 
      n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, 
      n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, 
      n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, 
      n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, 
      n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, 
      n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, 
      n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, 
      n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, 
      n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, 
      n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, 
      n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, 
      n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, 
      n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, 
      n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, 
      n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, 
      n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, 
      n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, 
      n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, 
      n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, 
      n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, 
      n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, 
      n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, 
      n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, 
      n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, 
      n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, 
      n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, 
      n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, 
      n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, 
      n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, 
      n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, 
      n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, 
      n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, 
      n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, 
      n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, 
      n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, 
      n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, 
      n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, 
      n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, 
      n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, 
      n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, 
      n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, 
      n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, 
      n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, 
      n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, 
      n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, 
      n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, 
      n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, 
      n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, 
      n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, 
      n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, 
      n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, 
      n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, 
      n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, 
      n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, 
      n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, 
      n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, 
      n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, 
      n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, 
      n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, 
      n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, 
      n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, 
      n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, 
      n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, 
      n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, 
      n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, 
      n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, 
      n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, 
      n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, 
      n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, 
      n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, 
      n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, 
      n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, 
      n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, 
      n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, 
      n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, 
      n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, 
      n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, 
      n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, 
      n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, 
      n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, 
      n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, 
      n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, 
      n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, 
      n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, 
      n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, 
      n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, 
      n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, 
      n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, 
      n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, 
      n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, 
      n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, 
      n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, 
      n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, 
      n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, 
      n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, 
      n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, 
      n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, 
      n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, 
      n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, 
      n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, 
      n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, 
      n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, 
      n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, 
      n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, 
      n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, 
      n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, 
      n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, 
      n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, 
      n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, 
      n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, 
      n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, 
      n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, 
      n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, 
      n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, 
      n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, 
      n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, 
      n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, 
      n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, 
      n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, 
      n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, 
      n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, 
      n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, 
      n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, 
      n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, 
      n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, 
      n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, 
      n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, 
      n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, 
      n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, 
      n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, 
      n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, 
      n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, 
      n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, 
      n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, 
      n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, 
      n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, 
      n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, 
      n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, 
      n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, 
      n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, 
      n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, 
      n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, 
      n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, 
      n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, 
      n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, 
      n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, 
      n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, 
      n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, 
      n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, 
      n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, 
      n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, 
      n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, 
      n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, 
      n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, 
      n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, 
      n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, 
      n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, 
      n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, 
      n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, 
      n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, 
      n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, 
      n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, 
      n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, 
      n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, 
      n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, 
      n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, 
      n11270, n11272, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
      n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
      n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
      n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
      n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
      n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
      n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
      n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
      n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
      n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
      n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
      n3567, n3568, n3569, n3570, n3571, n3572, n3574, n3575, n3576, n3577, 
      n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, 
      n3588, n3589, n3590, n3591, n13461, n13462, n13463, n13464, n13465, 
      n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, 
      n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, 
      n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, 
      n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, 
      n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, 
      n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, 
      n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, 
      n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, 
      n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, 
      n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, 
      n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, 
      n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, 
      n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, 
      n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, 
      n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, 
      n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, 
      n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, 
      n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, 
      n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, 
      n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, 
      n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, 
      n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, 
      n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, 
      n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, 
      n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, 
      n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, 
      n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, 
      n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, 
      n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, 
      n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, 
      n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, 
      n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, 
      n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, 
      n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, 
      n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, 
      n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, 
      n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, 
      n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, 
      n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, 
      n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, 
      n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, 
      n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, 
      n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, 
      n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, 
      n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, 
      n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, 
      n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, 
      n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, 
      n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, 
      n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, 
      n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, 
      n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, 
      n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, 
      n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, 
      n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, 
      n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, 
      n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, 
      n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, 
      n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, 
      n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, 
      n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, 
      n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, 
      n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, 
      n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, 
      n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, 
      n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, 
      n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, 
      n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, 
      n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, 
      n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, 
      n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, 
      n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, 
      n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, 
      n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, 
      n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, 
      n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, 
      n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, 
      n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, 
      n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, 
      n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, 
      n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, 
      n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, 
      n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, 
      n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, 
      n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, 
      n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, 
      n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, 
      n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, 
      n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, 
      n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, 
      n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, 
      n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, 
      n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, 
      n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, 
      n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, 
      n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, 
      n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, 
      n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, 
      n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, 
      n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, 
      n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, 
      n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, 
      n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, 
      n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, 
      n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, 
      n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, 
      n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, 
      n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, 
      n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, 
      n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, 
      n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, 
      n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, 
      n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, 
      n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, 
      n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, 
      n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, 
      n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, 
      n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, 
      n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, 
      n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, 
      n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, 
      n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, 
      n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, 
      n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, 
      n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, 
      n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, 
      n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, 
      n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, 
      n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, 
      n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, 
      n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, 
      n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, 
      n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, 
      n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, 
      n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, 
      n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, 
      n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, 
      n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, 
      n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, 
      n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, 
      n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, 
      n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, 
      n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, 
      n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, 
      n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, 
      n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, 
      n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, 
      n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, 
      n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, 
      n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, 
      n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, 
      n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, 
      n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, 
      n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, 
      n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, 
      n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, 
      n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, 
      n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, 
      n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, 
      n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, 
      n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, 
      n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, 
      n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, 
      n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, 
      n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, 
      n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, 
      n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, 
      n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, 
      n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, 
      n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, 
      n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, 
      n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, 
      n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, 
      n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, 
      n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, 
      n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, 
      n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, 
      n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, 
      n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, 
      n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, 
      n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, 
      n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, 
      n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, 
      n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, 
      n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, 
      n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, 
      n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, 
      n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, 
      n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, 
      n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, 
      n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, 
      n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, 
      n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, 
      n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, 
      n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, 
      n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, 
      n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, 
      n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, 
      n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, 
      n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, 
      n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, 
      n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, 
      n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, 
      n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, 
      n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, 
      n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, 
      n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, 
      n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, 
      n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, 
      n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, 
      n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, 
      n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, 
      n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, 
      n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, 
      n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, 
      n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, 
      n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, 
      n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, 
      n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, 
      n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, 
      n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, 
      n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, 
      n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, 
      n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, 
      n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, 
      n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, 
      n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, 
      n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, 
      n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, 
      n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, 
      n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, 
      n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, 
      n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, 
      n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, 
      n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, 
      n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, 
      n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, 
      n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, 
      n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, 
      n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, 
      n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, 
      n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, 
      n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, 
      n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, 
      n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, 
      n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, 
      n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, 
      n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, 
      n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, 
      n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, 
      n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, 
      n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, 
      n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, 
      n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, 
      n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, 
      n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, 
      n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, 
      n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, 
      n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, 
      n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, 
      n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, 
      n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, 
      n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, 
      n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, 
      n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, 
      n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, 
      n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, 
      n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, 
      n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, 
      n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, 
      n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, 
      n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, 
      n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, 
      n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, 
      n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, 
      n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, 
      n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, 
      n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, 
      n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, 
      n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, 
      n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, 
      n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, 
      n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, 
      n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, 
      n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, 
      n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, 
      n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, 
      n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, 
      n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, 
      n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, 
      n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, 
      n16085, n16086, n16087, n16088, n16089, n16090, n_1672, n_1673, n_1674, 
      n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, 
      n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, 
      n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, 
      n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, 
      n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, 
      n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, 
      n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, 
      n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, 
      n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, 
      n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, 
      n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, 
      n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, 
      n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, 
      n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, 
      n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, 
      n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, 
      n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, 
      n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, 
      n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, 
      n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, 
      n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, 
      n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, 
      n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, 
      n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, 
      n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, 
      n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, 
      n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, 
      n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, 
      n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, 
      n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, 
      n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, 
      n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, 
      n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, 
      n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, 
      n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, 
      n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, 
      n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, 
      n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, 
      n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, 
      n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, 
      n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, 
      n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, 
      n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, 
      n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, 
      n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, 
      n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, 
      n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, 
      n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, 
      n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, 
      n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, 
      n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, 
      n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, 
      n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, 
      n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, 
      n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, 
      n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, 
      n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, 
      n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, 
      n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, 
      n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, 
      n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, 
      n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, 
      n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, 
      n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, 
      n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, 
      n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, 
      n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, 
      n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, 
      n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, 
      n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, 
      n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, 
      n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, 
      n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, 
      n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, 
      n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, 
      n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, 
      n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, 
      n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, 
      n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, 
      n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, 
      n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, 
      n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, 
      n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, 
      n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, 
      n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, 
      n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, 
      n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, 
      n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, 
      n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, 
      n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, 
      n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, 
      n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, 
      n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, 
      n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, 
      n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, 
      n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, 
      n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, 
      n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, 
      n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, 
      n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, 
      n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, 
      n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, 
      n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, 
      n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, 
      n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, 
      n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, 
      n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, 
      n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, 
      n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, 
      n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, 
      n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, 
      n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, 
      n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, 
      n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, 
      n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, 
      n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, 
      n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, 
      n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, 
      n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, 
      n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, 
      n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, 
      n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, 
      n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, 
      n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, 
      n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, 
      n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, 
      n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, 
      n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, 
      n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, 
      n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, 
      n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, 
      n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, 
      n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, 
      n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, 
      n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, 
      n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, 
      n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, 
      n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, 
      n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, 
      n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, 
      n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, 
      n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, 
      n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, 
      n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, 
      n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, 
      n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, 
      n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, 
      n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, 
      n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, 
      n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, 
      n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, 
      n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, 
      n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, 
      n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, 
      n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, 
      n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, 
      n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, 
      n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, 
      n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, 
      n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, 
      n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, 
      n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, 
      n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, 
      n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, 
      n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, 
      n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, 
      n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, 
      n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, 
      n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, 
      n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, 
      n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, 
      n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, 
      n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, 
      n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, 
      n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, 
      n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, 
      n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, 
      n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, 
      n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, 
      n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, 
      n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, 
      n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, 
      n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, 
      n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, 
      n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, 
      n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, 
      n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, 
      n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, 
      n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, 
      n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, 
      n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, 
      n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402, 
      n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, 
      n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, 
      n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, 
      n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, 
      n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, 
      n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, 
      n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465, 
      n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, 
      n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, 
      n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, 
      n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, 
      n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, 
      n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, 
      n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, 
      n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, 
      n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, 
      n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, 
      n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, 
      n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, 
      n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, 
      n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, 
      n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, 
      n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, 
      n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, 
      n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, 
      n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, 
      n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645, 
      n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, n_3654, 
      n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, 
      n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, 
      n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, 
      n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, 
      n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, 
      n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, n_3708, 
      n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, n_3717, 
      n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, n_3726, 
      n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, 
      n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, 
      n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, 
      n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, 
      n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, 
      n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, 
      n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, 
      n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, 
      n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, 
      n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, 
      n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, 
      n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, 
      n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, n_3843, 
      n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, n_3852, 
      n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, 
      n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, n_3870, 
      n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, 
      n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, 
      n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, 
      n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906, 
      n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, 
      n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, n_3924, 
      n_3925, n_3926, n_3927, n_3928 : std_logic;

begin
   
   clk_r_REG3182_S2 : DFFR_X1 port map( D => ENABLE, CK => CLK, RN => RESET_BAR
                           , Q => n11272, QN => n_1672);
   clk_r_REG3247_S2 : DFFR_X1 port map( D => RD1, CK => CLK, RN => RESET_BAR, Q
                           => n11270, QN => n_1673);
   clk_r_REG3179_S1 : DFFR_X1 port map( D => RD2, CK => CLK, RN => RESET_BAR, Q
                           => n11269, QN => n_1674);
   clk_r_REG3491_S7 : DFFR_X1 port map( D => ADD_RD1(4), CK => CLK, RN => 
                           RESET_BAR, Q => n11268, QN => n_1675);
   clk_r_REG3493_S7 : DFFS_X1 port map( D => n3574, CK => CLK, SN => RESET_BAR,
                           Q => n_1676, QN => n11267);
   clk_r_REG3391_S7 : DFFR_X1 port map( D => ADD_RD2(4), CK => CLK, RN => 
                           RESET_BAR, Q => n11266, QN => n_1677);
   clk_r_REG3425_S7 : DFFS_X1 port map( D => n3583, CK => CLK, SN => RESET_BAR,
                           Q => n_1678, QN => n11265);
   clk_r_REG120_S53 : DFFR_X1 port map( D => DATAIN(31), CK => CLK, RN => 
                           RESET_BAR, Q => n11264, QN => n_1679);
   clk_r_REG2170_S52 : DFFR_X1 port map( D => DATAIN(30), CK => CLK, RN => 
                           RESET_BAR, Q => n11263, QN => n_1680);
   clk_r_REG2247_S50 : DFFR_X1 port map( D => DATAIN(29), CK => CLK, RN => 
                           RESET_BAR, Q => n11262, QN => n_1681);
   clk_r_REG2321_S49 : DFFR_X1 port map( D => DATAIN(28), CK => CLK, RN => 
                           RESET_BAR, Q => n11261, QN => n_1682);
   clk_r_REG2401_S47 : DFFR_X1 port map( D => DATAIN(27), CK => CLK, RN => 
                           RESET_BAR, Q => n11260, QN => n_1683);
   clk_r_REG2478_S46 : DFFR_X1 port map( D => DATAIN(26), CK => CLK, RN => 
                           RESET_BAR, Q => n11259, QN => n_1684);
   clk_r_REG2559_S44 : DFFR_X1 port map( D => DATAIN(25), CK => CLK, RN => 
                           RESET_BAR, Q => n11258, QN => n_1685);
   clk_r_REG2636_S43 : DFFR_X1 port map( D => DATAIN(24), CK => CLK, RN => 
                           RESET_BAR, Q => n11257, QN => n_1686);
   clk_r_REG1796_S43 : DFFR_X1 port map( D => DATAIN(23), CK => CLK, RN => 
                           RESET_BAR, Q => n11256, QN => n_1687);
   clk_r_REG1868_S42 : DFFR_X1 port map( D => DATAIN(22), CK => CLK, RN => 
                           RESET_BAR, Q => n11255, QN => n_1688);
   clk_r_REG1945_S36 : DFFR_X1 port map( D => DATAIN(21), CK => CLK, RN => 
                           RESET_BAR, Q => n11254, QN => n_1689);
   clk_r_REG2717_S39 : DFFR_X1 port map( D => DATAIN(20), CK => CLK, RN => 
                           RESET_BAR, Q => n11253, QN => n_1690);
   clk_r_REG2793_S37 : DFFR_X1 port map( D => DATAIN(19), CK => CLK, RN => 
                           RESET_BAR, Q => n11252, QN => n_1691);
   clk_r_REG2866_S36 : DFFR_X1 port map( D => DATAIN(18), CK => CLK, RN => 
                           RESET_BAR, Q => n11251, QN => n_1692);
   clk_r_REG2017_S36 : DFFR_X1 port map( D => DATAIN(17), CK => CLK, RN => 
                           RESET_BAR, Q => n11250, QN => n_1693);
   clk_r_REG2943_S33 : DFFR_X1 port map( D => DATAIN(16), CK => CLK, RN => 
                           RESET_BAR, Q => n11249, QN => n_1694);
   clk_r_REG1558_S9 : DFFR_X1 port map( D => DATAIN(15), CK => CLK, RN => 
                           RESET_BAR, Q => n11248, QN => n_1695);
   clk_r_REG1634_S8 : DFFR_X1 port map( D => DATAIN(14), CK => CLK, RN => 
                           RESET_BAR, Q => n11247, QN => n_1696);
   clk_r_REG1380_S8 : DFFR_X1 port map( D => DATAIN(13), CK => CLK, RN => 
                           RESET_BAR, Q => n11246, QN => n_1697);
   clk_r_REG1720_S8 : DFFR_X1 port map( D => DATAIN(12), CK => CLK, RN => 
                           RESET_BAR, Q => n11245, QN => n_1698);
   clk_r_REG999_S25 : DFFR_X1 port map( D => DATAIN(11), CK => CLK, RN => 
                           RESET_BAR, Q => n11244, QN => n_1699);
   clk_r_REG1074_S21 : DFFR_X1 port map( D => DATAIN(10), CK => CLK, RN => 
                           RESET_BAR, Q => n11243, QN => n_1700);
   clk_r_REG745_S7 : DFFR_X1 port map( D => DATAIN(9), CK => CLK, RN => 
                           RESET_BAR, Q => n11242, QN => n_1701);
   clk_r_REG823_S11 : DFFR_X1 port map( D => DATAIN(8), CK => CLK, RN => 
                           RESET_BAR, Q => n11241, QN => n_1702);
   clk_r_REG384_S11 : DFFR_X1 port map( D => DATAIN(7), CK => CLK, RN => 
                           RESET_BAR, Q => n11240, QN => n_1703);
   clk_r_REG1221_S8 : DFFR_X1 port map( D => DATAIN(6), CK => CLK, RN => 
                           RESET_BAR, Q => n11239, QN => n_1704);
   clk_r_REG520_S8 : DFFR_X1 port map( D => DATAIN(5), CK => CLK, RN => 
                           RESET_BAR, Q => n11238, QN => n_1705);
   clk_r_REG904_S9 : DFFR_X1 port map( D => DATAIN(4), CK => CLK, RN => 
                           RESET_BAR, Q => n11237, QN => n_1706);
   clk_r_REG357_S8 : DFFR_X1 port map( D => DATAIN(3), CK => CLK, RN => 
                           RESET_BAR, Q => n11236, QN => n_1707);
   clk_r_REG1485_S11 : DFFR_X1 port map( D => DATAIN(2), CK => CLK, RN => 
                           RESET_BAR, Q => n11235, QN => n_1708);
   clk_r_REG3037_S15 : DFFR_X1 port map( D => DATAIN(1), CK => CLK, RN => 
                           RESET_BAR, Q => n11234, QN => n_1709);
   clk_r_REG3112_S13 : DFFR_X1 port map( D => DATAIN(0), CK => CLK, RN => 
                           RESET_BAR, Q => n11233, QN => n_1710);
   clk_r_REG3246_S2 : DFFS_X1 port map( D => n3987, CK => CLK, SN => RESET_BAR,
                           Q => n11221, QN => n_1711);
   clk_r_REG3426_S7 : DFFS_X1 port map( D => n3583, CK => CLK, SN => RESET_BAR,
                           Q => n11192, QN => n_1712);
   clk_r_REG3403_S7 : DFFR_X1 port map( D => n4710, CK => CLK, RN => RESET_BAR,
                           Q => n11191, QN => n_1713);
   clk_r_REG3397_S7 : DFFR_X1 port map( D => n4881, CK => CLK, RN => RESET_BAR,
                           Q => n11190, QN => n_1714);
   clk_r_REG3393_S7 : DFFR_X1 port map( D => n4855, CK => CLK, RN => RESET_BAR,
                           Q => n11189, QN => n_1715);
   clk_r_REG3415_S7 : DFFR_X1 port map( D => n4883, CK => CLK, RN => RESET_BAR,
                           Q => n11188, QN => n_1716);
   clk_r_REG3413_S7 : DFFR_X1 port map( D => n4920, CK => CLK, RN => RESET_BAR,
                           Q => n11187, QN => n_1717);
   clk_r_REG3411_S7 : DFFR_X1 port map( D => n4876, CK => CLK, RN => RESET_BAR,
                           Q => n11186, QN => n_1718);
   clk_r_REG3433_S7 : DFFR_X1 port map( D => n3590, CK => CLK, RN => RESET_BAR,
                           Q => n11185, QN => n_1719);
   clk_r_REG3446_S7 : DFFR_X1 port map( D => n3586, CK => CLK, RN => RESET_BAR,
                           Q => n11184, QN => n_1720);
   clk_r_REG3443_S7 : DFFR_X1 port map( D => n3585, CK => CLK, RN => RESET_BAR,
                           Q => n11183, QN => n_1721);
   clk_r_REG3449_S7 : DFFR_X1 port map( D => n3587, CK => CLK, RN => RESET_BAR,
                           Q => n11182, QN => n_1722);
   clk_r_REG3430_S7 : DFFR_X1 port map( D => n3591, CK => CLK, RN => RESET_BAR,
                           Q => n11181, QN => n_1723);
   clk_r_REG3440_S7 : DFFR_X1 port map( D => n3584, CK => CLK, RN => RESET_BAR,
                           Q => n11180, QN => n_1724);
   clk_r_REG3442_S7 : DFFR_X1 port map( D => n3585, CK => CLK, RN => RESET_BAR,
                           Q => n11179, QN => n_1725);
   clk_r_REG3448_S7 : DFFR_X1 port map( D => n3587, CK => CLK, RN => RESET_BAR,
                           Q => n11178, QN => n_1726);
   clk_r_REG3439_S7 : DFFR_X1 port map( D => n3584, CK => CLK, RN => RESET_BAR,
                           Q => n11177, QN => n_1727);
   clk_r_REG3429_S7 : DFFR_X1 port map( D => n3591, CK => CLK, RN => RESET_BAR,
                           Q => n11176, QN => n_1728);
   clk_r_REG3423_S7 : DFFR_X1 port map( D => n4906, CK => CLK, RN => RESET_BAR,
                           Q => n11175, QN => n_1729);
   clk_r_REG3407_S7 : DFFR_X1 port map( D => n4754, CK => CLK, RN => RESET_BAR,
                           Q => n11174, QN => n_1730);
   clk_r_REG3405_S7 : DFFR_X1 port map( D => n4803, CK => CLK, RN => RESET_BAR,
                           Q => n11173, QN => n_1731);
   clk_r_REG3401_S7 : DFFR_X1 port map( D => n4621, CK => CLK, RN => RESET_BAR,
                           Q => n11172, QN => n_1732);
   clk_r_REG3445_S7 : DFFR_X1 port map( D => n3586, CK => CLK, RN => RESET_BAR,
                           Q => n11171, QN => n_1733);
   clk_r_REG3432_S7 : DFFR_X1 port map( D => n3590, CK => CLK, RN => RESET_BAR,
                           Q => n11170, QN => n_1734);
   clk_r_REG3428_S7 : DFFR_X1 port map( D => n3591, CK => CLK, RN => RESET_BAR,
                           Q => n11169, QN => n_1735);
   clk_r_REG3421_S7 : DFFR_X1 port map( D => n4882, CK => CLK, RN => RESET_BAR,
                           Q => n11168, QN => n_1736);
   clk_r_REG3417_S7 : DFFR_X1 port map( D => n4856, CK => CLK, RN => RESET_BAR,
                           Q => n11167, QN => n_1737);
   clk_r_REG3399_S7 : DFFR_X1 port map( D => n4825, CK => CLK, RN => RESET_BAR,
                           Q => n11166, QN => n_1738);
   clk_r_REG3419_S7 : DFFR_X1 port map( D => n4905, CK => CLK, RN => RESET_BAR,
                           Q => n11165, QN => n_1739);
   clk_r_REG3438_S7 : DFFR_X1 port map( D => n3584, CK => CLK, RN => RESET_BAR,
                           Q => n11164, QN => n_1740);
   clk_r_REG3441_S7 : DFFR_X1 port map( D => n3585, CK => CLK, RN => RESET_BAR,
                           Q => n11163, QN => n_1741);
   clk_r_REG3409_S7 : DFFR_X1 port map( D => n4804, CK => CLK, RN => RESET_BAR,
                           Q => n11162, QN => n_1742);
   clk_r_REG3447_S7 : DFFR_X1 port map( D => n3587, CK => CLK, RN => RESET_BAR,
                           Q => n11161, QN => n_1743);
   clk_r_REG3444_S7 : DFFR_X1 port map( D => n3586, CK => CLK, RN => RESET_BAR,
                           Q => n11160, QN => n_1744);
   clk_r_REG3431_S7 : DFFR_X1 port map( D => n3590, CK => CLK, RN => RESET_BAR,
                           Q => n11159, QN => n_1745);
   clk_r_REG3435_S7 : DFFS_X1 port map( D => n3589, CK => CLK, SN => RESET_BAR,
                           Q => n11158, QN => n_1746);
   clk_r_REG3395_S7 : DFFR_X1 port map( D => n4442, CK => CLK, RN => RESET_BAR,
                           Q => n11157, QN => n_1747);
   clk_r_REG3437_S7 : DFFR_X1 port map( D => n3588, CK => CLK, RN => RESET_BAR,
                           Q => n11156, QN => n_1748);
   clk_r_REG3494_S7 : DFFS_X1 port map( D => n3574, CK => CLK, SN => RESET_BAR,
                           Q => n11155, QN => n_1749);
   clk_r_REG3375_S7 : DFFR_X1 port map( D => n5599, CK => CLK, RN => RESET_BAR,
                           Q => n11154, QN => n_1750);
   clk_r_REG3379_S7 : DFFR_X1 port map( D => n5688, CK => CLK, RN => RESET_BAR,
                           Q => n11153, QN => n_1751);
   clk_r_REG3341_S7 : DFFR_X1 port map( D => n5697, CK => CLK, RN => RESET_BAR,
                           Q => n11152, QN => n_1752);
   clk_r_REG3377_S7 : DFFR_X1 port map( D => n5645, CK => CLK, RN => RESET_BAR,
                           Q => n11151, QN => n_1753);
   clk_r_REG3339_S7 : DFFR_X1 port map( D => n5624, CK => CLK, RN => RESET_BAR,
                           Q => n11150, QN => n_1754);
   clk_r_REG3360_S7 : DFFR_X1 port map( D => n5696, CK => CLK, RN => RESET_BAR,
                           Q => n11149, QN => n_1755);
   clk_r_REG3371_S7 : DFFR_X1 port map( D => n3578, CK => CLK, RN => RESET_BAR,
                           Q => n11148, QN => n_1756);
   clk_r_REG3358_S7 : DFFR_X1 port map( D => n3576, CK => CLK, RN => RESET_BAR,
                           Q => n11147, QN => n_1757);
   clk_r_REG3387_S7 : DFFS_X1 port map( D => n3579, CK => CLK, SN => RESET_BAR,
                           Q => n11146, QN => n_1758);
   clk_r_REG3357_S7 : DFFR_X1 port map( D => n3576, CK => CLK, RN => RESET_BAR,
                           Q => n11145, QN => n_1759);
   clk_r_REG3370_S7 : DFFR_X1 port map( D => n3578, CK => CLK, RN => RESET_BAR,
                           Q => n11144, QN => n_1760);
   clk_r_REG3351_S7 : DFFR_X1 port map( D => n5625, CK => CLK, RN => RESET_BAR,
                           Q => n11143, QN => n_1761);
   clk_r_REG3345_S7 : DFFR_X1 port map( D => n5655, CK => CLK, RN => RESET_BAR,
                           Q => n11142, QN => n_1762);
   clk_r_REG3366_S7 : DFFR_X1 port map( D => n5686, CK => CLK, RN => RESET_BAR,
                           Q => n11141, QN => n_1763);
   clk_r_REG3364_S7 : DFFR_X1 port map( D => n5694, CK => CLK, RN => RESET_BAR,
                           Q => n11140, QN => n_1764);
   clk_r_REG3347_S7 : DFFR_X1 port map( D => n5654, CK => CLK, RN => RESET_BAR,
                           Q => n11139, QN => n_1765);
   clk_r_REG3362_S7 : DFFR_X1 port map( D => n5594, CK => CLK, RN => RESET_BAR,
                           Q => n11138, QN => n_1766);
   clk_r_REG3373_S7 : DFFR_X1 port map( D => n5648, CK => CLK, RN => RESET_BAR,
                           Q => n11137, QN => n_1767);
   clk_r_REG3383_S7 : DFFR_X1 port map( D => n5700, CK => CLK, RN => RESET_BAR,
                           Q => n11136, QN => n_1768);
   clk_r_REG3368_S7 : DFFR_X1 port map( D => n3577, CK => CLK, RN => RESET_BAR,
                           Q => n11135, QN => n_1769);
   clk_r_REG3343_S7 : DFFR_X1 port map( D => n3582, CK => CLK, RN => RESET_BAR,
                           Q => n11134, QN => n_1770);
   clk_r_REG3353_S7 : DFFR_X1 port map( D => n5570, CK => CLK, RN => RESET_BAR,
                           Q => n11133, QN => n_1771);
   clk_r_REG3385_S7 : DFFR_X1 port map( D => n5699, CK => CLK, RN => RESET_BAR,
                           Q => n11132, QN => n_1772);
   clk_r_REG3349_S7 : DFFR_X1 port map( D => n3581, CK => CLK, RN => RESET_BAR,
                           Q => n11131, QN => n_1773);
   clk_r_REG3355_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR,
                           Q => n11130, QN => n_1774);
   clk_r_REG3381_S7 : DFFR_X1 port map( D => n3580, CK => CLK, RN => RESET_BAR,
                           Q => n11129, QN => n_1775);
   clk_r_REG3369_S7 : DFFR_X1 port map( D => n3578, CK => CLK, RN => RESET_BAR,
                           Q => n11128, QN => n_1776);
   clk_r_REG3356_S7 : DFFR_X1 port map( D => n3576, CK => CLK, RN => RESET_BAR,
                           Q => n11127, QN => n_1777);
   clk_r_REG1709_S1 : DFF_X1 port map( D => n3100, CK => CLK, Q => n11126, QN 
                           => n_1778);
   clk_r_REG2936_S1 : DFF_X1 port map( D => n2972, CK => CLK, Q => n11125, QN 
                           => n_1779);
   clk_r_REG122_S1 : DFF_X1 port map( D => n2549, CK => CLK, Q => n11124, QN =>
                           n_1780);
   clk_r_REG2692_S1 : DFF_X1 port map( D => n2773, CK => CLK, Q => n11123, QN 
                           => n_1781);
   clk_r_REG2116_S1 : DFF_X1 port map( D => n2554, CK => CLK, Q => n11122, QN 
                           => n_1782);
   clk_r_REG726_S1 : DFF_X1 port map( D => n3387, CK => CLK, Q => n11121, QN =>
                           n_1783);
   clk_r_REG724_S1 : DFF_X1 port map( D => n3388, CK => CLK, Q => n11120, QN =>
                           n_1784);
   clk_r_REG906_S1 : DFF_X1 port map( D => n3444, CK => CLK, Q => n11119, QN =>
                           n_1785);
   clk_r_REG937_S1 : DFF_X1 port map( D => n3443, CK => CLK, Q => n11118, QN =>
                           n_1786);
   clk_r_REG939_S1 : DFF_X1 port map( D => n3442, CK => CLK, Q => n11117, QN =>
                           n_1787);
   clk_r_REG941_S1 : DFF_X1 port map( D => n3441, CK => CLK, Q => n11116, QN =>
                           n_1788);
   clk_r_REG943_S1 : DFF_X1 port map( D => n3440, CK => CLK, Q => n11115, QN =>
                           n_1789);
   clk_r_REG945_S1 : DFF_X1 port map( D => n3439, CK => CLK, Q => n11114, QN =>
                           n_1790);
   clk_r_REG947_S1 : DFF_X1 port map( D => n3438, CK => CLK, Q => n11113, QN =>
                           n_1791);
   clk_r_REG714_S1 : DFF_X1 port map( D => n3393, CK => CLK, Q => n11112, QN =>
                           n_1792);
   clk_r_REG716_S1 : DFF_X1 port map( D => n3392, CK => CLK, Q => n11111, QN =>
                           n_1793);
   clk_r_REG718_S1 : DFF_X1 port map( D => n3391, CK => CLK, Q => n11110, QN =>
                           n_1794);
   clk_r_REG720_S1 : DFF_X1 port map( D => n3390, CK => CLK, Q => n11109, QN =>
                           n_1795);
   clk_r_REG722_S1 : DFF_X1 port map( D => n3389, CK => CLK, Q => n11108, QN =>
                           n_1796);
   clk_r_REG738_S1 : DFF_X1 port map( D => n3381, CK => CLK, Q => n11107, QN =>
                           n_1797);
   clk_r_REG736_S1 : DFF_X1 port map( D => n3382, CK => CLK, Q => n11106, QN =>
                           n_1798);
   clk_r_REG734_S1 : DFF_X1 port map( D => n3383, CK => CLK, Q => n11105, QN =>
                           n_1799);
   clk_r_REG732_S1 : DFF_X1 port map( D => n3384, CK => CLK, Q => n11104, QN =>
                           n_1800);
   clk_r_REG730_S1 : DFF_X1 port map( D => n3385, CK => CLK, Q => n11103, QN =>
                           n_1801);
   clk_r_REG728_S1 : DFF_X1 port map( D => n3386, CK => CLK, Q => n11102, QN =>
                           n_1802);
   clk_r_REG692_S1 : DFF_X1 port map( D => n3404, CK => CLK, Q => n11101, QN =>
                           n_1803);
   clk_r_REG694_S1 : DFF_X1 port map( D => n3403, CK => CLK, Q => n11100, QN =>
                           n_1804);
   clk_r_REG696_S1 : DFF_X1 port map( D => n3402, CK => CLK, Q => n11099, QN =>
                           n_1805);
   clk_r_REG698_S1 : DFF_X1 port map( D => n3401, CK => CLK, Q => n11098, QN =>
                           n_1806);
   clk_r_REG700_S1 : DFF_X1 port map( D => n3400, CK => CLK, Q => n11097, QN =>
                           n_1807);
   clk_r_REG702_S1 : DFF_X1 port map( D => n3399, CK => CLK, Q => n11096, QN =>
                           n_1808);
   clk_r_REG704_S1 : DFF_X1 port map( D => n3398, CK => CLK, Q => n11095, QN =>
                           n_1809);
   clk_r_REG706_S1 : DFF_X1 port map( D => n3397, CK => CLK, Q => n11094, QN =>
                           n_1810);
   clk_r_REG708_S1 : DFF_X1 port map( D => n3396, CK => CLK, Q => n11093, QN =>
                           n_1811);
   clk_r_REG710_S1 : DFF_X1 port map( D => n3395, CK => CLK, Q => n11092, QN =>
                           n_1812);
   clk_r_REG712_S1 : DFF_X1 port map( D => n3394, CK => CLK, Q => n11091, QN =>
                           n_1813);
   clk_r_REG1277_S1 : DFF_X1 port map( D => n3356, CK => CLK, Q => n11090, QN 
                           => n_1814);
   clk_r_REG522_S1 : DFF_X1 port map( D => n3412, CK => CLK, Q => n11089, QN =>
                           n_1815);
   clk_r_REG678_S1 : DFF_X1 port map( D => n3411, CK => CLK, Q => n11088, QN =>
                           n_1816);
   clk_r_REG680_S1 : DFF_X1 port map( D => n3410, CK => CLK, Q => n11087, QN =>
                           n_1817);
   clk_r_REG682_S1 : DFF_X1 port map( D => n3409, CK => CLK, Q => n11086, QN =>
                           n_1818);
   clk_r_REG684_S1 : DFF_X1 port map( D => n3408, CK => CLK, Q => n11085, QN =>
                           n_1819);
   clk_r_REG686_S1 : DFF_X1 port map( D => n3407, CK => CLK, Q => n11084, QN =>
                           n_1820);
   clk_r_REG688_S1 : DFF_X1 port map( D => n3406, CK => CLK, Q => n11083, QN =>
                           n_1821);
   clk_r_REG690_S1 : DFF_X1 port map( D => n3405, CK => CLK, Q => n11082, QN =>
                           n_1822);
   clk_r_REG1269_S1 : DFF_X1 port map( D => n3360, CK => CLK, Q => n11081, QN 
                           => n_1823);
   clk_r_REG1271_S1 : DFF_X1 port map( D => n3359, CK => CLK, Q => n11080, QN 
                           => n_1824);
   clk_r_REG1273_S1 : DFF_X1 port map( D => n3358, CK => CLK, Q => n11079, QN 
                           => n_1825);
   clk_r_REG1275_S1 : DFF_X1 port map( D => n3357, CK => CLK, Q => n11078, QN 
                           => n_1826);
   clk_r_REG1291_S1 : DFF_X1 port map( D => n3349, CK => CLK, Q => n11077, QN 
                           => n_1827);
   clk_r_REG1289_S1 : DFF_X1 port map( D => n3350, CK => CLK, Q => n11076, QN 
                           => n_1828);
   clk_r_REG1287_S1 : DFF_X1 port map( D => n3351, CK => CLK, Q => n11075, QN 
                           => n_1829);
   clk_r_REG1285_S1 : DFF_X1 port map( D => n3352, CK => CLK, Q => n11074, QN 
                           => n_1830);
   clk_r_REG1283_S1 : DFF_X1 port map( D => n3353, CK => CLK, Q => n11073, QN 
                           => n_1831);
   clk_r_REG1281_S1 : DFF_X1 port map( D => n3354, CK => CLK, Q => n11072, QN 
                           => n_1832);
   clk_r_REG1279_S1 : DFF_X1 port map( D => n3355, CK => CLK, Q => n11071, QN 
                           => n_1833);
   clk_r_REG1247_S1 : DFF_X1 port map( D => n3371, CK => CLK, Q => n11070, QN 
                           => n_1834);
   clk_r_REG1249_S1 : DFF_X1 port map( D => n3370, CK => CLK, Q => n11069, QN 
                           => n_1835);
   clk_r_REG1251_S1 : DFF_X1 port map( D => n3369, CK => CLK, Q => n11068, QN 
                           => n_1836);
   clk_r_REG1253_S1 : DFF_X1 port map( D => n3368, CK => CLK, Q => n11067, QN 
                           => n_1837);
   clk_r_REG1255_S1 : DFF_X1 port map( D => n3367, CK => CLK, Q => n11066, QN 
                           => n_1838);
   clk_r_REG1257_S1 : DFF_X1 port map( D => n3366, CK => CLK, Q => n11065, QN 
                           => n_1839);
   clk_r_REG1259_S1 : DFF_X1 port map( D => n3365, CK => CLK, Q => n11064, QN 
                           => n_1840);
   clk_r_REG1261_S1 : DFF_X1 port map( D => n3364, CK => CLK, Q => n11063, QN 
                           => n_1841);
   clk_r_REG1263_S1 : DFF_X1 port map( D => n3363, CK => CLK, Q => n11062, QN 
                           => n_1842);
   clk_r_REG1265_S1 : DFF_X1 port map( D => n3362, CK => CLK, Q => n11061, QN 
                           => n_1843);
   clk_r_REG1267_S1 : DFF_X1 port map( D => n3361, CK => CLK, Q => n11060, QN 
                           => n_1844);
   clk_r_REG1223_S1 : DFF_X1 port map( D => n3380, CK => CLK, Q => n11059, QN 
                           => n_1845);
   clk_r_REG1231_S1 : DFF_X1 port map( D => n3379, CK => CLK, Q => n11058, QN 
                           => n_1846);
   clk_r_REG1233_S1 : DFF_X1 port map( D => n3378, CK => CLK, Q => n11057, QN 
                           => n_1847);
   clk_r_REG1235_S1 : DFF_X1 port map( D => n3377, CK => CLK, Q => n11056, QN 
                           => n_1848);
   clk_r_REG1237_S1 : DFF_X1 port map( D => n3376, CK => CLK, Q => n11055, QN 
                           => n_1849);
   clk_r_REG1239_S1 : DFF_X1 port map( D => n3375, CK => CLK, Q => n11054, QN 
                           => n_1850);
   clk_r_REG1241_S1 : DFF_X1 port map( D => n3374, CK => CLK, Q => n11053, QN 
                           => n_1851);
   clk_r_REG1243_S1 : DFF_X1 port map( D => n3373, CK => CLK, Q => n11052, QN 
                           => n_1852);
   clk_r_REG1245_S1 : DFF_X1 port map( D => n3372, CK => CLK, Q => n11051, QN 
                           => n_1853);
   clk_r_REG1191_S1 : DFF_X1 port map( D => n3327, CK => CLK, Q => n11050, QN 
                           => n_1854);
   clk_r_REG1193_S1 : DFF_X1 port map( D => n3326, CK => CLK, Q => n11049, QN 
                           => n_1855);
   clk_r_REG1195_S1 : DFF_X1 port map( D => n3325, CK => CLK, Q => n11048, QN 
                           => n_1856);
   clk_r_REG1197_S1 : DFF_X1 port map( D => n3317, CK => CLK, Q => n11047, QN 
                           => n_1857);
   clk_r_REG1199_S1 : DFF_X1 port map( D => n3318, CK => CLK, Q => n11046, QN 
                           => n_1858);
   clk_r_REG1201_S1 : DFF_X1 port map( D => n3319, CK => CLK, Q => n11045, QN 
                           => n_1859);
   clk_r_REG1203_S1 : DFF_X1 port map( D => n3320, CK => CLK, Q => n11044, QN 
                           => n_1860);
   clk_r_REG1205_S1 : DFF_X1 port map( D => n3321, CK => CLK, Q => n11043, QN 
                           => n_1861);
   clk_r_REG1207_S1 : DFF_X1 port map( D => n3322, CK => CLK, Q => n11042, QN 
                           => n_1862);
   clk_r_REG1209_S1 : DFF_X1 port map( D => n3323, CK => CLK, Q => n11041, QN 
                           => n_1863);
   clk_r_REG1211_S1 : DFF_X1 port map( D => n3324, CK => CLK, Q => n11040, QN 
                           => n_1864);
   clk_r_REG1169_S1 : DFF_X1 port map( D => n3338, CK => CLK, Q => n11039, QN 
                           => n_1865);
   clk_r_REG1171_S1 : DFF_X1 port map( D => n3337, CK => CLK, Q => n11038, QN 
                           => n_1866);
   clk_r_REG1173_S1 : DFF_X1 port map( D => n3336, CK => CLK, Q => n11037, QN 
                           => n_1867);
   clk_r_REG1175_S1 : DFF_X1 port map( D => n3335, CK => CLK, Q => n11036, QN 
                           => n_1868);
   clk_r_REG1177_S1 : DFF_X1 port map( D => n3334, CK => CLK, Q => n11035, QN 
                           => n_1869);
   clk_r_REG1179_S1 : DFF_X1 port map( D => n3333, CK => CLK, Q => n11034, QN 
                           => n_1870);
   clk_r_REG1181_S1 : DFF_X1 port map( D => n3332, CK => CLK, Q => n11033, QN 
                           => n_1871);
   clk_r_REG1183_S1 : DFF_X1 port map( D => n3331, CK => CLK, Q => n11032, QN 
                           => n_1872);
   clk_r_REG1185_S1 : DFF_X1 port map( D => n3330, CK => CLK, Q => n11031, QN 
                           => n_1873);
   clk_r_REG1187_S1 : DFF_X1 port map( D => n3329, CK => CLK, Q => n11030, QN 
                           => n_1874);
   clk_r_REG1189_S1 : DFF_X1 port map( D => n3328, CK => CLK, Q => n11029, QN 
                           => n_1875);
   clk_r_REG386_S1 : DFF_X1 port map( D => n3348, CK => CLK, Q => n11028, QN =>
                           n_1876);
   clk_r_REG1151_S1 : DFF_X1 port map( D => n3347, CK => CLK, Q => n11027, QN 
                           => n_1877);
   clk_r_REG1153_S1 : DFF_X1 port map( D => n3346, CK => CLK, Q => n11026, QN 
                           => n_1878);
   clk_r_REG1155_S1 : DFF_X1 port map( D => n3345, CK => CLK, Q => n11025, QN 
                           => n_1879);
   clk_r_REG1157_S1 : DFF_X1 port map( D => n3344, CK => CLK, Q => n11024, QN 
                           => n_1880);
   clk_r_REG1159_S1 : DFF_X1 port map( D => n3343, CK => CLK, Q => n11023, QN 
                           => n_1881);
   clk_r_REG1161_S1 : DFF_X1 port map( D => n3342, CK => CLK, Q => n11022, QN 
                           => n_1882);
   clk_r_REG1163_S1 : DFF_X1 port map( D => n3341, CK => CLK, Q => n11021, QN 
                           => n_1883);
   clk_r_REG1165_S1 : DFF_X1 port map( D => n3340, CK => CLK, Q => n11020, QN 
                           => n_1884);
   clk_r_REG1167_S1 : DFF_X1 port map( D => n3339, CK => CLK, Q => n11019, QN 
                           => n_1885);
   clk_r_REG880_S1 : DFF_X1 port map( D => n3294, CK => CLK, Q => n11018, QN =>
                           n_1886);
   clk_r_REG882_S1 : DFF_X1 port map( D => n3293, CK => CLK, Q => n11017, QN =>
                           n_1887);
   clk_r_REG884_S1 : DFF_X1 port map( D => n3285, CK => CLK, Q => n11016, QN =>
                           n_1888);
   clk_r_REG886_S1 : DFF_X1 port map( D => n3286, CK => CLK, Q => n11015, QN =>
                           n_1889);
   clk_r_REG888_S1 : DFF_X1 port map( D => n3287, CK => CLK, Q => n11014, QN =>
                           n_1890);
   clk_r_REG890_S1 : DFF_X1 port map( D => n3288, CK => CLK, Q => n11013, QN =>
                           n_1891);
   clk_r_REG892_S1 : DFF_X1 port map( D => n3289, CK => CLK, Q => n11012, QN =>
                           n_1892);
   clk_r_REG894_S1 : DFF_X1 port map( D => n3290, CK => CLK, Q => n11011, QN =>
                           n_1893);
   clk_r_REG896_S1 : DFF_X1 port map( D => n3291, CK => CLK, Q => n11010, QN =>
                           n_1894);
   clk_r_REG898_S1 : DFF_X1 port map( D => n3292, CK => CLK, Q => n11009, QN =>
                           n_1895);
   clk_r_REG858_S1 : DFF_X1 port map( D => n3305, CK => CLK, Q => n11008, QN =>
                           n_1896);
   clk_r_REG860_S1 : DFF_X1 port map( D => n3304, CK => CLK, Q => n11007, QN =>
                           n_1897);
   clk_r_REG862_S1 : DFF_X1 port map( D => n3303, CK => CLK, Q => n11006, QN =>
                           n_1898);
   clk_r_REG864_S1 : DFF_X1 port map( D => n3302, CK => CLK, Q => n11005, QN =>
                           n_1899);
   clk_r_REG866_S1 : DFF_X1 port map( D => n3301, CK => CLK, Q => n11004, QN =>
                           n_1900);
   clk_r_REG868_S1 : DFF_X1 port map( D => n3300, CK => CLK, Q => n11003, QN =>
                           n_1901);
   clk_r_REG870_S1 : DFF_X1 port map( D => n3299, CK => CLK, Q => n11002, QN =>
                           n_1902);
   clk_r_REG872_S1 : DFF_X1 port map( D => n3298, CK => CLK, Q => n11001, QN =>
                           n_1903);
   clk_r_REG874_S1 : DFF_X1 port map( D => n3297, CK => CLK, Q => n11000, QN =>
                           n_1904);
   clk_r_REG876_S1 : DFF_X1 port map( D => n3296, CK => CLK, Q => n10999, QN =>
                           n_1905);
   clk_r_REG878_S1 : DFF_X1 port map( D => n3295, CK => CLK, Q => n10998, QN =>
                           n_1906);
   clk_r_REG825_S1 : DFF_X1 port map( D => n3316, CK => CLK, Q => n10997, QN =>
                           n_1907);
   clk_r_REG838_S1 : DFF_X1 port map( D => n3315, CK => CLK, Q => n10996, QN =>
                           n_1908);
   clk_r_REG840_S1 : DFF_X1 port map( D => n3314, CK => CLK, Q => n10995, QN =>
                           n_1909);
   clk_r_REG842_S1 : DFF_X1 port map( D => n3313, CK => CLK, Q => n10994, QN =>
                           n_1910);
   clk_r_REG844_S1 : DFF_X1 port map( D => n3312, CK => CLK, Q => n10993, QN =>
                           n_1911);
   clk_r_REG846_S1 : DFF_X1 port map( D => n3311, CK => CLK, Q => n10992, QN =>
                           n_1912);
   clk_r_REG848_S1 : DFF_X1 port map( D => n3310, CK => CLK, Q => n10991, QN =>
                           n_1913);
   clk_r_REG850_S1 : DFF_X1 port map( D => n3309, CK => CLK, Q => n10990, QN =>
                           n_1914);
   clk_r_REG852_S1 : DFF_X1 port map( D => n3308, CK => CLK, Q => n10989, QN =>
                           n_1915);
   clk_r_REG854_S1 : DFF_X1 port map( D => n3307, CK => CLK, Q => n10988, QN =>
                           n_1916);
   clk_r_REG856_S1 : DFF_X1 port map( D => n3306, CK => CLK, Q => n10987, QN =>
                           n_1917);
   clk_r_REG805_S1 : DFF_X1 port map( D => n3261, CK => CLK, Q => n10986, QN =>
                           n_1918);
   clk_r_REG807_S1 : DFF_X1 port map( D => n3253, CK => CLK, Q => n10985, QN =>
                           n_1919);
   clk_r_REG809_S1 : DFF_X1 port map( D => n3254, CK => CLK, Q => n10984, QN =>
                           n_1920);
   clk_r_REG811_S1 : DFF_X1 port map( D => n3255, CK => CLK, Q => n10983, QN =>
                           n_1921);
   clk_r_REG813_S1 : DFF_X1 port map( D => n3256, CK => CLK, Q => n10982, QN =>
                           n_1922);
   clk_r_REG815_S1 : DFF_X1 port map( D => n3257, CK => CLK, Q => n10981, QN =>
                           n_1923);
   clk_r_REG817_S1 : DFF_X1 port map( D => n3258, CK => CLK, Q => n10980, QN =>
                           n_1924);
   clk_r_REG819_S1 : DFF_X1 port map( D => n3259, CK => CLK, Q => n10979, QN =>
                           n_1925);
   clk_r_REG821_S1 : DFF_X1 port map( D => n3260, CK => CLK, Q => n10978, QN =>
                           n_1926);
   clk_r_REG783_S1 : DFF_X1 port map( D => n3272, CK => CLK, Q => n10977, QN =>
                           n_1927);
   clk_r_REG785_S1 : DFF_X1 port map( D => n3271, CK => CLK, Q => n10976, QN =>
                           n_1928);
   clk_r_REG787_S1 : DFF_X1 port map( D => n3270, CK => CLK, Q => n10975, QN =>
                           n_1929);
   clk_r_REG789_S1 : DFF_X1 port map( D => n3269, CK => CLK, Q => n10974, QN =>
                           n_1930);
   clk_r_REG791_S1 : DFF_X1 port map( D => n3268, CK => CLK, Q => n10973, QN =>
                           n_1931);
   clk_r_REG793_S1 : DFF_X1 port map( D => n3267, CK => CLK, Q => n10972, QN =>
                           n_1932);
   clk_r_REG795_S1 : DFF_X1 port map( D => n3266, CK => CLK, Q => n10971, QN =>
                           n_1933);
   clk_r_REG797_S1 : DFF_X1 port map( D => n3265, CK => CLK, Q => n10970, QN =>
                           n_1934);
   clk_r_REG799_S1 : DFF_X1 port map( D => n3264, CK => CLK, Q => n10969, QN =>
                           n_1935);
   clk_r_REG801_S1 : DFF_X1 port map( D => n3263, CK => CLK, Q => n10968, QN =>
                           n_1936);
   clk_r_REG803_S1 : DFF_X1 port map( D => n3262, CK => CLK, Q => n10967, QN =>
                           n_1937);
   clk_r_REG761_S1 : DFF_X1 port map( D => n3283, CK => CLK, Q => n10966, QN =>
                           n_1938);
   clk_r_REG763_S1 : DFF_X1 port map( D => n3282, CK => CLK, Q => n10965, QN =>
                           n_1939);
   clk_r_REG765_S1 : DFF_X1 port map( D => n3281, CK => CLK, Q => n10964, QN =>
                           n_1940);
   clk_r_REG767_S1 : DFF_X1 port map( D => n3280, CK => CLK, Q => n10963, QN =>
                           n_1941);
   clk_r_REG769_S1 : DFF_X1 port map( D => n3279, CK => CLK, Q => n10962, QN =>
                           n_1942);
   clk_r_REG771_S1 : DFF_X1 port map( D => n3278, CK => CLK, Q => n10961, QN =>
                           n_1943);
   clk_r_REG773_S1 : DFF_X1 port map( D => n3277, CK => CLK, Q => n10960, QN =>
                           n_1944);
   clk_r_REG775_S1 : DFF_X1 port map( D => n3276, CK => CLK, Q => n10959, QN =>
                           n_1945);
   clk_r_REG777_S1 : DFF_X1 port map( D => n3275, CK => CLK, Q => n10958, QN =>
                           n_1946);
   clk_r_REG779_S1 : DFF_X1 port map( D => n3274, CK => CLK, Q => n10957, QN =>
                           n_1947);
   clk_r_REG781_S1 : DFF_X1 port map( D => n3273, CK => CLK, Q => n10956, QN =>
                           n_1948);
   clk_r_REG1133_S1 : DFF_X1 port map( D => n3221, CK => CLK, Q => n10955, QN 
                           => n_1949);
   clk_r_REG1135_S1 : DFF_X1 port map( D => n3222, CK => CLK, Q => n10954, QN 
                           => n_1950);
   clk_r_REG1137_S1 : DFF_X1 port map( D => n3223, CK => CLK, Q => n10953, QN 
                           => n_1951);
   clk_r_REG1139_S1 : DFF_X1 port map( D => n3224, CK => CLK, Q => n10952, QN 
                           => n_1952);
   clk_r_REG1141_S1 : DFF_X1 port map( D => n3225, CK => CLK, Q => n10951, QN 
                           => n_1953);
   clk_r_REG1143_S1 : DFF_X1 port map( D => n3226, CK => CLK, Q => n10950, QN 
                           => n_1954);
   clk_r_REG1145_S1 : DFF_X1 port map( D => n3227, CK => CLK, Q => n10949, QN 
                           => n_1955);
   clk_r_REG1147_S1 : DFF_X1 port map( D => n3228, CK => CLK, Q => n10948, QN 
                           => n_1956);
   clk_r_REG747_S1 : DFF_X1 port map( D => n3284, CK => CLK, Q => n10947, QN =>
                           n_1957);
   clk_r_REG1111_S1 : DFF_X1 port map( D => n3239, CK => CLK, Q => n10946, QN 
                           => n_1958);
   clk_r_REG1113_S1 : DFF_X1 port map( D => n3238, CK => CLK, Q => n10945, QN 
                           => n_1959);
   clk_r_REG1115_S1 : DFF_X1 port map( D => n3237, CK => CLK, Q => n10944, QN 
                           => n_1960);
   clk_r_REG1117_S1 : DFF_X1 port map( D => n3236, CK => CLK, Q => n10943, QN 
                           => n_1961);
   clk_r_REG1119_S1 : DFF_X1 port map( D => n3235, CK => CLK, Q => n10942, QN 
                           => n_1962);
   clk_r_REG1121_S1 : DFF_X1 port map( D => n3234, CK => CLK, Q => n10941, QN 
                           => n_1963);
   clk_r_REG1123_S1 : DFF_X1 port map( D => n3233, CK => CLK, Q => n10940, QN 
                           => n_1964);
   clk_r_REG1125_S1 : DFF_X1 port map( D => n3232, CK => CLK, Q => n10939, QN 
                           => n_1965);
   clk_r_REG1127_S1 : DFF_X1 port map( D => n3231, CK => CLK, Q => n10938, QN 
                           => n_1966);
   clk_r_REG1129_S1 : DFF_X1 port map( D => n3230, CK => CLK, Q => n10937, QN 
                           => n_1967);
   clk_r_REG1131_S1 : DFF_X1 port map( D => n3229, CK => CLK, Q => n10936, QN 
                           => n_1968);
   clk_r_REG1089_S1 : DFF_X1 port map( D => n3250, CK => CLK, Q => n10935, QN 
                           => n_1969);
   clk_r_REG1091_S1 : DFF_X1 port map( D => n3249, CK => CLK, Q => n10934, QN 
                           => n_1970);
   clk_r_REG1093_S1 : DFF_X1 port map( D => n3248, CK => CLK, Q => n10933, QN 
                           => n_1971);
   clk_r_REG1095_S1 : DFF_X1 port map( D => n3247, CK => CLK, Q => n10932, QN 
                           => n_1972);
   clk_r_REG1097_S1 : DFF_X1 port map( D => n3246, CK => CLK, Q => n10931, QN 
                           => n_1973);
   clk_r_REG1099_S1 : DFF_X1 port map( D => n3245, CK => CLK, Q => n10930, QN 
                           => n_1974);
   clk_r_REG1101_S1 : DFF_X1 port map( D => n3244, CK => CLK, Q => n10929, QN 
                           => n_1975);
   clk_r_REG1103_S1 : DFF_X1 port map( D => n3243, CK => CLK, Q => n10928, QN 
                           => n_1976);
   clk_r_REG1105_S1 : DFF_X1 port map( D => n3242, CK => CLK, Q => n10927, QN 
                           => n_1977);
   clk_r_REG1107_S1 : DFF_X1 port map( D => n3241, CK => CLK, Q => n10926, QN 
                           => n_1978);
   clk_r_REG1109_S1 : DFF_X1 port map( D => n3240, CK => CLK, Q => n10925, QN 
                           => n_1979);
   clk_r_REG1060_S1 : DFF_X1 port map( D => n3190, CK => CLK, Q => n10924, QN 
                           => n_1980);
   clk_r_REG1062_S1 : DFF_X1 port map( D => n3191, CK => CLK, Q => n10923, QN 
                           => n_1981);
   clk_r_REG1064_S1 : DFF_X1 port map( D => n3192, CK => CLK, Q => n10922, QN 
                           => n_1982);
   clk_r_REG1066_S1 : DFF_X1 port map( D => n3193, CK => CLK, Q => n10921, QN 
                           => n_1983);
   clk_r_REG1068_S1 : DFF_X1 port map( D => n3194, CK => CLK, Q => n10920, QN 
                           => n_1984);
   clk_r_REG1070_S1 : DFF_X1 port map( D => n3195, CK => CLK, Q => n10919, QN 
                           => n_1985);
   clk_r_REG1072_S1 : DFF_X1 port map( D => n3196, CK => CLK, Q => n10918, QN 
                           => n_1986);
   clk_r_REG1076_S1 : DFF_X1 port map( D => n3252, CK => CLK, Q => n10917, QN 
                           => n_1987);
   clk_r_REG1087_S1 : DFF_X1 port map( D => n3251, CK => CLK, Q => n10916, QN 
                           => n_1988);
   clk_r_REG1038_S1 : DFF_X1 port map( D => n3206, CK => CLK, Q => n10915, QN 
                           => n_1989);
   clk_r_REG1040_S1 : DFF_X1 port map( D => n3205, CK => CLK, Q => n10914, QN 
                           => n_1990);
   clk_r_REG1042_S1 : DFF_X1 port map( D => n3204, CK => CLK, Q => n10913, QN 
                           => n_1991);
   clk_r_REG1044_S1 : DFF_X1 port map( D => n3203, CK => CLK, Q => n10912, QN 
                           => n_1992);
   clk_r_REG1046_S1 : DFF_X1 port map( D => n3202, CK => CLK, Q => n10911, QN 
                           => n_1993);
   clk_r_REG1048_S1 : DFF_X1 port map( D => n3201, CK => CLK, Q => n10910, QN 
                           => n_1994);
   clk_r_REG1050_S1 : DFF_X1 port map( D => n3200, CK => CLK, Q => n10909, QN 
                           => n_1995);
   clk_r_REG1052_S1 : DFF_X1 port map( D => n3199, CK => CLK, Q => n10908, QN 
                           => n_1996);
   clk_r_REG1054_S1 : DFF_X1 port map( D => n3198, CK => CLK, Q => n10907, QN 
                           => n_1997);
   clk_r_REG1056_S1 : DFF_X1 port map( D => n3197, CK => CLK, Q => n10906, QN 
                           => n_1998);
   clk_r_REG1058_S1 : DFF_X1 port map( D => n3189, CK => CLK, Q => n10905, QN 
                           => n_1999);
   clk_r_REG1016_S1 : DFF_X1 port map( D => n3217, CK => CLK, Q => n10904, QN 
                           => n_2000);
   clk_r_REG1018_S1 : DFF_X1 port map( D => n3216, CK => CLK, Q => n10903, QN 
                           => n_2001);
   clk_r_REG1020_S1 : DFF_X1 port map( D => n3215, CK => CLK, Q => n10902, QN 
                           => n_2002);
   clk_r_REG1022_S1 : DFF_X1 port map( D => n3214, CK => CLK, Q => n10901, QN 
                           => n_2003);
   clk_r_REG1024_S1 : DFF_X1 port map( D => n3213, CK => CLK, Q => n10900, QN 
                           => n_2004);
   clk_r_REG1026_S1 : DFF_X1 port map( D => n3212, CK => CLK, Q => n10899, QN 
                           => n_2005);
   clk_r_REG1028_S1 : DFF_X1 port map( D => n3211, CK => CLK, Q => n10898, QN 
                           => n_2006);
   clk_r_REG1030_S1 : DFF_X1 port map( D => n3210, CK => CLK, Q => n10897, QN 
                           => n_2007);
   clk_r_REG1032_S1 : DFF_X1 port map( D => n3209, CK => CLK, Q => n10896, QN 
                           => n_2008);
   clk_r_REG1034_S1 : DFF_X1 port map( D => n3208, CK => CLK, Q => n10895, QN 
                           => n_2009);
   clk_r_REG1036_S1 : DFF_X1 port map( D => n3207, CK => CLK, Q => n10894, QN 
                           => n_2010);
   clk_r_REG1783_S1 : DFF_X1 port map( D => n3159, CK => CLK, Q => n10893, QN 
                           => n_2011);
   clk_r_REG1785_S1 : DFF_X1 port map( D => n3160, CK => CLK, Q => n10892, QN 
                           => n_2012);
   clk_r_REG1787_S1 : DFF_X1 port map( D => n3161, CK => CLK, Q => n10891, QN 
                           => n_2013);
   clk_r_REG1789_S1 : DFF_X1 port map( D => n3162, CK => CLK, Q => n10890, QN 
                           => n_2014);
   clk_r_REG1791_S1 : DFF_X1 port map( D => n3163, CK => CLK, Q => n10889, QN 
                           => n_2015);
   clk_r_REG1793_S1 : DFF_X1 port map( D => n3164, CK => CLK, Q => n10888, QN 
                           => n_2016);
   clk_r_REG1001_S1 : DFF_X1 port map( D => n3220, CK => CLK, Q => n10887, QN 
                           => n_2017);
   clk_r_REG1012_S1 : DFF_X1 port map( D => n3219, CK => CLK, Q => n10886, QN 
                           => n_2018);
   clk_r_REG1014_S1 : DFF_X1 port map( D => n3218, CK => CLK, Q => n10885, QN 
                           => n_2019);
   clk_r_REG1761_S1 : DFF_X1 port map( D => n3173, CK => CLK, Q => n10884, QN 
                           => n_2020);
   clk_r_REG1763_S1 : DFF_X1 port map( D => n3172, CK => CLK, Q => n10883, QN 
                           => n_2021);
   clk_r_REG1765_S1 : DFF_X1 port map( D => n3171, CK => CLK, Q => n10882, QN 
                           => n_2022);
   clk_r_REG1767_S1 : DFF_X1 port map( D => n3170, CK => CLK, Q => n10881, QN 
                           => n_2023);
   clk_r_REG1769_S1 : DFF_X1 port map( D => n3169, CK => CLK, Q => n10880, QN 
                           => n_2024);
   clk_r_REG1771_S1 : DFF_X1 port map( D => n3168, CK => CLK, Q => n10879, QN 
                           => n_2025);
   clk_r_REG1773_S1 : DFF_X1 port map( D => n3167, CK => CLK, Q => n10878, QN 
                           => n_2026);
   clk_r_REG1775_S1 : DFF_X1 port map( D => n3166, CK => CLK, Q => n10877, QN 
                           => n_2027);
   clk_r_REG1777_S1 : DFF_X1 port map( D => n3165, CK => CLK, Q => n10876, QN 
                           => n_2028);
   clk_r_REG1779_S1 : DFF_X1 port map( D => n3157, CK => CLK, Q => n10875, QN 
                           => n_2029);
   clk_r_REG1781_S1 : DFF_X1 port map( D => n3158, CK => CLK, Q => n10874, QN 
                           => n_2030);
   clk_r_REG1739_S1 : DFF_X1 port map( D => n3184, CK => CLK, Q => n10873, QN 
                           => n_2031);
   clk_r_REG1741_S1 : DFF_X1 port map( D => n3183, CK => CLK, Q => n10872, QN 
                           => n_2032);
   clk_r_REG1743_S1 : DFF_X1 port map( D => n3182, CK => CLK, Q => n10871, QN 
                           => n_2033);
   clk_r_REG1745_S1 : DFF_X1 port map( D => n3181, CK => CLK, Q => n10870, QN 
                           => n_2034);
   clk_r_REG1747_S1 : DFF_X1 port map( D => n3180, CK => CLK, Q => n10869, QN 
                           => n_2035);
   clk_r_REG1749_S1 : DFF_X1 port map( D => n3179, CK => CLK, Q => n10868, QN 
                           => n_2036);
   clk_r_REG1751_S1 : DFF_X1 port map( D => n3178, CK => CLK, Q => n10867, QN 
                           => n_2037);
   clk_r_REG1753_S1 : DFF_X1 port map( D => n3177, CK => CLK, Q => n10866, QN 
                           => n_2038);
   clk_r_REG1755_S1 : DFF_X1 port map( D => n3176, CK => CLK, Q => n10865, QN 
                           => n_2039);
   clk_r_REG1757_S1 : DFF_X1 port map( D => n3175, CK => CLK, Q => n10864, QN 
                           => n_2040);
   clk_r_REG1759_S1 : DFF_X1 port map( D => n3174, CK => CLK, Q => n10863, QN 
                           => n_2041);
   clk_r_REG1448_S1 : DFF_X1 port map( D => n3128, CK => CLK, Q => n10862, QN 
                           => n_2042);
   clk_r_REG1450_S1 : DFF_X1 port map( D => n3129, CK => CLK, Q => n10861, QN 
                           => n_2043);
   clk_r_REG1452_S1 : DFF_X1 port map( D => n3130, CK => CLK, Q => n10860, QN 
                           => n_2044);
   clk_r_REG1454_S1 : DFF_X1 port map( D => n3131, CK => CLK, Q => n10859, QN 
                           => n_2045);
   clk_r_REG1456_S1 : DFF_X1 port map( D => n3132, CK => CLK, Q => n10858, QN 
                           => n_2046);
   clk_r_REG1722_S1 : DFF_X1 port map( D => n3188, CK => CLK, Q => n10857, QN 
                           => n_2047);
   clk_r_REG1733_S1 : DFF_X1 port map( D => n3187, CK => CLK, Q => n10856, QN 
                           => n_2048);
   clk_r_REG1735_S1 : DFF_X1 port map( D => n3186, CK => CLK, Q => n10855, QN 
                           => n_2049);
   clk_r_REG1737_S1 : DFF_X1 port map( D => n3185, CK => CLK, Q => n10854, QN 
                           => n_2050);
   clk_r_REG1426_S1 : DFF_X1 port map( D => n3140, CK => CLK, Q => n10853, QN 
                           => n_2051);
   clk_r_REG1428_S1 : DFF_X1 port map( D => n3139, CK => CLK, Q => n10852, QN 
                           => n_2052);
   clk_r_REG1430_S1 : DFF_X1 port map( D => n3138, CK => CLK, Q => n10851, QN 
                           => n_2053);
   clk_r_REG1432_S1 : DFF_X1 port map( D => n3137, CK => CLK, Q => n10850, QN 
                           => n_2054);
   clk_r_REG1434_S1 : DFF_X1 port map( D => n3136, CK => CLK, Q => n10849, QN 
                           => n_2055);
   clk_r_REG1436_S1 : DFF_X1 port map( D => n3135, CK => CLK, Q => n10848, QN 
                           => n_2056);
   clk_r_REG1438_S1 : DFF_X1 port map( D => n3134, CK => CLK, Q => n10847, QN 
                           => n_2057);
   clk_r_REG1440_S1 : DFF_X1 port map( D => n3133, CK => CLK, Q => n10846, QN 
                           => n_2058);
   clk_r_REG1442_S1 : DFF_X1 port map( D => n3125, CK => CLK, Q => n10845, QN 
                           => n_2059);
   clk_r_REG1444_S1 : DFF_X1 port map( D => n3126, CK => CLK, Q => n10844, QN 
                           => n_2060);
   clk_r_REG1446_S1 : DFF_X1 port map( D => n3127, CK => CLK, Q => n10843, QN 
                           => n_2061);
   clk_r_REG1404_S1 : DFF_X1 port map( D => n3151, CK => CLK, Q => n10842, QN 
                           => n_2062);
   clk_r_REG1406_S1 : DFF_X1 port map( D => n3150, CK => CLK, Q => n10841, QN 
                           => n_2063);
   clk_r_REG1408_S1 : DFF_X1 port map( D => n3149, CK => CLK, Q => n10840, QN 
                           => n_2064);
   clk_r_REG1410_S1 : DFF_X1 port map( D => n3148, CK => CLK, Q => n10839, QN 
                           => n_2065);
   clk_r_REG1412_S1 : DFF_X1 port map( D => n3147, CK => CLK, Q => n10838, QN 
                           => n_2066);
   clk_r_REG1414_S1 : DFF_X1 port map( D => n3146, CK => CLK, Q => n10837, QN 
                           => n_2067);
   clk_r_REG1416_S1 : DFF_X1 port map( D => n3145, CK => CLK, Q => n10836, QN 
                           => n_2068);
   clk_r_REG1418_S1 : DFF_X1 port map( D => n3144, CK => CLK, Q => n10835, QN 
                           => n_2069);
   clk_r_REG1420_S1 : DFF_X1 port map( D => n3143, CK => CLK, Q => n10834, QN 
                           => n_2070);
   clk_r_REG1422_S1 : DFF_X1 port map( D => n3142, CK => CLK, Q => n10833, QN 
                           => n_2071);
   clk_r_REG1424_S1 : DFF_X1 port map( D => n3141, CK => CLK, Q => n10832, QN 
                           => n_2072);
   clk_r_REG1626_S1 : DFF_X1 port map( D => n3065, CK => CLK, Q => n10831, QN 
                           => n_2073);
   clk_r_REG1628_S1 : DFF_X1 port map( D => n3066, CK => CLK, Q => n10830, QN 
                           => n_2074);
   clk_r_REG1630_S1 : DFF_X1 port map( D => n3067, CK => CLK, Q => n10829, QN 
                           => n_2075);
   clk_r_REG1632_S1 : DFF_X1 port map( D => n3068, CK => CLK, Q => n10828, QN 
                           => n_2076);
   clk_r_REG1382_S1 : DFF_X1 port map( D => n3156, CK => CLK, Q => n10827, QN 
                           => n_2077);
   clk_r_REG1396_S1 : DFF_X1 port map( D => n3155, CK => CLK, Q => n10826, QN 
                           => n_2078);
   clk_r_REG1398_S1 : DFF_X1 port map( D => n3154, CK => CLK, Q => n10825, QN 
                           => n_2079);
   clk_r_REG1400_S1 : DFF_X1 port map( D => n3153, CK => CLK, Q => n10824, QN 
                           => n_2080);
   clk_r_REG1402_S1 : DFF_X1 port map( D => n3152, CK => CLK, Q => n10823, QN 
                           => n_2081);
   clk_r_REG1604_S1 : DFF_X1 port map( D => n3075, CK => CLK, Q => n10822, QN 
                           => n_2082);
   clk_r_REG1606_S1 : DFF_X1 port map( D => n3074, CK => CLK, Q => n10821, QN 
                           => n_2083);
   clk_r_REG1608_S1 : DFF_X1 port map( D => n3073, CK => CLK, Q => n10820, QN 
                           => n_2084);
   clk_r_REG1610_S1 : DFF_X1 port map( D => n3072, CK => CLK, Q => n10819, QN 
                           => n_2085);
   clk_r_REG1612_S1 : DFF_X1 port map( D => n3071, CK => CLK, Q => n10818, QN 
                           => n_2086);
   clk_r_REG1614_S1 : DFF_X1 port map( D => n3070, CK => CLK, Q => n10817, QN 
                           => n_2087);
   clk_r_REG1616_S1 : DFF_X1 port map( D => n3069, CK => CLK, Q => n10816, QN 
                           => n_2088);
   clk_r_REG1618_S1 : DFF_X1 port map( D => n3061, CK => CLK, Q => n10815, QN 
                           => n_2089);
   clk_r_REG1620_S1 : DFF_X1 port map( D => n3062, CK => CLK, Q => n10814, QN 
                           => n_2090);
   clk_r_REG1622_S1 : DFF_X1 port map( D => n3063, CK => CLK, Q => n10813, QN 
                           => n_2091);
   clk_r_REG1624_S1 : DFF_X1 port map( D => n3064, CK => CLK, Q => n10812, QN 
                           => n_2092);
   clk_r_REG1582_S1 : DFF_X1 port map( D => n3086, CK => CLK, Q => n10811, QN 
                           => n_2093);
   clk_r_REG1584_S1 : DFF_X1 port map( D => n3085, CK => CLK, Q => n10810, QN 
                           => n_2094);
   clk_r_REG1586_S1 : DFF_X1 port map( D => n3084, CK => CLK, Q => n10809, QN 
                           => n_2095);
   clk_r_REG1588_S1 : DFF_X1 port map( D => n3083, CK => CLK, Q => n10808, QN 
                           => n_2096);
   clk_r_REG1590_S1 : DFF_X1 port map( D => n3082, CK => CLK, Q => n10807, QN 
                           => n_2097);
   clk_r_REG1592_S1 : DFF_X1 port map( D => n3081, CK => CLK, Q => n10806, QN 
                           => n_2098);
   clk_r_REG1594_S1 : DFF_X1 port map( D => n3080, CK => CLK, Q => n10805, QN 
                           => n_2099);
   clk_r_REG1596_S1 : DFF_X1 port map( D => n3079, CK => CLK, Q => n10804, QN 
                           => n_2100);
   clk_r_REG1598_S1 : DFF_X1 port map( D => n3078, CK => CLK, Q => n10803, QN 
                           => n_2101);
   clk_r_REG1600_S1 : DFF_X1 port map( D => n3077, CK => CLK, Q => n10802, QN 
                           => n_2102);
   clk_r_REG1602_S1 : DFF_X1 port map( D => n3076, CK => CLK, Q => n10801, QN 
                           => n_2103);
   clk_r_REG1705_S1 : DFF_X1 port map( D => n3098, CK => CLK, Q => n10800, QN 
                           => n_2104);
   clk_r_REG1707_S1 : DFF_X1 port map( D => n3099, CK => CLK, Q => n10799, QN 
                           => n_2105);
   clk_r_REG1560_S1 : DFF_X1 port map( D => n3092, CK => CLK, Q => n10798, QN 
                           => n_2106);
   clk_r_REG1572_S1 : DFF_X1 port map( D => n3091, CK => CLK, Q => n10797, QN 
                           => n_2107);
   clk_r_REG1574_S1 : DFF_X1 port map( D => n3090, CK => CLK, Q => n10796, QN 
                           => n_2108);
   clk_r_REG1576_S1 : DFF_X1 port map( D => n3089, CK => CLK, Q => n10795, QN 
                           => n_2109);
   clk_r_REG1578_S1 : DFF_X1 port map( D => n3088, CK => CLK, Q => n10794, QN 
                           => n_2110);
   clk_r_REG1580_S1 : DFF_X1 port map( D => n3087, CK => CLK, Q => n10793, QN 
                           => n_2111);
   clk_r_REG1683_S1 : DFF_X1 port map( D => n3106, CK => CLK, Q => n10792, QN 
                           => n_2112);
   clk_r_REG1685_S1 : DFF_X1 port map( D => n3105, CK => CLK, Q => n10791, QN 
                           => n_2113);
   clk_r_REG1687_S1 : DFF_X1 port map( D => n3104, CK => CLK, Q => n10790, QN 
                           => n_2114);
   clk_r_REG1689_S1 : DFF_X1 port map( D => n3103, CK => CLK, Q => n10789, QN 
                           => n_2115);
   clk_r_REG1691_S1 : DFF_X1 port map( D => n3102, CK => CLK, Q => n10788, QN 
                           => n_2116);
   clk_r_REG1693_S1 : DFF_X1 port map( D => n3101, CK => CLK, Q => n10787, QN 
                           => n_2117);
   clk_r_REG1695_S1 : DFF_X1 port map( D => n3093, CK => CLK, Q => n10786, QN 
                           => n_2118);
   clk_r_REG1697_S1 : DFF_X1 port map( D => n3094, CK => CLK, Q => n10785, QN 
                           => n_2119);
   clk_r_REG1699_S1 : DFF_X1 port map( D => n3095, CK => CLK, Q => n10784, QN 
                           => n_2120);
   clk_r_REG1701_S1 : DFF_X1 port map( D => n3096, CK => CLK, Q => n10783, QN 
                           => n_2121);
   clk_r_REG1703_S1 : DFF_X1 port map( D => n3097, CK => CLK, Q => n10782, QN 
                           => n_2122);
   clk_r_REG1661_S1 : DFF_X1 port map( D => n3117, CK => CLK, Q => n10781, QN 
                           => n_2123);
   clk_r_REG1663_S1 : DFF_X1 port map( D => n3116, CK => CLK, Q => n10780, QN 
                           => n_2124);
   clk_r_REG1665_S1 : DFF_X1 port map( D => n3115, CK => CLK, Q => n10779, QN 
                           => n_2125);
   clk_r_REG1667_S1 : DFF_X1 port map( D => n3114, CK => CLK, Q => n10778, QN 
                           => n_2126);
   clk_r_REG1669_S1 : DFF_X1 port map( D => n3113, CK => CLK, Q => n10777, QN 
                           => n_2127);
   clk_r_REG1671_S1 : DFF_X1 port map( D => n3112, CK => CLK, Q => n10776, QN 
                           => n_2128);
   clk_r_REG1673_S1 : DFF_X1 port map( D => n3111, CK => CLK, Q => n10775, QN 
                           => n_2129);
   clk_r_REG1675_S1 : DFF_X1 port map( D => n3110, CK => CLK, Q => n10774, QN 
                           => n_2130);
   clk_r_REG1677_S1 : DFF_X1 port map( D => n3109, CK => CLK, Q => n10773, QN 
                           => n_2131);
   clk_r_REG1679_S1 : DFF_X1 port map( D => n3108, CK => CLK, Q => n10772, QN 
                           => n_2132);
   clk_r_REG1681_S1 : DFF_X1 port map( D => n3107, CK => CLK, Q => n10771, QN 
                           => n_2133);
   clk_r_REG2785_S1 : DFF_X1 port map( D => n2906, CK => CLK, Q => n10770, QN 
                           => n_2134);
   clk_r_REG2787_S1 : DFF_X1 port map( D => n2907, CK => CLK, Q => n10769, QN 
                           => n_2135);
   clk_r_REG2789_S1 : DFF_X1 port map( D => n2908, CK => CLK, Q => n10768, QN 
                           => n_2136);
   clk_r_REG1636_S1 : DFF_X1 port map( D => n3124, CK => CLK, Q => n10767, QN 
                           => n_2137);
   clk_r_REG1649_S1 : DFF_X1 port map( D => n3123, CK => CLK, Q => n10766, QN 
                           => n_2138);
   clk_r_REG1651_S1 : DFF_X1 port map( D => n3122, CK => CLK, Q => n10765, QN 
                           => n_2139);
   clk_r_REG1653_S1 : DFF_X1 port map( D => n3121, CK => CLK, Q => n10764, QN 
                           => n_2140);
   clk_r_REG1655_S1 : DFF_X1 port map( D => n3120, CK => CLK, Q => n10763, QN 
                           => n_2141);
   clk_r_REG1657_S1 : DFF_X1 port map( D => n3119, CK => CLK, Q => n10762, QN 
                           => n_2142);
   clk_r_REG1659_S1 : DFF_X1 port map( D => n3118, CK => CLK, Q => n10761, QN 
                           => n_2143);
   clk_r_REG2763_S1 : DFF_X1 port map( D => n2914, CK => CLK, Q => n10760, QN 
                           => n_2144);
   clk_r_REG2765_S1 : DFF_X1 port map( D => n2913, CK => CLK, Q => n10759, QN 
                           => n_2145);
   clk_r_REG2767_S1 : DFF_X1 port map( D => n2912, CK => CLK, Q => n10758, QN 
                           => n_2146);
   clk_r_REG2769_S1 : DFF_X1 port map( D => n2911, CK => CLK, Q => n10757, QN 
                           => n_2147);
   clk_r_REG2771_S1 : DFF_X1 port map( D => n2910, CK => CLK, Q => n10756, QN 
                           => n_2148);
   clk_r_REG2773_S1 : DFF_X1 port map( D => n2909, CK => CLK, Q => n10755, QN 
                           => n_2149);
   clk_r_REG2775_S1 : DFF_X1 port map( D => n2901, CK => CLK, Q => n10754, QN 
                           => n_2150);
   clk_r_REG2777_S1 : DFF_X1 port map( D => n2902, CK => CLK, Q => n10753, QN 
                           => n_2151);
   clk_r_REG2779_S1 : DFF_X1 port map( D => n2903, CK => CLK, Q => n10752, QN 
                           => n_2152);
   clk_r_REG2781_S1 : DFF_X1 port map( D => n2904, CK => CLK, Q => n10751, QN 
                           => n_2153);
   clk_r_REG2783_S1 : DFF_X1 port map( D => n2905, CK => CLK, Q => n10750, QN 
                           => n_2154);
   clk_r_REG1372_S1 : DFF_X1 port map( D => n3449, CK => CLK, Q => n10749, QN 
                           => n_2155);
   clk_r_REG1374_S1 : DFF_X1 port map( D => n3450, CK => CLK, Q => n10748, QN 
                           => n_2156);
   clk_r_REG1376_S1 : DFF_X1 port map( D => n3451, CK => CLK, Q => n10747, QN 
                           => n_2157);
   clk_r_REG1378_S1 : DFF_X1 port map( D => n3452, CK => CLK, Q => n10746, QN 
                           => n_2158);
   clk_r_REG3039_S1 : DFF_X1 port map( D => n3540, CK => CLK, Q => n10745, QN 
                           => n_2159);
   clk_r_REG3045_S1 : DFF_X1 port map( D => n3539, CK => CLK, Q => n10744, QN 
                           => n_2160);
   clk_r_REG3047_S1 : DFF_X1 port map( D => n3538, CK => CLK, Q => n10743, QN 
                           => n_2161);
   clk_r_REG3049_S1 : DFF_X1 port map( D => n3537, CK => CLK, Q => n10742, QN 
                           => n_2162);
   clk_r_REG3051_S1 : DFF_X1 port map( D => n3536, CK => CLK, Q => n10741, QN 
                           => n_2163);
   clk_r_REG1350_S1 : DFF_X1 port map( D => n3459, CK => CLK, Q => n10740, QN 
                           => n_2164);
   clk_r_REG1352_S1 : DFF_X1 port map( D => n3458, CK => CLK, Q => n10739, QN 
                           => n_2165);
   clk_r_REG1354_S1 : DFF_X1 port map( D => n3457, CK => CLK, Q => n10738, QN 
                           => n_2166);
   clk_r_REG1356_S1 : DFF_X1 port map( D => n3456, CK => CLK, Q => n10737, QN 
                           => n_2167);
   clk_r_REG1358_S1 : DFF_X1 port map( D => n3455, CK => CLK, Q => n10736, QN 
                           => n_2168);
   clk_r_REG1360_S1 : DFF_X1 port map( D => n3454, CK => CLK, Q => n10735, QN 
                           => n_2169);
   clk_r_REG1362_S1 : DFF_X1 port map( D => n3453, CK => CLK, Q => n10734, QN 
                           => n_2170);
   clk_r_REG1364_S1 : DFF_X1 port map( D => n3445, CK => CLK, Q => n10733, QN 
                           => n_2171);
   clk_r_REG1366_S1 : DFF_X1 port map( D => n3446, CK => CLK, Q => n10732, QN 
                           => n_2172);
   clk_r_REG1368_S1 : DFF_X1 port map( D => n3447, CK => CLK, Q => n10731, QN 
                           => n_2173);
   clk_r_REG1370_S1 : DFF_X1 port map( D => n3448, CK => CLK, Q => n10730, QN 
                           => n_2174);
   clk_r_REG1328_S1 : DFF_X1 port map( D => n3470, CK => CLK, Q => n10729, QN 
                           => n_2175);
   clk_r_REG1330_S1 : DFF_X1 port map( D => n3469, CK => CLK, Q => n10728, QN 
                           => n_2176);
   clk_r_REG1332_S1 : DFF_X1 port map( D => n3468, CK => CLK, Q => n10727, QN 
                           => n_2177);
   clk_r_REG1334_S1 : DFF_X1 port map( D => n3467, CK => CLK, Q => n10726, QN 
                           => n_2178);
   clk_r_REG1336_S1 : DFF_X1 port map( D => n3466, CK => CLK, Q => n10725, QN 
                           => n_2179);
   clk_r_REG1338_S1 : DFF_X1 port map( D => n3465, CK => CLK, Q => n10724, QN 
                           => n_2180);
   clk_r_REG1340_S1 : DFF_X1 port map( D => n3464, CK => CLK, Q => n10723, QN 
                           => n_2181);
   clk_r_REG1342_S1 : DFF_X1 port map( D => n3463, CK => CLK, Q => n10722, QN 
                           => n_2182);
   clk_r_REG1344_S1 : DFF_X1 port map( D => n3462, CK => CLK, Q => n10721, QN 
                           => n_2183);
   clk_r_REG1346_S1 : DFF_X1 port map( D => n3461, CK => CLK, Q => n10720, QN 
                           => n_2184);
   clk_r_REG1348_S1 : DFF_X1 port map( D => n3460, CK => CLK, Q => n10719, QN 
                           => n_2185);
   clk_r_REG993_S1 : DFF_X1 port map( D => n3418, CK => CLK, Q => n10718, QN =>
                           n_2186);
   clk_r_REG995_S1 : DFF_X1 port map( D => n3419, CK => CLK, Q => n10717, QN =>
                           n_2187);
   clk_r_REG997_S1 : DFF_X1 port map( D => n3420, CK => CLK, Q => n10716, QN =>
                           n_2188);
   clk_r_REG359_S1 : DFF_X1 port map( D => n3476, CK => CLK, Q => n10715, QN =>
                           n_2189);
   clk_r_REG1318_S1 : DFF_X1 port map( D => n3475, CK => CLK, Q => n10714, QN 
                           => n_2190);
   clk_r_REG1320_S1 : DFF_X1 port map( D => n3474, CK => CLK, Q => n10713, QN 
                           => n_2191);
   clk_r_REG1322_S1 : DFF_X1 port map( D => n3473, CK => CLK, Q => n10712, QN 
                           => n_2192);
   clk_r_REG1324_S1 : DFF_X1 port map( D => n3472, CK => CLK, Q => n10711, QN 
                           => n_2193);
   clk_r_REG1326_S1 : DFF_X1 port map( D => n3471, CK => CLK, Q => n10710, QN 
                           => n_2194);
   clk_r_REG971_S1 : DFF_X1 port map( D => n3426, CK => CLK, Q => n10709, QN =>
                           n_2195);
   clk_r_REG973_S1 : DFF_X1 port map( D => n3425, CK => CLK, Q => n10708, QN =>
                           n_2196);
   clk_r_REG975_S1 : DFF_X1 port map( D => n3424, CK => CLK, Q => n10707, QN =>
                           n_2197);
   clk_r_REG977_S1 : DFF_X1 port map( D => n3423, CK => CLK, Q => n10706, QN =>
                           n_2198);
   clk_r_REG979_S1 : DFF_X1 port map( D => n3422, CK => CLK, Q => n10705, QN =>
                           n_2199);
   clk_r_REG981_S1 : DFF_X1 port map( D => n3421, CK => CLK, Q => n10704, QN =>
                           n_2200);
   clk_r_REG983_S1 : DFF_X1 port map( D => n3413, CK => CLK, Q => n10703, QN =>
                           n_2201);
   clk_r_REG985_S1 : DFF_X1 port map( D => n3414, CK => CLK, Q => n10702, QN =>
                           n_2202);
   clk_r_REG987_S1 : DFF_X1 port map( D => n3415, CK => CLK, Q => n10701, QN =>
                           n_2203);
   clk_r_REG989_S1 : DFF_X1 port map( D => n3416, CK => CLK, Q => n10700, QN =>
                           n_2204);
   clk_r_REG991_S1 : DFF_X1 port map( D => n3417, CK => CLK, Q => n10699, QN =>
                           n_2205);
   clk_r_REG949_S1 : DFF_X1 port map( D => n3437, CK => CLK, Q => n10698, QN =>
                           n_2206);
   clk_r_REG951_S1 : DFF_X1 port map( D => n3436, CK => CLK, Q => n10697, QN =>
                           n_2207);
   clk_r_REG953_S1 : DFF_X1 port map( D => n3435, CK => CLK, Q => n10696, QN =>
                           n_2208);
   clk_r_REG955_S1 : DFF_X1 port map( D => n3434, CK => CLK, Q => n10695, QN =>
                           n_2209);
   clk_r_REG957_S1 : DFF_X1 port map( D => n3433, CK => CLK, Q => n10694, QN =>
                           n_2210);
   clk_r_REG959_S1 : DFF_X1 port map( D => n3432, CK => CLK, Q => n10693, QN =>
                           n_2211);
   clk_r_REG961_S1 : DFF_X1 port map( D => n3431, CK => CLK, Q => n10692, QN =>
                           n_2212);
   clk_r_REG963_S1 : DFF_X1 port map( D => n3430, CK => CLK, Q => n10691, QN =>
                           n_2213);
   clk_r_REG965_S1 : DFF_X1 port map( D => n3429, CK => CLK, Q => n10690, QN =>
                           n_2214);
   clk_r_REG967_S1 : DFF_X1 port map( D => n3428, CK => CLK, Q => n10689, QN =>
                           n_2215);
   clk_r_REG969_S1 : DFF_X1 port map( D => n3427, CK => CLK, Q => n10688, QN =>
                           n_2216);
   clk_r_REG3097_S1 : DFF_X1 port map( D => n3512, CK => CLK, Q => n10687, QN 
                           => n_2217);
   clk_r_REG3099_S1 : DFF_X1 port map( D => n3513, CK => CLK, Q => n10686, QN 
                           => n_2218);
   clk_r_REG3101_S1 : DFF_X1 port map( D => n3514, CK => CLK, Q => n10685, QN 
                           => n_2219);
   clk_r_REG3103_S1 : DFF_X1 port map( D => n3515, CK => CLK, Q => n10684, QN 
                           => n_2220);
   clk_r_REG3105_S1 : DFF_X1 port map( D => n3516, CK => CLK, Q => n10683, QN 
                           => n_2221);
   clk_r_REG3075_S1 : DFF_X1 port map( D => n3524, CK => CLK, Q => n10682, QN 
                           => n_2222);
   clk_r_REG3077_S1 : DFF_X1 port map( D => n3523, CK => CLK, Q => n10681, QN 
                           => n_2223);
   clk_r_REG3079_S1 : DFF_X1 port map( D => n3522, CK => CLK, Q => n10680, QN 
                           => n_2224);
   clk_r_REG3081_S1 : DFF_X1 port map( D => n3521, CK => CLK, Q => n10679, QN 
                           => n_2225);
   clk_r_REG3083_S1 : DFF_X1 port map( D => n3520, CK => CLK, Q => n10678, QN 
                           => n_2226);
   clk_r_REG3085_S1 : DFF_X1 port map( D => n3519, CK => CLK, Q => n10677, QN 
                           => n_2227);
   clk_r_REG3087_S1 : DFF_X1 port map( D => n3518, CK => CLK, Q => n10676, QN 
                           => n_2228);
   clk_r_REG3089_S1 : DFF_X1 port map( D => n3517, CK => CLK, Q => n10675, QN 
                           => n_2229);
   clk_r_REG3091_S1 : DFF_X1 port map( D => n3509, CK => CLK, Q => n10674, QN 
                           => n_2230);
   clk_r_REG3093_S1 : DFF_X1 port map( D => n3510, CK => CLK, Q => n10673, QN 
                           => n_2231);
   clk_r_REG3095_S1 : DFF_X1 port map( D => n3511, CK => CLK, Q => n10672, QN 
                           => n_2232);
   clk_r_REG3053_S1 : DFF_X1 port map( D => n3535, CK => CLK, Q => n10671, QN 
                           => n_2233);
   clk_r_REG3055_S1 : DFF_X1 port map( D => n3534, CK => CLK, Q => n10670, QN 
                           => n_2234);
   clk_r_REG3057_S1 : DFF_X1 port map( D => n3533, CK => CLK, Q => n10669, QN 
                           => n_2235);
   clk_r_REG3059_S1 : DFF_X1 port map( D => n3532, CK => CLK, Q => n10668, QN 
                           => n_2236);
   clk_r_REG3061_S1 : DFF_X1 port map( D => n3531, CK => CLK, Q => n10667, QN 
                           => n_2237);
   clk_r_REG3063_S1 : DFF_X1 port map( D => n3530, CK => CLK, Q => n10666, QN 
                           => n_2238);
   clk_r_REG3065_S1 : DFF_X1 port map( D => n3529, CK => CLK, Q => n10665, QN 
                           => n_2239);
   clk_r_REG3067_S1 : DFF_X1 port map( D => n3528, CK => CLK, Q => n10664, QN 
                           => n_2240);
   clk_r_REG3069_S1 : DFF_X1 port map( D => n3527, CK => CLK, Q => n10663, QN 
                           => n_2241);
   clk_r_REG3071_S1 : DFF_X1 port map( D => n3526, CK => CLK, Q => n10662, QN 
                           => n_2242);
   clk_r_REG3073_S1 : DFF_X1 port map( D => n3525, CK => CLK, Q => n10661, QN 
                           => n_2243);
   clk_r_REG2741_S1 : DFF_X1 port map( D => n2925, CK => CLK, Q => n10660, QN 
                           => n_2244);
   clk_r_REG2743_S1 : DFF_X1 port map( D => n2924, CK => CLK, Q => n10659, QN 
                           => n_2245);
   clk_r_REG2745_S1 : DFF_X1 port map( D => n2923, CK => CLK, Q => n10658, QN 
                           => n_2246);
   clk_r_REG2747_S1 : DFF_X1 port map( D => n2922, CK => CLK, Q => n10657, QN 
                           => n_2247);
   clk_r_REG2749_S1 : DFF_X1 port map( D => n2921, CK => CLK, Q => n10656, QN 
                           => n_2248);
   clk_r_REG2751_S1 : DFF_X1 port map( D => n2920, CK => CLK, Q => n10655, QN 
                           => n_2249);
   clk_r_REG2753_S1 : DFF_X1 port map( D => n2919, CK => CLK, Q => n10654, QN 
                           => n_2250);
   clk_r_REG2755_S1 : DFF_X1 port map( D => n2918, CK => CLK, Q => n10653, QN 
                           => n_2251);
   clk_r_REG2757_S1 : DFF_X1 port map( D => n2917, CK => CLK, Q => n10652, QN 
                           => n_2252);
   clk_r_REG2759_S1 : DFF_X1 port map( D => n2916, CK => CLK, Q => n10651, QN 
                           => n_2253);
   clk_r_REG2761_S1 : DFF_X1 port map( D => n2915, CK => CLK, Q => n10650, QN 
                           => n_2254);
   clk_r_REG2862_S1 : DFF_X1 port map( D => n2939, CK => CLK, Q => n10649, QN 
                           => n_2255);
   clk_r_REG2864_S1 : DFF_X1 port map( D => n2940, CK => CLK, Q => n10648, QN 
                           => n_2256);
   clk_r_REG2719_S1 : DFF_X1 port map( D => n2932, CK => CLK, Q => n10647, QN 
                           => n_2257);
   clk_r_REG2729_S1 : DFF_X1 port map( D => n2931, CK => CLK, Q => n10646, QN 
                           => n_2258);
   clk_r_REG2731_S1 : DFF_X1 port map( D => n2930, CK => CLK, Q => n10645, QN 
                           => n_2259);
   clk_r_REG2733_S1 : DFF_X1 port map( D => n2929, CK => CLK, Q => n10644, QN 
                           => n_2260);
   clk_r_REG2735_S1 : DFF_X1 port map( D => n2928, CK => CLK, Q => n10643, QN 
                           => n_2261);
   clk_r_REG2737_S1 : DFF_X1 port map( D => n2927, CK => CLK, Q => n10642, QN 
                           => n_2262);
   clk_r_REG2739_S1 : DFF_X1 port map( D => n2926, CK => CLK, Q => n10641, QN 
                           => n_2263);
   clk_r_REG2840_S1 : DFF_X1 port map( D => n2945, CK => CLK, Q => n10640, QN 
                           => n_2264);
   clk_r_REG2842_S1 : DFF_X1 port map( D => n2944, CK => CLK, Q => n10639, QN 
                           => n_2265);
   clk_r_REG2844_S1 : DFF_X1 port map( D => n2943, CK => CLK, Q => n10638, QN 
                           => n_2266);
   clk_r_REG2846_S1 : DFF_X1 port map( D => n2942, CK => CLK, Q => n10637, QN 
                           => n_2267);
   clk_r_REG2848_S1 : DFF_X1 port map( D => n2941, CK => CLK, Q => n10636, QN 
                           => n_2268);
   clk_r_REG2850_S1 : DFF_X1 port map( D => n2933, CK => CLK, Q => n10635, QN 
                           => n_2269);
   clk_r_REG2852_S1 : DFF_X1 port map( D => n2934, CK => CLK, Q => n10634, QN 
                           => n_2270);
   clk_r_REG2854_S1 : DFF_X1 port map( D => n2935, CK => CLK, Q => n10633, QN 
                           => n_2271);
   clk_r_REG2856_S1 : DFF_X1 port map( D => n2936, CK => CLK, Q => n10632, QN 
                           => n_2272);
   clk_r_REG2858_S1 : DFF_X1 port map( D => n2937, CK => CLK, Q => n10631, QN 
                           => n_2273);
   clk_r_REG2860_S1 : DFF_X1 port map( D => n2938, CK => CLK, Q => n10630, QN 
                           => n_2274);
   clk_r_REG2818_S1 : DFF_X1 port map( D => n2956, CK => CLK, Q => n10629, QN 
                           => n_2275);
   clk_r_REG2820_S1 : DFF_X1 port map( D => n2955, CK => CLK, Q => n10628, QN 
                           => n_2276);
   clk_r_REG2822_S1 : DFF_X1 port map( D => n2954, CK => CLK, Q => n10627, QN 
                           => n_2277);
   clk_r_REG2824_S1 : DFF_X1 port map( D => n2953, CK => CLK, Q => n10626, QN 
                           => n_2278);
   clk_r_REG2826_S1 : DFF_X1 port map( D => n2952, CK => CLK, Q => n10625, QN 
                           => n_2279);
   clk_r_REG2828_S1 : DFF_X1 port map( D => n2951, CK => CLK, Q => n10624, QN 
                           => n_2280);
   clk_r_REG2830_S1 : DFF_X1 port map( D => n2950, CK => CLK, Q => n10623, QN 
                           => n_2281);
   clk_r_REG2832_S1 : DFF_X1 port map( D => n2949, CK => CLK, Q => n10622, QN 
                           => n_2282);
   clk_r_REG2834_S1 : DFF_X1 port map( D => n2948, CK => CLK, Q => n10621, QN 
                           => n_2283);
   clk_r_REG2836_S1 : DFF_X1 port map( D => n2947, CK => CLK, Q => n10620, QN 
                           => n_2284);
   clk_r_REG2838_S1 : DFF_X1 port map( D => n2946, CK => CLK, Q => n10619, QN 
                           => n_2285);
   clk_r_REG2795_S1 : DFF_X1 port map( D => n2964, CK => CLK, Q => n10618, QN 
                           => n_2286);
   clk_r_REG2804_S1 : DFF_X1 port map( D => n2963, CK => CLK, Q => n10617, QN 
                           => n_2287);
   clk_r_REG2806_S1 : DFF_X1 port map( D => n2962, CK => CLK, Q => n10616, QN 
                           => n_2288);
   clk_r_REG2808_S1 : DFF_X1 port map( D => n2961, CK => CLK, Q => n10615, QN 
                           => n_2289);
   clk_r_REG2810_S1 : DFF_X1 port map( D => n2960, CK => CLK, Q => n10614, QN 
                           => n_2290);
   clk_r_REG2812_S1 : DFF_X1 port map( D => n2959, CK => CLK, Q => n10613, QN 
                           => n_2291);
   clk_r_REG2814_S1 : DFF_X1 port map( D => n2958, CK => CLK, Q => n10612, QN 
                           => n_2292);
   clk_r_REG2816_S1 : DFF_X1 port map( D => n2957, CK => CLK, Q => n10611, QN 
                           => n_2293);
   clk_r_REG2914_S1 : DFF_X1 port map( D => n2976, CK => CLK, Q => n10610, QN 
                           => n_2294);
   clk_r_REG2916_S1 : DFF_X1 port map( D => n2975, CK => CLK, Q => n10609, QN 
                           => n_2295);
   clk_r_REG2918_S1 : DFF_X1 port map( D => n2974, CK => CLK, Q => n10608, QN 
                           => n_2296);
   clk_r_REG2920_S1 : DFF_X1 port map( D => n2973, CK => CLK, Q => n10607, QN 
                           => n_2297);
   clk_r_REG2922_S1 : DFF_X1 port map( D => n2965, CK => CLK, Q => n10606, QN 
                           => n_2298);
   clk_r_REG2924_S1 : DFF_X1 port map( D => n2966, CK => CLK, Q => n10605, QN 
                           => n_2299);
   clk_r_REG2926_S1 : DFF_X1 port map( D => n2967, CK => CLK, Q => n10604, QN 
                           => n_2300);
   clk_r_REG2928_S1 : DFF_X1 port map( D => n2968, CK => CLK, Q => n10603, QN 
                           => n_2301);
   clk_r_REG2930_S1 : DFF_X1 port map( D => n2969, CK => CLK, Q => n10602, QN 
                           => n_2302);
   clk_r_REG2932_S1 : DFF_X1 port map( D => n2970, CK => CLK, Q => n10601, QN 
                           => n_2303);
   clk_r_REG2934_S1 : DFF_X1 port map( D => n2971, CK => CLK, Q => n10600, QN 
                           => n_2304);
   clk_r_REG1824_S1 : DFF_X1 port map( D => n2826, CK => CLK, Q => n10599, QN 
                           => n_2305);
   clk_r_REG1826_S1 : DFF_X1 port map( D => n2825, CK => CLK, Q => n10598, QN 
                           => n_2306);
   clk_r_REG1828_S1 : DFF_X1 port map( D => n2824, CK => CLK, Q => n10597, QN 
                           => n_2307);
   clk_r_REG1830_S1 : DFF_X1 port map( D => n2823, CK => CLK, Q => n10596, QN 
                           => n_2308);
   clk_r_REG1832_S1 : DFF_X1 port map( D => n2822, CK => CLK, Q => n10595, QN 
                           => n_2309);
   clk_r_REG1834_S1 : DFF_X1 port map( D => n2821, CK => CLK, Q => n10594, QN 
                           => n_2310);
   clk_r_REG1836_S1 : DFF_X1 port map( D => n2820, CK => CLK, Q => n10593, QN 
                           => n_2311);
   clk_r_REG1838_S1 : DFF_X1 port map( D => n2819, CK => CLK, Q => n10592, QN 
                           => n_2312);
   clk_r_REG1840_S1 : DFF_X1 port map( D => n2818, CK => CLK, Q => n10591, QN 
                           => n_2313);
   clk_r_REG1842_S1 : DFF_X1 port map( D => n2817, CK => CLK, Q => n10590, QN 
                           => n_2314);
   clk_r_REG1844_S1 : DFF_X1 port map( D => n2816, CK => CLK, Q => n10589, QN 
                           => n_2315);
   clk_r_REG1798_S1 : DFF_X1 port map( D => n2836, CK => CLK, Q => n10588, QN 
                           => n_2316);
   clk_r_REG1806_S1 : DFF_X1 port map( D => n2835, CK => CLK, Q => n10587, QN 
                           => n_2317);
   clk_r_REG1808_S1 : DFF_X1 port map( D => n2834, CK => CLK, Q => n10586, QN 
                           => n_2318);
   clk_r_REG1810_S1 : DFF_X1 port map( D => n2833, CK => CLK, Q => n10585, QN 
                           => n_2319);
   clk_r_REG1812_S1 : DFF_X1 port map( D => n2832, CK => CLK, Q => n10584, QN 
                           => n_2320);
   clk_r_REG1814_S1 : DFF_X1 port map( D => n2831, CK => CLK, Q => n10583, QN 
                           => n_2321);
   clk_r_REG1816_S1 : DFF_X1 port map( D => n2830, CK => CLK, Q => n10582, QN 
                           => n_2322);
   clk_r_REG1818_S1 : DFF_X1 port map( D => n2829, CK => CLK, Q => n10581, QN 
                           => n_2323);
   clk_r_REG1820_S1 : DFF_X1 port map( D => n2828, CK => CLK, Q => n10580, QN 
                           => n_2324);
   clk_r_REG1822_S1 : DFF_X1 port map( D => n2827, CK => CLK, Q => n10579, QN 
                           => n_2325);
   clk_r_REG1922_S1 : DFF_X1 port map( D => n2846, CK => CLK, Q => n10578, QN 
                           => n_2326);
   clk_r_REG1924_S1 : DFF_X1 port map( D => n2845, CK => CLK, Q => n10577, QN 
                           => n_2327);
   clk_r_REG1926_S1 : DFF_X1 port map( D => n2837, CK => CLK, Q => n10576, QN 
                           => n_2328);
   clk_r_REG1928_S1 : DFF_X1 port map( D => n2838, CK => CLK, Q => n10575, QN 
                           => n_2329);
   clk_r_REG1930_S1 : DFF_X1 port map( D => n2839, CK => CLK, Q => n10574, QN 
                           => n_2330);
   clk_r_REG1932_S1 : DFF_X1 port map( D => n2840, CK => CLK, Q => n10573, QN 
                           => n_2331);
   clk_r_REG1934_S1 : DFF_X1 port map( D => n2841, CK => CLK, Q => n10572, QN 
                           => n_2332);
   clk_r_REG1936_S1 : DFF_X1 port map( D => n2842, CK => CLK, Q => n10571, QN 
                           => n_2333);
   clk_r_REG1938_S1 : DFF_X1 port map( D => n2843, CK => CLK, Q => n10570, QN 
                           => n_2334);
   clk_r_REG1940_S1 : DFF_X1 port map( D => n2844, CK => CLK, Q => n10569, QN 
                           => n_2335);
   clk_r_REG1900_S1 : DFF_X1 port map( D => n2857, CK => CLK, Q => n10568, QN 
                           => n_2336);
   clk_r_REG1902_S1 : DFF_X1 port map( D => n2856, CK => CLK, Q => n10567, QN 
                           => n_2337);
   clk_r_REG1904_S1 : DFF_X1 port map( D => n2855, CK => CLK, Q => n10566, QN 
                           => n_2338);
   clk_r_REG1906_S1 : DFF_X1 port map( D => n2854, CK => CLK, Q => n10565, QN 
                           => n_2339);
   clk_r_REG1908_S1 : DFF_X1 port map( D => n2853, CK => CLK, Q => n10564, QN 
                           => n_2340);
   clk_r_REG1910_S1 : DFF_X1 port map( D => n2852, CK => CLK, Q => n10563, QN 
                           => n_2341);
   clk_r_REG1912_S1 : DFF_X1 port map( D => n2851, CK => CLK, Q => n10562, QN 
                           => n_2342);
   clk_r_REG1914_S1 : DFF_X1 port map( D => n2850, CK => CLK, Q => n10561, QN 
                           => n_2343);
   clk_r_REG1916_S1 : DFF_X1 port map( D => n2849, CK => CLK, Q => n10560, QN 
                           => n_2344);
   clk_r_REG1918_S1 : DFF_X1 port map( D => n2848, CK => CLK, Q => n10559, QN 
                           => n_2345);
   clk_r_REG1920_S1 : DFF_X1 port map( D => n2847, CK => CLK, Q => n10558, QN 
                           => n_2346);
   clk_r_REG1870_S1 : DFF_X1 port map( D => n2868, CK => CLK, Q => n10557, QN 
                           => n_2347);
   clk_r_REG1880_S1 : DFF_X1 port map( D => n2867, CK => CLK, Q => n10556, QN 
                           => n_2348);
   clk_r_REG1882_S1 : DFF_X1 port map( D => n2866, CK => CLK, Q => n10555, QN 
                           => n_2349);
   clk_r_REG1884_S1 : DFF_X1 port map( D => n2865, CK => CLK, Q => n10554, QN 
                           => n_2350);
   clk_r_REG1886_S1 : DFF_X1 port map( D => n2864, CK => CLK, Q => n10553, QN 
                           => n_2351);
   clk_r_REG1888_S1 : DFF_X1 port map( D => n2863, CK => CLK, Q => n10552, QN 
                           => n_2352);
   clk_r_REG1890_S1 : DFF_X1 port map( D => n2862, CK => CLK, Q => n10551, QN 
                           => n_2353);
   clk_r_REG1892_S1 : DFF_X1 port map( D => n2861, CK => CLK, Q => n10550, QN 
                           => n_2354);
   clk_r_REG1894_S1 : DFF_X1 port map( D => n2860, CK => CLK, Q => n10549, QN 
                           => n_2355);
   clk_r_REG1896_S1 : DFF_X1 port map( D => n2859, CK => CLK, Q => n10548, QN 
                           => n_2356);
   clk_r_REG1898_S1 : DFF_X1 port map( D => n2858, CK => CLK, Q => n10547, QN 
                           => n_2357);
   clk_r_REG1999_S1 : DFF_X1 port map( D => n2877, CK => CLK, Q => n10546, QN 
                           => n_2358);
   clk_r_REG2001_S1 : DFF_X1 port map( D => n2869, CK => CLK, Q => n10545, QN 
                           => n_2359);
   clk_r_REG2003_S1 : DFF_X1 port map( D => n2870, CK => CLK, Q => n10544, QN 
                           => n_2360);
   clk_r_REG2005_S1 : DFF_X1 port map( D => n2871, CK => CLK, Q => n10543, QN 
                           => n_2361);
   clk_r_REG2007_S1 : DFF_X1 port map( D => n2872, CK => CLK, Q => n10542, QN 
                           => n_2362);
   clk_r_REG2009_S1 : DFF_X1 port map( D => n2873, CK => CLK, Q => n10541, QN 
                           => n_2363);
   clk_r_REG2011_S1 : DFF_X1 port map( D => n2874, CK => CLK, Q => n10540, QN 
                           => n_2364);
   clk_r_REG2013_S1 : DFF_X1 port map( D => n2875, CK => CLK, Q => n10539, QN 
                           => n_2365);
   clk_r_REG2015_S1 : DFF_X1 port map( D => n2876, CK => CLK, Q => n10538, QN 
                           => n_2366);
   clk_r_REG2892_S1 : DFF_X1 port map( D => n2987, CK => CLK, Q => n10537, QN 
                           => n_2367);
   clk_r_REG2894_S1 : DFF_X1 port map( D => n2986, CK => CLK, Q => n10536, QN 
                           => n_2368);
   clk_r_REG2896_S1 : DFF_X1 port map( D => n2985, CK => CLK, Q => n10535, QN 
                           => n_2369);
   clk_r_REG2898_S1 : DFF_X1 port map( D => n2984, CK => CLK, Q => n10534, QN 
                           => n_2370);
   clk_r_REG2900_S1 : DFF_X1 port map( D => n2983, CK => CLK, Q => n10533, QN 
                           => n_2371);
   clk_r_REG2902_S1 : DFF_X1 port map( D => n2982, CK => CLK, Q => n10532, QN 
                           => n_2372);
   clk_r_REG2904_S1 : DFF_X1 port map( D => n2981, CK => CLK, Q => n10531, QN 
                           => n_2373);
   clk_r_REG2906_S1 : DFF_X1 port map( D => n2980, CK => CLK, Q => n10530, QN 
                           => n_2374);
   clk_r_REG2908_S1 : DFF_X1 port map( D => n2979, CK => CLK, Q => n10529, QN 
                           => n_2375);
   clk_r_REG2910_S1 : DFF_X1 port map( D => n2978, CK => CLK, Q => n10528, QN 
                           => n_2376);
   clk_r_REG2912_S1 : DFF_X1 port map( D => n2977, CK => CLK, Q => n10527, QN 
                           => n_2377);
   clk_r_REG2868_S1 : DFF_X1 port map( D => n2996, CK => CLK, Q => n10526, QN 
                           => n_2378);
   clk_r_REG2876_S1 : DFF_X1 port map( D => n2995, CK => CLK, Q => n10525, QN 
                           => n_2379);
   clk_r_REG2878_S1 : DFF_X1 port map( D => n2994, CK => CLK, Q => n10524, QN 
                           => n_2380);
   clk_r_REG2880_S1 : DFF_X1 port map( D => n2993, CK => CLK, Q => n10523, QN 
                           => n_2381);
   clk_r_REG2882_S1 : DFF_X1 port map( D => n2992, CK => CLK, Q => n10522, QN 
                           => n_2382);
   clk_r_REG2884_S1 : DFF_X1 port map( D => n2991, CK => CLK, Q => n10521, QN 
                           => n_2383);
   clk_r_REG2886_S1 : DFF_X1 port map( D => n2990, CK => CLK, Q => n10520, QN 
                           => n_2384);
   clk_r_REG2888_S1 : DFF_X1 port map( D => n2989, CK => CLK, Q => n10519, QN 
                           => n_2385);
   clk_r_REG2890_S1 : DFF_X1 port map( D => n2988, CK => CLK, Q => n10518, QN 
                           => n_2386);
   clk_r_REG2993_S1 : DFF_X1 port map( D => n3039, CK => CLK, Q => n10517, QN 
                           => n_2387);
   clk_r_REG2995_S1 : DFF_X1 port map( D => n3038, CK => CLK, Q => n10516, QN 
                           => n_2388);
   clk_r_REG2997_S1 : DFF_X1 port map( D => n3037, CK => CLK, Q => n10515, QN 
                           => n_2389);
   clk_r_REG2999_S1 : DFF_X1 port map( D => n3029, CK => CLK, Q => n10514, QN 
                           => n_2390);
   clk_r_REG3001_S1 : DFF_X1 port map( D => n3030, CK => CLK, Q => n10513, QN 
                           => n_2391);
   clk_r_REG3003_S1 : DFF_X1 port map( D => n3031, CK => CLK, Q => n10512, QN 
                           => n_2392);
   clk_r_REG3005_S1 : DFF_X1 port map( D => n3032, CK => CLK, Q => n10511, QN 
                           => n_2393);
   clk_r_REG3007_S1 : DFF_X1 port map( D => n3033, CK => CLK, Q => n10510, QN 
                           => n_2394);
   clk_r_REG3009_S1 : DFF_X1 port map( D => n3034, CK => CLK, Q => n10509, QN 
                           => n_2395);
   clk_r_REG3011_S1 : DFF_X1 port map( D => n3035, CK => CLK, Q => n10508, QN 
                           => n_2396);
   clk_r_REG3013_S1 : DFF_X1 port map( D => n3036, CK => CLK, Q => n10507, QN 
                           => n_2397);
   clk_r_REG2971_S1 : DFF_X1 port map( D => n3050, CK => CLK, Q => n10506, QN 
                           => n_2398);
   clk_r_REG2973_S1 : DFF_X1 port map( D => n3049, CK => CLK, Q => n10505, QN 
                           => n_2399);
   clk_r_REG2975_S1 : DFF_X1 port map( D => n3048, CK => CLK, Q => n10504, QN 
                           => n_2400);
   clk_r_REG2977_S1 : DFF_X1 port map( D => n3047, CK => CLK, Q => n10503, QN 
                           => n_2401);
   clk_r_REG2979_S1 : DFF_X1 port map( D => n3046, CK => CLK, Q => n10502, QN 
                           => n_2402);
   clk_r_REG2981_S1 : DFF_X1 port map( D => n3045, CK => CLK, Q => n10501, QN 
                           => n_2403);
   clk_r_REG2983_S1 : DFF_X1 port map( D => n3044, CK => CLK, Q => n10500, QN 
                           => n_2404);
   clk_r_REG2985_S1 : DFF_X1 port map( D => n3043, CK => CLK, Q => n10499, QN 
                           => n_2405);
   clk_r_REG2987_S1 : DFF_X1 port map( D => n3042, CK => CLK, Q => n10498, QN 
                           => n_2406);
   clk_r_REG2989_S1 : DFF_X1 port map( D => n3041, CK => CLK, Q => n10497, QN 
                           => n_2407);
   clk_r_REG2991_S1 : DFF_X1 port map( D => n3040, CK => CLK, Q => n10496, QN 
                           => n_2408);
   clk_r_REG2945_S1 : DFF_X1 port map( D => n3060, CK => CLK, Q => n10495, QN 
                           => n_2409);
   clk_r_REG2953_S1 : DFF_X1 port map( D => n3059, CK => CLK, Q => n10494, QN 
                           => n_2410);
   clk_r_REG2955_S1 : DFF_X1 port map( D => n3058, CK => CLK, Q => n10493, QN 
                           => n_2411);
   clk_r_REG2957_S1 : DFF_X1 port map( D => n3057, CK => CLK, Q => n10492, QN 
                           => n_2412);
   clk_r_REG2959_S1 : DFF_X1 port map( D => n3056, CK => CLK, Q => n10491, QN 
                           => n_2413);
   clk_r_REG2961_S1 : DFF_X1 port map( D => n3055, CK => CLK, Q => n10490, QN 
                           => n_2414);
   clk_r_REG2963_S1 : DFF_X1 port map( D => n3054, CK => CLK, Q => n10489, QN 
                           => n_2415);
   clk_r_REG2965_S1 : DFF_X1 port map( D => n3053, CK => CLK, Q => n10488, QN 
                           => n_2416);
   clk_r_REG2967_S1 : DFF_X1 port map( D => n3052, CK => CLK, Q => n10487, QN 
                           => n_2417);
   clk_r_REG2969_S1 : DFF_X1 port map( D => n3051, CK => CLK, Q => n10486, QN 
                           => n_2418);
   clk_r_REG1846_S1 : DFF_X1 port map( D => n2815, CK => CLK, Q => n10485, QN 
                           => n_2419);
   clk_r_REG1848_S1 : DFF_X1 port map( D => n2814, CK => CLK, Q => n10484, QN 
                           => n_2420);
   clk_r_REG1850_S1 : DFF_X1 port map( D => n2813, CK => CLK, Q => n10483, QN 
                           => n_2421);
   clk_r_REG1852_S1 : DFF_X1 port map( D => n2805, CK => CLK, Q => n10482, QN 
                           => n_2422);
   clk_r_REG1854_S1 : DFF_X1 port map( D => n2806, CK => CLK, Q => n10481, QN 
                           => n_2423);
   clk_r_REG1856_S1 : DFF_X1 port map( D => n2807, CK => CLK, Q => n10480, QN 
                           => n_2424);
   clk_r_REG1858_S1 : DFF_X1 port map( D => n2808, CK => CLK, Q => n10479, QN 
                           => n_2425);
   clk_r_REG1860_S1 : DFF_X1 port map( D => n2809, CK => CLK, Q => n10478, QN 
                           => n_2426);
   clk_r_REG1862_S1 : DFF_X1 port map( D => n2810, CK => CLK, Q => n10477, QN 
                           => n_2427);
   clk_r_REG1864_S1 : DFF_X1 port map( D => n2811, CK => CLK, Q => n10476, QN 
                           => n_2428);
   clk_r_REG1866_S1 : DFF_X1 port map( D => n2812, CK => CLK, Q => n10475, QN 
                           => n_2429);
   clk_r_REG2672_S1 : DFF_X1 port map( D => n2792, CK => CLK, Q => n10474, QN 
                           => n_2430);
   clk_r_REG2674_S1 : DFF_X1 port map( D => n2791, CK => CLK, Q => n10473, QN 
                           => n_2431);
   clk_r_REG2676_S1 : DFF_X1 port map( D => n2790, CK => CLK, Q => n10472, QN 
                           => n_2432);
   clk_r_REG2678_S1 : DFF_X1 port map( D => n2789, CK => CLK, Q => n10471, QN 
                           => n_2433);
   clk_r_REG2680_S1 : DFF_X1 port map( D => n2788, CK => CLK, Q => n10470, QN 
                           => n_2434);
   clk_r_REG2694_S1 : DFF_X1 port map( D => n2774, CK => CLK, Q => n10469, QN 
                           => n_2435);
   clk_r_REG2682_S1 : DFF_X1 port map( D => n2787, CK => CLK, Q => n10468, QN 
                           => n_2436);
   clk_r_REG2684_S1 : DFF_X1 port map( D => n2786, CK => CLK, Q => n10467, QN 
                           => n_2437);
   clk_r_REG2686_S1 : DFF_X1 port map( D => n2785, CK => CLK, Q => n10466, QN 
                           => n_2438);
   clk_r_REG2688_S1 : DFF_X1 port map( D => n2784, CK => CLK, Q => n10465, QN 
                           => n_2439);
   clk_r_REG2690_S1 : DFF_X1 port map( D => n2783, CK => CLK, Q => n10464, QN 
                           => n_2440);
   clk_r_REG2652_S1 : DFF_X1 port map( D => n2802, CK => CLK, Q => n10463, QN 
                           => n_2441);
   clk_r_REG2654_S1 : DFF_X1 port map( D => n2801, CK => CLK, Q => n10462, QN 
                           => n_2442);
   clk_r_REG2656_S1 : DFF_X1 port map( D => n2800, CK => CLK, Q => n10461, QN 
                           => n_2443);
   clk_r_REG2658_S1 : DFF_X1 port map( D => n2799, CK => CLK, Q => n10460, QN 
                           => n_2444);
   clk_r_REG2660_S1 : DFF_X1 port map( D => n2798, CK => CLK, Q => n10459, QN 
                           => n_2445);
   clk_r_REG2662_S1 : DFF_X1 port map( D => n2797, CK => CLK, Q => n10458, QN 
                           => n_2446);
   clk_r_REG2664_S1 : DFF_X1 port map( D => n2796, CK => CLK, Q => n10457, QN 
                           => n_2447);
   clk_r_REG2666_S1 : DFF_X1 port map( D => n2795, CK => CLK, Q => n10456, QN 
                           => n_2448);
   clk_r_REG2668_S1 : DFF_X1 port map( D => n2794, CK => CLK, Q => n10455, QN 
                           => n_2449);
   clk_r_REG2670_S1 : DFF_X1 port map( D => n2793, CK => CLK, Q => n10454, QN 
                           => n_2450);
   clk_r_REG2084_S1 : DFF_X1 port map( D => n2998, CK => CLK, Q => n10453, QN 
                           => n_2451);
   clk_r_REG2082_S1 : DFF_X1 port map( D => n2999, CK => CLK, Q => n10452, QN 
                           => n_2452);
   clk_r_REG2080_S1 : DFF_X1 port map( D => n3000, CK => CLK, Q => n10451, QN 
                           => n_2453);
   clk_r_REG2078_S1 : DFF_X1 port map( D => n3001, CK => CLK, Q => n10450, QN 
                           => n_2454);
   clk_r_REG2076_S1 : DFF_X1 port map( D => n3002, CK => CLK, Q => n10449, QN 
                           => n_2455);
   clk_r_REG2074_S1 : DFF_X1 port map( D => n3003, CK => CLK, Q => n10448, QN 
                           => n_2456);
   clk_r_REG2072_S1 : DFF_X1 port map( D => n3004, CK => CLK, Q => n10447, QN 
                           => n_2457);
   clk_r_REG2638_S1 : DFF_X1 port map( D => n2804, CK => CLK, Q => n10446, QN 
                           => n_2458);
   clk_r_REG2650_S1 : DFF_X1 port map( D => n2803, CK => CLK, Q => n10445, QN 
                           => n_2459);
   clk_r_REG2052_S1 : DFF_X1 port map( D => n3014, CK => CLK, Q => n10444, QN 
                           => n_2460);
   clk_r_REG2054_S1 : DFF_X1 port map( D => n3013, CK => CLK, Q => n10443, QN 
                           => n_2461);
   clk_r_REG2056_S1 : DFF_X1 port map( D => n3012, CK => CLK, Q => n10442, QN 
                           => n_2462);
   clk_r_REG2058_S1 : DFF_X1 port map( D => n3011, CK => CLK, Q => n10441, QN 
                           => n_2463);
   clk_r_REG2060_S1 : DFF_X1 port map( D => n3010, CK => CLK, Q => n10440, QN 
                           => n_2464);
   clk_r_REG2062_S1 : DFF_X1 port map( D => n3009, CK => CLK, Q => n10439, QN 
                           => n_2465);
   clk_r_REG2064_S1 : DFF_X1 port map( D => n3008, CK => CLK, Q => n10438, QN 
                           => n_2466);
   clk_r_REG2066_S1 : DFF_X1 port map( D => n3007, CK => CLK, Q => n10437, QN 
                           => n_2467);
   clk_r_REG2068_S1 : DFF_X1 port map( D => n3006, CK => CLK, Q => n10436, QN 
                           => n_2468);
   clk_r_REG2070_S1 : DFF_X1 port map( D => n3005, CK => CLK, Q => n10435, QN 
                           => n_2469);
   clk_r_REG2086_S1 : DFF_X1 port map( D => n2997, CK => CLK, Q => n10434, QN 
                           => n_2470);
   clk_r_REG2030_S1 : DFF_X1 port map( D => n3025, CK => CLK, Q => n10433, QN 
                           => n_2471);
   clk_r_REG2032_S1 : DFF_X1 port map( D => n3024, CK => CLK, Q => n10432, QN 
                           => n_2472);
   clk_r_REG2034_S1 : DFF_X1 port map( D => n3023, CK => CLK, Q => n10431, QN 
                           => n_2473);
   clk_r_REG2036_S1 : DFF_X1 port map( D => n3022, CK => CLK, Q => n10430, QN 
                           => n_2474);
   clk_r_REG2038_S1 : DFF_X1 port map( D => n3021, CK => CLK, Q => n10429, QN 
                           => n_2475);
   clk_r_REG2040_S1 : DFF_X1 port map( D => n3020, CK => CLK, Q => n10428, QN 
                           => n_2476);
   clk_r_REG2042_S1 : DFF_X1 port map( D => n3019, CK => CLK, Q => n10427, QN 
                           => n_2477);
   clk_r_REG2044_S1 : DFF_X1 port map( D => n3018, CK => CLK, Q => n10426, QN 
                           => n_2478);
   clk_r_REG2046_S1 : DFF_X1 port map( D => n3017, CK => CLK, Q => n10425, QN 
                           => n_2479);
   clk_r_REG2048_S1 : DFF_X1 port map( D => n3016, CK => CLK, Q => n10424, QN 
                           => n_2480);
   clk_r_REG2050_S1 : DFF_X1 port map( D => n3015, CK => CLK, Q => n10423, QN 
                           => n_2481);
   clk_r_REG1550_S1 : DFF_X1 port map( D => n3479, CK => CLK, Q => n10422, QN 
                           => n_2482);
   clk_r_REG1548_S1 : DFF_X1 port map( D => n3480, CK => CLK, Q => n10421, QN 
                           => n_2483);
   clk_r_REG1546_S1 : DFF_X1 port map( D => n3481, CK => CLK, Q => n10420, QN 
                           => n_2484);
   clk_r_REG1544_S1 : DFF_X1 port map( D => n3482, CK => CLK, Q => n10419, QN 
                           => n_2485);
   clk_r_REG1542_S1 : DFF_X1 port map( D => n3483, CK => CLK, Q => n10418, QN 
                           => n_2486);
   clk_r_REG1540_S1 : DFF_X1 port map( D => n3484, CK => CLK, Q => n10417, QN 
                           => n_2487);
   clk_r_REG2019_S1 : DFF_X1 port map( D => n3028, CK => CLK, Q => n10416, QN 
                           => n_2488);
   clk_r_REG2026_S1 : DFF_X1 port map( D => n3027, CK => CLK, Q => n10415, QN 
                           => n_2489);
   clk_r_REG2028_S1 : DFF_X1 port map( D => n3026, CK => CLK, Q => n10414, QN 
                           => n_2490);
   clk_r_REG1977_S1 : DFF_X1 port map( D => n2888, CK => CLK, Q => n10413, QN 
                           => n_2491);
   clk_r_REG1979_S1 : DFF_X1 port map( D => n2887, CK => CLK, Q => n10412, QN 
                           => n_2492);
   clk_r_REG1981_S1 : DFF_X1 port map( D => n2886, CK => CLK, Q => n10411, QN 
                           => n_2493);
   clk_r_REG1983_S1 : DFF_X1 port map( D => n2885, CK => CLK, Q => n10410, QN 
                           => n_2494);
   clk_r_REG1985_S1 : DFF_X1 port map( D => n2884, CK => CLK, Q => n10409, QN 
                           => n_2495);
   clk_r_REG1987_S1 : DFF_X1 port map( D => n2883, CK => CLK, Q => n10408, QN 
                           => n_2496);
   clk_r_REG1989_S1 : DFF_X1 port map( D => n2882, CK => CLK, Q => n10407, QN 
                           => n_2497);
   clk_r_REG1991_S1 : DFF_X1 port map( D => n2881, CK => CLK, Q => n10406, QN 
                           => n_2498);
   clk_r_REG1993_S1 : DFF_X1 port map( D => n2880, CK => CLK, Q => n10405, QN 
                           => n_2499);
   clk_r_REG1995_S1 : DFF_X1 port map( D => n2879, CK => CLK, Q => n10404, QN 
                           => n_2500);
   clk_r_REG1997_S1 : DFF_X1 port map( D => n2878, CK => CLK, Q => n10403, QN 
                           => n_2501);
   clk_r_REG1955_S1 : DFF_X1 port map( D => n2899, CK => CLK, Q => n10402, QN 
                           => n_2502);
   clk_r_REG1957_S1 : DFF_X1 port map( D => n2898, CK => CLK, Q => n10401, QN 
                           => n_2503);
   clk_r_REG1959_S1 : DFF_X1 port map( D => n2897, CK => CLK, Q => n10400, QN 
                           => n_2504);
   clk_r_REG1961_S1 : DFF_X1 port map( D => n2896, CK => CLK, Q => n10399, QN 
                           => n_2505);
   clk_r_REG1963_S1 : DFF_X1 port map( D => n2895, CK => CLK, Q => n10398, QN 
                           => n_2506);
   clk_r_REG1965_S1 : DFF_X1 port map( D => n2894, CK => CLK, Q => n10397, QN 
                           => n_2507);
   clk_r_REG1967_S1 : DFF_X1 port map( D => n2893, CK => CLK, Q => n10396, QN 
                           => n_2508);
   clk_r_REG1969_S1 : DFF_X1 port map( D => n2892, CK => CLK, Q => n10395, QN 
                           => n_2509);
   clk_r_REG1971_S1 : DFF_X1 port map( D => n2891, CK => CLK, Q => n10394, QN 
                           => n_2510);
   clk_r_REG1973_S1 : DFF_X1 port map( D => n2890, CK => CLK, Q => n10393, QN 
                           => n_2511);
   clk_r_REG1975_S1 : DFF_X1 port map( D => n2889, CK => CLK, Q => n10392, QN 
                           => n_2512);
   clk_r_REG2614_S1 : DFF_X1 port map( D => n2751, CK => CLK, Q => n10391, QN 
                           => n_2513);
   clk_r_REG2620_S1 : DFF_X1 port map( D => n2743, CK => CLK, Q => n10390, QN 
                           => n_2514);
   clk_r_REG2622_S1 : DFF_X1 port map( D => n2744, CK => CLK, Q => n10389, QN 
                           => n_2515);
   clk_r_REG2624_S1 : DFF_X1 port map( D => n2745, CK => CLK, Q => n10388, QN 
                           => n_2516);
   clk_r_REG2626_S1 : DFF_X1 port map( D => n2746, CK => CLK, Q => n10387, QN 
                           => n_2517);
   clk_r_REG2628_S1 : DFF_X1 port map( D => n2747, CK => CLK, Q => n10386, QN 
                           => n_2518);
   clk_r_REG2630_S1 : DFF_X1 port map( D => n2748, CK => CLK, Q => n10385, QN 
                           => n_2519);
   clk_r_REG2632_S1 : DFF_X1 port map( D => n2749, CK => CLK, Q => n10384, QN 
                           => n_2520);
   clk_r_REG2634_S1 : DFF_X1 port map( D => n2750, CK => CLK, Q => n10383, QN 
                           => n_2521);
   clk_r_REG1947_S1 : DFF_X1 port map( D => n2900, CK => CLK, Q => n10382, QN 
                           => n_2522);
   clk_r_REG2594_S1 : DFF_X1 port map( D => n2761, CK => CLK, Q => n10381, QN 
                           => n_2523);
   clk_r_REG2596_S1 : DFF_X1 port map( D => n2760, CK => CLK, Q => n10380, QN 
                           => n_2524);
   clk_r_REG2598_S1 : DFF_X1 port map( D => n2759, CK => CLK, Q => n10379, QN 
                           => n_2525);
   clk_r_REG2600_S1 : DFF_X1 port map( D => n2758, CK => CLK, Q => n10378, QN 
                           => n_2526);
   clk_r_REG2602_S1 : DFF_X1 port map( D => n2757, CK => CLK, Q => n10377, QN 
                           => n_2527);
   clk_r_REG2604_S1 : DFF_X1 port map( D => n2756, CK => CLK, Q => n10376, QN 
                           => n_2528);
   clk_r_REG2618_S1 : DFF_X1 port map( D => n2742, CK => CLK, Q => n10375, QN 
                           => n_2529);
   clk_r_REG2606_S1 : DFF_X1 port map( D => n2755, CK => CLK, Q => n10374, QN 
                           => n_2530);
   clk_r_REG2608_S1 : DFF_X1 port map( D => n2754, CK => CLK, Q => n10373, QN 
                           => n_2531);
   clk_r_REG2610_S1 : DFF_X1 port map( D => n2753, CK => CLK, Q => n10372, QN 
                           => n_2532);
   clk_r_REG2612_S1 : DFF_X1 port map( D => n2752, CK => CLK, Q => n10371, QN 
                           => n_2533);
   clk_r_REG2574_S1 : DFF_X1 port map( D => n2771, CK => CLK, Q => n10370, QN 
                           => n_2534);
   clk_r_REG2576_S1 : DFF_X1 port map( D => n2770, CK => CLK, Q => n10369, QN 
                           => n_2535);
   clk_r_REG2578_S1 : DFF_X1 port map( D => n2769, CK => CLK, Q => n10368, QN 
                           => n_2536);
   clk_r_REG2580_S1 : DFF_X1 port map( D => n2768, CK => CLK, Q => n10367, QN 
                           => n_2537);
   clk_r_REG2582_S1 : DFF_X1 port map( D => n2767, CK => CLK, Q => n10366, QN 
                           => n_2538);
   clk_r_REG2584_S1 : DFF_X1 port map( D => n2766, CK => CLK, Q => n10365, QN 
                           => n_2539);
   clk_r_REG2586_S1 : DFF_X1 port map( D => n2765, CK => CLK, Q => n10364, QN 
                           => n_2540);
   clk_r_REG2588_S1 : DFF_X1 port map( D => n2764, CK => CLK, Q => n10363, QN 
                           => n_2541);
   clk_r_REG2590_S1 : DFF_X1 port map( D => n2763, CK => CLK, Q => n10362, QN 
                           => n_2542);
   clk_r_REG2592_S1 : DFF_X1 port map( D => n2762, CK => CLK, Q => n10361, QN 
                           => n_2543);
   clk_r_REG2616_S1 : DFF_X1 port map( D => n2741, CK => CLK, Q => n10360, QN 
                           => n_2544);
   clk_r_REG2696_S1 : DFF_X1 port map( D => n2775, CK => CLK, Q => n10359, QN 
                           => n_2545);
   clk_r_REG2698_S1 : DFF_X1 port map( D => n2776, CK => CLK, Q => n10358, QN 
                           => n_2546);
   clk_r_REG2700_S1 : DFF_X1 port map( D => n2777, CK => CLK, Q => n10357, QN 
                           => n_2547);
   clk_r_REG2702_S1 : DFF_X1 port map( D => n2778, CK => CLK, Q => n10356, QN 
                           => n_2548);
   clk_r_REG2704_S1 : DFF_X1 port map( D => n2779, CK => CLK, Q => n10355, QN 
                           => n_2549);
   clk_r_REG2706_S1 : DFF_X1 port map( D => n2780, CK => CLK, Q => n10354, QN 
                           => n_2550);
   clk_r_REG2708_S1 : DFF_X1 port map( D => n2781, CK => CLK, Q => n10353, QN 
                           => n_2551);
   clk_r_REG2710_S1 : DFF_X1 port map( D => n2782, CK => CLK, Q => n10352, QN 
                           => n_2552);
   clk_r_REG2561_S1 : DFF_X1 port map( D => n2772, CK => CLK, Q => n10351, QN 
                           => n_2553);
   clk_r_REG1522_S1 : DFF_X1 port map( D => n3493, CK => CLK, Q => n10350, QN 
                           => n_2554);
   clk_r_REG1524_S1 : DFF_X1 port map( D => n3492, CK => CLK, Q => n10349, QN 
                           => n_2555);
   clk_r_REG1526_S1 : DFF_X1 port map( D => n3491, CK => CLK, Q => n10348, QN 
                           => n_2556);
   clk_r_REG1528_S1 : DFF_X1 port map( D => n3490, CK => CLK, Q => n10347, QN 
                           => n_2557);
   clk_r_REG1530_S1 : DFF_X1 port map( D => n3489, CK => CLK, Q => n10346, QN 
                           => n_2558);
   clk_r_REG1532_S1 : DFF_X1 port map( D => n3488, CK => CLK, Q => n10345, QN 
                           => n_2559);
   clk_r_REG1534_S1 : DFF_X1 port map( D => n3487, CK => CLK, Q => n10344, QN 
                           => n_2560);
   clk_r_REG1536_S1 : DFF_X1 port map( D => n3486, CK => CLK, Q => n10343, QN 
                           => n_2561);
   clk_r_REG1538_S1 : DFF_X1 port map( D => n3485, CK => CLK, Q => n10342, QN 
                           => n_2562);
   clk_r_REG1554_S1 : DFF_X1 port map( D => n3477, CK => CLK, Q => n10341, QN 
                           => n_2563);
   clk_r_REG1552_S1 : DFF_X1 port map( D => n3478, CK => CLK, Q => n10340, QN 
                           => n_2564);
   clk_r_REG1500_S1 : DFF_X1 port map( D => n3504, CK => CLK, Q => n10339, QN 
                           => n_2565);
   clk_r_REG1502_S1 : DFF_X1 port map( D => n3503, CK => CLK, Q => n10338, QN 
                           => n_2566);
   clk_r_REG1504_S1 : DFF_X1 port map( D => n3502, CK => CLK, Q => n10337, QN 
                           => n_2567);
   clk_r_REG1506_S1 : DFF_X1 port map( D => n3501, CK => CLK, Q => n10336, QN 
                           => n_2568);
   clk_r_REG1508_S1 : DFF_X1 port map( D => n3500, CK => CLK, Q => n10335, QN 
                           => n_2569);
   clk_r_REG1510_S1 : DFF_X1 port map( D => n3499, CK => CLK, Q => n10334, QN 
                           => n_2570);
   clk_r_REG1512_S1 : DFF_X1 port map( D => n3498, CK => CLK, Q => n10333, QN 
                           => n_2571);
   clk_r_REG1514_S1 : DFF_X1 port map( D => n3497, CK => CLK, Q => n10332, QN 
                           => n_2572);
   clk_r_REG1516_S1 : DFF_X1 port map( D => n3496, CK => CLK, Q => n10331, QN 
                           => n_2573);
   clk_r_REG1518_S1 : DFF_X1 port map( D => n3495, CK => CLK, Q => n10330, QN 
                           => n_2574);
   clk_r_REG1520_S1 : DFF_X1 port map( D => n3494, CK => CLK, Q => n10329, QN 
                           => n_2575);
   clk_r_REG2544_S1 : DFF_X1 port map( D => n2713, CK => CLK, Q => n10328, QN 
                           => n_2576);
   clk_r_REG2546_S1 : DFF_X1 port map( D => n2714, CK => CLK, Q => n10327, QN 
                           => n_2577);
   clk_r_REG2548_S1 : DFF_X1 port map( D => n2715, CK => CLK, Q => n10326, QN 
                           => n_2578);
   clk_r_REG2550_S1 : DFF_X1 port map( D => n2716, CK => CLK, Q => n10325, QN 
                           => n_2579);
   clk_r_REG2552_S1 : DFF_X1 port map( D => n2717, CK => CLK, Q => n10324, QN 
                           => n_2580);
   clk_r_REG2554_S1 : DFF_X1 port map( D => n2718, CK => CLK, Q => n10323, QN 
                           => n_2581);
   clk_r_REG1487_S1 : DFF_X1 port map( D => n3508, CK => CLK, Q => n10322, QN 
                           => n_2582);
   clk_r_REG1494_S1 : DFF_X1 port map( D => n3507, CK => CLK, Q => n10321, QN 
                           => n_2583);
   clk_r_REG1496_S1 : DFF_X1 port map( D => n3506, CK => CLK, Q => n10320, QN 
                           => n_2584);
   clk_r_REG1498_S1 : DFF_X1 port map( D => n3505, CK => CLK, Q => n10319, QN 
                           => n_2585);
   clk_r_REG2520_S1 : DFF_X1 port map( D => n2726, CK => CLK, Q => n10318, QN 
                           => n_2586);
   clk_r_REG2522_S1 : DFF_X1 port map( D => n2725, CK => CLK, Q => n10317, QN 
                           => n_2587);
   clk_r_REG2524_S1 : DFF_X1 port map( D => n2724, CK => CLK, Q => n10316, QN 
                           => n_2588);
   clk_r_REG2538_S1 : DFF_X1 port map( D => n2710, CK => CLK, Q => n10315, QN 
                           => n_2589);
   clk_r_REG2526_S1 : DFF_X1 port map( D => n2723, CK => CLK, Q => n10314, QN 
                           => n_2590);
   clk_r_REG2528_S1 : DFF_X1 port map( D => n2722, CK => CLK, Q => n10313, QN 
                           => n_2591);
   clk_r_REG2530_S1 : DFF_X1 port map( D => n2721, CK => CLK, Q => n10312, QN 
                           => n_2592);
   clk_r_REG2532_S1 : DFF_X1 port map( D => n2720, CK => CLK, Q => n10311, QN 
                           => n_2593);
   clk_r_REG2534_S1 : DFF_X1 port map( D => n2719, CK => CLK, Q => n10310, QN 
                           => n_2594);
   clk_r_REG2540_S1 : DFF_X1 port map( D => n2711, CK => CLK, Q => n10309, QN 
                           => n_2595);
   clk_r_REG2542_S1 : DFF_X1 port map( D => n2712, CK => CLK, Q => n10308, QN 
                           => n_2596);
   clk_r_REG2500_S1 : DFF_X1 port map( D => n2736, CK => CLK, Q => n10307, QN 
                           => n_2597);
   clk_r_REG2502_S1 : DFF_X1 port map( D => n2735, CK => CLK, Q => n10306, QN 
                           => n_2598);
   clk_r_REG2504_S1 : DFF_X1 port map( D => n2734, CK => CLK, Q => n10305, QN 
                           => n_2599);
   clk_r_REG2506_S1 : DFF_X1 port map( D => n2733, CK => CLK, Q => n10304, QN 
                           => n_2600);
   clk_r_REG2508_S1 : DFF_X1 port map( D => n2732, CK => CLK, Q => n10303, QN 
                           => n_2601);
   clk_r_REG2510_S1 : DFF_X1 port map( D => n2731, CK => CLK, Q => n10302, QN 
                           => n_2602);
   clk_r_REG2512_S1 : DFF_X1 port map( D => n2730, CK => CLK, Q => n10301, QN 
                           => n_2603);
   clk_r_REG2536_S1 : DFF_X1 port map( D => n2709, CK => CLK, Q => n10300, QN 
                           => n_2604);
   clk_r_REG2514_S1 : DFF_X1 port map( D => n2729, CK => CLK, Q => n10299, QN 
                           => n_2605);
   clk_r_REG2516_S1 : DFF_X1 port map( D => n2728, CK => CLK, Q => n10298, QN 
                           => n_2606);
   clk_r_REG2518_S1 : DFF_X1 port map( D => n2727, CK => CLK, Q => n10297, QN 
                           => n_2607);
   clk_r_REG3169_S1 : DFF_X1 port map( D => n3544, CK => CLK, Q => n10296, QN 
                           => n_2608);
   clk_r_REG3171_S1 : DFF_X1 port map( D => n3545, CK => CLK, Q => n10295, QN 
                           => n_2609);
   clk_r_REG3173_S1 : DFF_X1 port map( D => n3546, CK => CLK, Q => n10294, QN 
                           => n_2610);
   clk_r_REG3175_S1 : DFF_X1 port map( D => n3547, CK => CLK, Q => n10293, QN 
                           => n_2611);
   clk_r_REG3177_S1 : DFF_X1 port map( D => n3548, CK => CLK, Q => n10292, QN 
                           => n_2612);
   clk_r_REG2480_S1 : DFF_X1 port map( D => n2740, CK => CLK, Q => n10291, QN 
                           => n_2613);
   clk_r_REG2494_S1 : DFF_X1 port map( D => n2739, CK => CLK, Q => n10290, QN 
                           => n_2614);
   clk_r_REG2496_S1 : DFF_X1 port map( D => n2738, CK => CLK, Q => n10289, QN 
                           => n_2615);
   clk_r_REG2498_S1 : DFF_X1 port map( D => n2737, CK => CLK, Q => n10288, QN 
                           => n_2616);
   clk_r_REG2369_S1 : DFF_X1 port map( D => n2658, CK => CLK, Q => n10287, QN 
                           => n_2617);
   clk_r_REG2371_S1 : DFF_X1 port map( D => n2657, CK => CLK, Q => n10286, QN 
                           => n_2618);
   clk_r_REG2373_S1 : DFF_X1 port map( D => n2656, CK => CLK, Q => n10285, QN 
                           => n_2619);
   clk_r_REG2375_S1 : DFF_X1 port map( D => n2655, CK => CLK, Q => n10284, QN 
                           => n_2620);
   clk_r_REG2381_S1 : DFF_X1 port map( D => n2647, CK => CLK, Q => n10283, QN 
                           => n_2621);
   clk_r_REG2383_S1 : DFF_X1 port map( D => n2648, CK => CLK, Q => n10282, QN 
                           => n_2622);
   clk_r_REG2385_S1 : DFF_X1 port map( D => n2649, CK => CLK, Q => n10281, QN 
                           => n_2623);
   clk_r_REG2387_S1 : DFF_X1 port map( D => n2650, CK => CLK, Q => n10280, QN 
                           => n_2624);
   clk_r_REG2389_S1 : DFF_X1 port map( D => n2651, CK => CLK, Q => n10279, QN 
                           => n_2625);
   clk_r_REG2391_S1 : DFF_X1 port map( D => n2652, CK => CLK, Q => n10278, QN 
                           => n_2626);
   clk_r_REG2393_S1 : DFF_X1 port map( D => n2653, CK => CLK, Q => n10277, QN 
                           => n_2627);
   clk_r_REG2351_S1 : DFF_X1 port map( D => n2667, CK => CLK, Q => n10276, QN 
                           => n_2628);
   clk_r_REG2353_S1 : DFF_X1 port map( D => n2666, CK => CLK, Q => n10275, QN 
                           => n_2629);
   clk_r_REG2377_S1 : DFF_X1 port map( D => n2645, CK => CLK, Q => n10274, QN 
                           => n_2630);
   clk_r_REG2355_S1 : DFF_X1 port map( D => n2665, CK => CLK, Q => n10273, QN 
                           => n_2631);
   clk_r_REG2357_S1 : DFF_X1 port map( D => n2664, CK => CLK, Q => n10272, QN 
                           => n_2632);
   clk_r_REG2359_S1 : DFF_X1 port map( D => n2663, CK => CLK, Q => n10271, QN 
                           => n_2633);
   clk_r_REG2361_S1 : DFF_X1 port map( D => n2662, CK => CLK, Q => n10270, QN 
                           => n_2634);
   clk_r_REG2363_S1 : DFF_X1 port map( D => n2661, CK => CLK, Q => n10269, QN 
                           => n_2635);
   clk_r_REG2365_S1 : DFF_X1 port map( D => n2660, CK => CLK, Q => n10268, QN 
                           => n_2636);
   clk_r_REG2379_S1 : DFF_X1 port map( D => n2646, CK => CLK, Q => n10267, QN 
                           => n_2637);
   clk_r_REG2367_S1 : DFF_X1 port map( D => n2659, CK => CLK, Q => n10266, QN 
                           => n_2638);
   clk_r_REG2323_S1 : DFF_X1 port map( D => n2676, CK => CLK, Q => n10265, QN 
                           => n_2639);
   clk_r_REG2335_S1 : DFF_X1 port map( D => n2675, CK => CLK, Q => n10264, QN 
                           => n_2640);
   clk_r_REG2337_S1 : DFF_X1 port map( D => n2674, CK => CLK, Q => n10263, QN 
                           => n_2641);
   clk_r_REG2339_S1 : DFF_X1 port map( D => n2673, CK => CLK, Q => n10262, QN 
                           => n_2642);
   clk_r_REG2341_S1 : DFF_X1 port map( D => n2672, CK => CLK, Q => n10261, QN 
                           => n_2643);
   clk_r_REG2343_S1 : DFF_X1 port map( D => n2671, CK => CLK, Q => n10260, QN 
                           => n_2644);
   clk_r_REG2345_S1 : DFF_X1 port map( D => n2670, CK => CLK, Q => n10259, QN 
                           => n_2645);
   clk_r_REG2347_S1 : DFF_X1 port map( D => n2669, CK => CLK, Q => n10258, QN 
                           => n_2646);
   clk_r_REG2349_S1 : DFF_X1 port map( D => n2668, CK => CLK, Q => n10257, QN 
                           => n_2647);
   clk_r_REG2452_S1 : DFF_X1 port map( D => n2689, CK => CLK, Q => n10256, QN 
                           => n_2648);
   clk_r_REG2454_S1 : DFF_X1 port map( D => n2688, CK => CLK, Q => n10255, QN 
                           => n_2649);
   clk_r_REG2456_S1 : DFF_X1 port map( D => n2687, CK => CLK, Q => n10254, QN 
                           => n_2650);
   clk_r_REG2462_S1 : DFF_X1 port map( D => n2679, CK => CLK, Q => n10253, QN 
                           => n_2651);
   clk_r_REG2464_S1 : DFF_X1 port map( D => n2680, CK => CLK, Q => n10252, QN 
                           => n_2652);
   clk_r_REG2466_S1 : DFF_X1 port map( D => n2681, CK => CLK, Q => n10251, QN 
                           => n_2653);
   clk_r_REG2468_S1 : DFF_X1 port map( D => n2682, CK => CLK, Q => n10250, QN 
                           => n_2654);
   clk_r_REG2470_S1 : DFF_X1 port map( D => n2683, CK => CLK, Q => n10249, QN 
                           => n_2655);
   clk_r_REG2472_S1 : DFF_X1 port map( D => n2684, CK => CLK, Q => n10248, QN 
                           => n_2656);
   clk_r_REG2474_S1 : DFF_X1 port map( D => n2685, CK => CLK, Q => n10247, QN 
                           => n_2657);
   clk_r_REG2476_S1 : DFF_X1 port map( D => n2686, CK => CLK, Q => n10246, QN 
                           => n_2658);
   clk_r_REG2434_S1 : DFF_X1 port map( D => n2698, CK => CLK, Q => n10245, QN 
                           => n_2659);
   clk_r_REG2458_S1 : DFF_X1 port map( D => n2677, CK => CLK, Q => n10244, QN 
                           => n_2660);
   clk_r_REG2436_S1 : DFF_X1 port map( D => n2697, CK => CLK, Q => n10243, QN 
                           => n_2661);
   clk_r_REG2438_S1 : DFF_X1 port map( D => n2696, CK => CLK, Q => n10242, QN 
                           => n_2662);
   clk_r_REG2440_S1 : DFF_X1 port map( D => n2695, CK => CLK, Q => n10241, QN 
                           => n_2663);
   clk_r_REG2442_S1 : DFF_X1 port map( D => n2694, CK => CLK, Q => n10240, QN 
                           => n_2664);
   clk_r_REG2444_S1 : DFF_X1 port map( D => n2693, CK => CLK, Q => n10239, QN 
                           => n_2665);
   clk_r_REG2446_S1 : DFF_X1 port map( D => n2692, CK => CLK, Q => n10238, QN 
                           => n_2666);
   clk_r_REG2460_S1 : DFF_X1 port map( D => n2678, CK => CLK, Q => n10237, QN 
                           => n_2667);
   clk_r_REG2448_S1 : DFF_X1 port map( D => n2691, CK => CLK, Q => n10236, QN 
                           => n_2668);
   clk_r_REG2450_S1 : DFF_X1 port map( D => n2690, CK => CLK, Q => n10235, QN 
                           => n_2669);
   clk_r_REG2403_S1 : DFF_X1 port map( D => n2708, CK => CLK, Q => n10234, QN 
                           => n_2670);
   clk_r_REG2416_S1 : DFF_X1 port map( D => n2707, CK => CLK, Q => n10233, QN 
                           => n_2671);
   clk_r_REG2418_S1 : DFF_X1 port map( D => n2706, CK => CLK, Q => n10232, QN 
                           => n_2672);
   clk_r_REG2420_S1 : DFF_X1 port map( D => n2705, CK => CLK, Q => n10231, QN 
                           => n_2673);
   clk_r_REG2422_S1 : DFF_X1 port map( D => n2704, CK => CLK, Q => n10230, QN 
                           => n_2674);
   clk_r_REG2424_S1 : DFF_X1 port map( D => n2703, CK => CLK, Q => n10229, QN 
                           => n_2675);
   clk_r_REG2426_S1 : DFF_X1 port map( D => n2702, CK => CLK, Q => n10228, QN 
                           => n_2676);
   clk_r_REG2428_S1 : DFF_X1 port map( D => n2701, CK => CLK, Q => n10227, QN 
                           => n_2677);
   clk_r_REG2430_S1 : DFF_X1 port map( D => n2700, CK => CLK, Q => n10226, QN 
                           => n_2678);
   clk_r_REG2432_S1 : DFF_X1 port map( D => n2699, CK => CLK, Q => n10225, QN 
                           => n_2679);
   clk_r_REG2227_S1 : DFF_X1 port map( D => n2582, CK => CLK, Q => n10224, QN 
                           => n_2680);
   clk_r_REG2215_S1 : DFF_X1 port map( D => n2595, CK => CLK, Q => n10223, QN 
                           => n_2681);
   clk_r_REG2217_S1 : DFF_X1 port map( D => n2594, CK => CLK, Q => n10222, QN 
                           => n_2682);
   clk_r_REG2219_S1 : DFF_X1 port map( D => n2593, CK => CLK, Q => n10221, QN 
                           => n_2683);
   clk_r_REG2221_S1 : DFF_X1 port map( D => n2592, CK => CLK, Q => n10220, QN 
                           => n_2684);
   clk_r_REG2223_S1 : DFF_X1 port map( D => n2591, CK => CLK, Q => n10219, QN 
                           => n_2685);
   clk_r_REG2229_S1 : DFF_X1 port map( D => n2583, CK => CLK, Q => n10218, QN 
                           => n_2686);
   clk_r_REG2231_S1 : DFF_X1 port map( D => n2584, CK => CLK, Q => n10217, QN 
                           => n_2687);
   clk_r_REG2233_S1 : DFF_X1 port map( D => n2585, CK => CLK, Q => n10216, QN 
                           => n_2688);
   clk_r_REG2235_S1 : DFF_X1 port map( D => n2586, CK => CLK, Q => n10215, QN 
                           => n_2689);
   clk_r_REG2237_S1 : DFF_X1 port map( D => n2587, CK => CLK, Q => n10214, QN 
                           => n_2690);
   clk_r_REG2195_S1 : DFF_X1 port map( D => n2605, CK => CLK, Q => n10213, QN 
                           => n_2691);
   clk_r_REG2197_S1 : DFF_X1 port map( D => n2604, CK => CLK, Q => n10212, QN 
                           => n_2692);
   clk_r_REG2199_S1 : DFF_X1 port map( D => n2603, CK => CLK, Q => n10211, QN 
                           => n_2693);
   clk_r_REG2201_S1 : DFF_X1 port map( D => n2602, CK => CLK, Q => n10210, QN 
                           => n_2694);
   clk_r_REG2225_S1 : DFF_X1 port map( D => n2581, CK => CLK, Q => n10209, QN 
                           => n_2695);
   clk_r_REG2203_S1 : DFF_X1 port map( D => n2601, CK => CLK, Q => n10208, QN 
                           => n_2696);
   clk_r_REG2205_S1 : DFF_X1 port map( D => n2600, CK => CLK, Q => n10207, QN 
                           => n_2697);
   clk_r_REG2207_S1 : DFF_X1 port map( D => n2599, CK => CLK, Q => n10206, QN 
                           => n_2698);
   clk_r_REG2209_S1 : DFF_X1 port map( D => n2598, CK => CLK, Q => n10205, QN 
                           => n_2699);
   clk_r_REG2211_S1 : DFF_X1 port map( D => n2597, CK => CLK, Q => n10204, QN 
                           => n_2700);
   clk_r_REG2213_S1 : DFF_X1 port map( D => n2596, CK => CLK, Q => n10203, QN 
                           => n_2701);
   clk_r_REG2317_S1 : DFF_X1 port map( D => n2621, CK => CLK, Q => n10202, QN 
                           => n_2702);
   clk_r_REG2319_S1 : DFF_X1 port map( D => n2622, CK => CLK, Q => n10201, QN 
                           => n_2703);
   clk_r_REG2172_S1 : DFF_X1 port map( D => n2612, CK => CLK, Q => n10200, QN 
                           => n_2704);
   clk_r_REG2183_S1 : DFF_X1 port map( D => n2611, CK => CLK, Q => n10199, QN 
                           => n_2705);
   clk_r_REG2185_S1 : DFF_X1 port map( D => n2610, CK => CLK, Q => n10198, QN 
                           => n_2706);
   clk_r_REG2187_S1 : DFF_X1 port map( D => n2609, CK => CLK, Q => n10197, QN 
                           => n_2707);
   clk_r_REG2189_S1 : DFF_X1 port map( D => n2608, CK => CLK, Q => n10196, QN 
                           => n_2708);
   clk_r_REG2191_S1 : DFF_X1 port map( D => n2607, CK => CLK, Q => n10195, QN 
                           => n_2709);
   clk_r_REG2193_S1 : DFF_X1 port map( D => n2606, CK => CLK, Q => n10194, QN 
                           => n_2710);
   clk_r_REG2291_S1 : DFF_X1 port map( D => n2627, CK => CLK, Q => n10193, QN 
                           => n_2711);
   clk_r_REG2293_S1 : DFF_X1 port map( D => n2626, CK => CLK, Q => n10192, QN 
                           => n_2712);
   clk_r_REG2295_S1 : DFF_X1 port map( D => n2625, CK => CLK, Q => n10191, QN 
                           => n_2713);
   clk_r_REG2297_S1 : DFF_X1 port map( D => n2624, CK => CLK, Q => n10190, QN 
                           => n_2714);
   clk_r_REG2299_S1 : DFF_X1 port map( D => n2623, CK => CLK, Q => n10189, QN 
                           => n_2715);
   clk_r_REG2305_S1 : DFF_X1 port map( D => n2615, CK => CLK, Q => n10188, QN 
                           => n_2716);
   clk_r_REG2307_S1 : DFF_X1 port map( D => n2616, CK => CLK, Q => n10187, QN 
                           => n_2717);
   clk_r_REG2309_S1 : DFF_X1 port map( D => n2617, CK => CLK, Q => n10186, QN 
                           => n_2718);
   clk_r_REG2311_S1 : DFF_X1 port map( D => n2618, CK => CLK, Q => n10185, QN 
                           => n_2719);
   clk_r_REG2313_S1 : DFF_X1 port map( D => n2619, CK => CLK, Q => n10184, QN 
                           => n_2720);
   clk_r_REG2315_S1 : DFF_X1 port map( D => n2620, CK => CLK, Q => n10183, QN 
                           => n_2721);
   clk_r_REG2273_S1 : DFF_X1 port map( D => n2636, CK => CLK, Q => n10182, QN 
                           => n_2722);
   clk_r_REG2275_S1 : DFF_X1 port map( D => n2635, CK => CLK, Q => n10181, QN 
                           => n_2723);
   clk_r_REG2277_S1 : DFF_X1 port map( D => n2634, CK => CLK, Q => n10180, QN 
                           => n_2724);
   clk_r_REG2301_S1 : DFF_X1 port map( D => n2613, CK => CLK, Q => n10179, QN 
                           => n_2725);
   clk_r_REG2279_S1 : DFF_X1 port map( D => n2633, CK => CLK, Q => n10178, QN 
                           => n_2726);
   clk_r_REG2281_S1 : DFF_X1 port map( D => n2632, CK => CLK, Q => n10177, QN 
                           => n_2727);
   clk_r_REG2283_S1 : DFF_X1 port map( D => n2631, CK => CLK, Q => n10176, QN 
                           => n_2728);
   clk_r_REG2285_S1 : DFF_X1 port map( D => n2630, CK => CLK, Q => n10175, QN 
                           => n_2729);
   clk_r_REG2287_S1 : DFF_X1 port map( D => n2629, CK => CLK, Q => n10174, QN 
                           => n_2730);
   clk_r_REG2289_S1 : DFF_X1 port map( D => n2628, CK => CLK, Q => n10173, QN 
                           => n_2731);
   clk_r_REG2303_S1 : DFF_X1 port map( D => n2614, CK => CLK, Q => n10172, QN 
                           => n_2732);
   clk_r_REG2395_S1 : DFF_X1 port map( D => n2654, CK => CLK, Q => n10171, QN 
                           => n_2733);
   clk_r_REG2249_S1 : DFF_X1 port map( D => n2644, CK => CLK, Q => n10170, QN 
                           => n_2734);
   clk_r_REG2259_S1 : DFF_X1 port map( D => n2643, CK => CLK, Q => n10169, QN 
                           => n_2735);
   clk_r_REG2261_S1 : DFF_X1 port map( D => n2642, CK => CLK, Q => n10168, QN 
                           => n_2736);
   clk_r_REG2263_S1 : DFF_X1 port map( D => n2641, CK => CLK, Q => n10167, QN 
                           => n_2737);
   clk_r_REG2265_S1 : DFF_X1 port map( D => n2640, CK => CLK, Q => n10166, QN 
                           => n_2738);
   clk_r_REG2267_S1 : DFF_X1 port map( D => n2639, CK => CLK, Q => n10165, QN 
                           => n_2739);
   clk_r_REG2269_S1 : DFF_X1 port map( D => n2638, CK => CLK, Q => n10164, QN 
                           => n_2740);
   clk_r_REG2271_S1 : DFF_X1 port map( D => n2637, CK => CLK, Q => n10163, QN 
                           => n_2741);
   clk_r_REG3147_S1 : DFF_X1 port map( D => n3556, CK => CLK, Q => n10162, QN 
                           => n_2742);
   clk_r_REG3149_S1 : DFF_X1 port map( D => n3555, CK => CLK, Q => n10161, QN 
                           => n_2743);
   clk_r_REG3151_S1 : DFF_X1 port map( D => n3554, CK => CLK, Q => n10160, QN 
                           => n_2744);
   clk_r_REG3153_S1 : DFF_X1 port map( D => n3553, CK => CLK, Q => n10159, QN 
                           => n_2745);
   clk_r_REG3155_S1 : DFF_X1 port map( D => n3552, CK => CLK, Q => n10158, QN 
                           => n_2746);
   clk_r_REG3157_S1 : DFF_X1 port map( D => n3551, CK => CLK, Q => n10157, QN 
                           => n_2747);
   clk_r_REG3159_S1 : DFF_X1 port map( D => n3550, CK => CLK, Q => n10156, QN 
                           => n_2748);
   clk_r_REG3161_S1 : DFF_X1 port map( D => n3549, CK => CLK, Q => n10155, QN 
                           => n_2749);
   clk_r_REG3163_S1 : DFF_X1 port map( D => n3541, CK => CLK, Q => n10154, QN 
                           => n_2750);
   clk_r_REG3165_S1 : DFF_X1 port map( D => n3542, CK => CLK, Q => n10153, QN 
                           => n_2751);
   clk_r_REG3167_S1 : DFF_X1 port map( D => n3543, CK => CLK, Q => n10152, QN 
                           => n_2752);
   clk_r_REG3125_S1 : DFF_X1 port map( D => n3567, CK => CLK, Q => n10151, QN 
                           => n_2753);
   clk_r_REG3127_S1 : DFF_X1 port map( D => n3566, CK => CLK, Q => n10150, QN 
                           => n_2754);
   clk_r_REG3129_S1 : DFF_X1 port map( D => n3565, CK => CLK, Q => n10149, QN 
                           => n_2755);
   clk_r_REG3131_S1 : DFF_X1 port map( D => n3564, CK => CLK, Q => n10148, QN 
                           => n_2756);
   clk_r_REG3133_S1 : DFF_X1 port map( D => n3563, CK => CLK, Q => n10147, QN 
                           => n_2757);
   clk_r_REG3135_S1 : DFF_X1 port map( D => n3562, CK => CLK, Q => n10146, QN 
                           => n_2758);
   clk_r_REG3137_S1 : DFF_X1 port map( D => n3561, CK => CLK, Q => n10145, QN 
                           => n_2759);
   clk_r_REG3139_S1 : DFF_X1 port map( D => n3560, CK => CLK, Q => n10144, QN 
                           => n_2760);
   clk_r_REG3141_S1 : DFF_X1 port map( D => n3559, CK => CLK, Q => n10143, QN 
                           => n_2761);
   clk_r_REG3143_S1 : DFF_X1 port map( D => n3558, CK => CLK, Q => n10142, QN 
                           => n_2762);
   clk_r_REG3145_S1 : DFF_X1 port map( D => n3557, CK => CLK, Q => n10141, QN 
                           => n_2763);
   clk_r_REG2162_S1 : DFF_X1 port map( D => n2560, CK => CLK, Q => n10140, QN 
                           => n_2764);
   clk_r_REG2164_S1 : DFF_X1 port map( D => n2559, CK => CLK, Q => n10139, QN 
                           => n_2765);
   clk_r_REG2166_S1 : DFF_X1 port map( D => n2558, CK => CLK, Q => n10138, QN 
                           => n_2766);
   clk_r_REG2168_S1 : DFF_X1 port map( D => n2557, CK => CLK, Q => n10137, QN 
                           => n_2767);
   clk_r_REG3114_S1 : DFF_X1 port map( D => n3572, CK => CLK, Q => n10136, QN 
                           => n_2768);
   clk_r_REG3117_S1 : DFF_X1 port map( D => n3571, CK => CLK, Q => n10135, QN 
                           => n_2769);
   clk_r_REG3119_S1 : DFF_X1 port map( D => n3570, CK => CLK, Q => n10134, QN 
                           => n_2770);
   clk_r_REG3121_S1 : DFF_X1 port map( D => n3569, CK => CLK, Q => n10133, QN 
                           => n_2771);
   clk_r_REG3123_S1 : DFF_X1 port map( D => n3568, CK => CLK, Q => n10132, QN 
                           => n_2772);
   clk_r_REG2140_S1 : DFF_X1 port map( D => n2571, CK => CLK, Q => n10131, QN 
                           => n_2773);
   clk_r_REG2142_S1 : DFF_X1 port map( D => n2570, CK => CLK, Q => n10130, QN 
                           => n_2774);
   clk_r_REG2144_S1 : DFF_X1 port map( D => n2569, CK => CLK, Q => n10129, QN 
                           => n_2775);
   clk_r_REG2146_S1 : DFF_X1 port map( D => n2568, CK => CLK, Q => n10128, QN 
                           => n_2776);
   clk_r_REG2148_S1 : DFF_X1 port map( D => n2567, CK => CLK, Q => n10127, QN 
                           => n_2777);
   clk_r_REG2150_S1 : DFF_X1 port map( D => n2566, CK => CLK, Q => n10126, QN 
                           => n_2778);
   clk_r_REG2152_S1 : DFF_X1 port map( D => n2565, CK => CLK, Q => n10125, QN 
                           => n_2779);
   clk_r_REG2154_S1 : DFF_X1 port map( D => n2564, CK => CLK, Q => n10124, QN 
                           => n_2780);
   clk_r_REG2156_S1 : DFF_X1 port map( D => n2563, CK => CLK, Q => n10123, QN 
                           => n_2781);
   clk_r_REG2158_S1 : DFF_X1 port map( D => n2562, CK => CLK, Q => n10122, QN 
                           => n_2782);
   clk_r_REG2160_S1 : DFF_X1 port map( D => n2561, CK => CLK, Q => n10121, QN 
                           => n_2783);
   clk_r_REG2118_S1 : DFF_X1 port map( D => n2555, CK => CLK, Q => n10120, QN 
                           => n_2784);
   clk_r_REG2120_S1 : DFF_X1 port map( D => n2556, CK => CLK, Q => n10119, QN 
                           => n_2785);
   clk_r_REG2122_S1 : DFF_X1 port map( D => n2580, CK => CLK, Q => n10118, QN 
                           => n_2786);
   clk_r_REG2124_S1 : DFF_X1 port map( D => n2579, CK => CLK, Q => n10117, QN 
                           => n_2787);
   clk_r_REG2126_S1 : DFF_X1 port map( D => n2578, CK => CLK, Q => n10116, QN 
                           => n_2788);
   clk_r_REG2128_S1 : DFF_X1 port map( D => n2577, CK => CLK, Q => n10115, QN 
                           => n_2789);
   clk_r_REG2130_S1 : DFF_X1 port map( D => n2576, CK => CLK, Q => n10114, QN 
                           => n_2790);
   clk_r_REG2132_S1 : DFF_X1 port map( D => n2575, CK => CLK, Q => n10113, QN 
                           => n_2791);
   clk_r_REG2134_S1 : DFF_X1 port map( D => n2574, CK => CLK, Q => n10112, QN 
                           => n_2792);
   clk_r_REG2136_S1 : DFF_X1 port map( D => n2573, CK => CLK, Q => n10111, QN 
                           => n_2793);
   clk_r_REG2138_S1 : DFF_X1 port map( D => n2572, CK => CLK, Q => n10110, QN 
                           => n_2794);
   clk_r_REG2239_S1 : DFF_X1 port map( D => n2588, CK => CLK, Q => n10109, QN 
                           => n_2795);
   clk_r_REG2241_S1 : DFF_X1 port map( D => n2589, CK => CLK, Q => n10108, QN 
                           => n_2796);
   clk_r_REG2243_S1 : DFF_X1 port map( D => n2590, CK => CLK, Q => n10107, QN 
                           => n_2797);
   clk_r_REG2108_S1 : DFF_X1 port map( D => n2550, CK => CLK, Q => n10106, QN 
                           => n_2798);
   clk_r_REG2110_S1 : DFF_X1 port map( D => n2551, CK => CLK, Q => n10105, QN 
                           => n_2799);
   clk_r_REG2112_S1 : DFF_X1 port map( D => n2552, CK => CLK, Q => n10104, QN 
                           => n_2800);
   clk_r_REG2114_S1 : DFF_X1 port map( D => n2553, CK => CLK, Q => n10103, QN 
                           => n_2801);
   clk_r_REG3422_S7 : DFFR_X1 port map( D => n4906, CK => CLK, RN => RESET_BAR,
                           Q => n10070, QN => n_2802);
   clk_r_REG3406_S7 : DFFR_X1 port map( D => n4754, CK => CLK, RN => RESET_BAR,
                           Q => n10069, QN => n_2803);
   clk_r_REG3404_S7 : DFFR_X1 port map( D => n4803, CK => CLK, RN => RESET_BAR,
                           Q => n10068, QN => n_2804);
   clk_r_REG3402_S7 : DFFR_X1 port map( D => n4710, CK => CLK, RN => RESET_BAR,
                           Q => n10067, QN => n_2805);
   clk_r_REG3420_S7 : DFFR_X1 port map( D => n4882, CK => CLK, RN => RESET_BAR,
                           Q => n10066, QN => n_2806);
   clk_r_REG3400_S7 : DFFR_X1 port map( D => n4621, CK => CLK, RN => RESET_BAR,
                           Q => n10065, QN => n_2807);
   clk_r_REG3398_S7 : DFFR_X1 port map( D => n4825, CK => CLK, RN => RESET_BAR,
                           Q => n10064, QN => n_2808);
   clk_r_REG3418_S7 : DFFR_X1 port map( D => n4905, CK => CLK, RN => RESET_BAR,
                           Q => n10063, QN => n_2809);
   clk_r_REG3416_S7 : DFFR_X1 port map( D => n4856, CK => CLK, RN => RESET_BAR,
                           Q => n10062, QN => n_2810);
   clk_r_REG3396_S7 : DFFR_X1 port map( D => n4881, CK => CLK, RN => RESET_BAR,
                           Q => n10061, QN => n_2811);
   clk_r_REG3394_S7 : DFFR_X1 port map( D => n4442, CK => CLK, RN => RESET_BAR,
                           Q => n10060, QN => n_2812);
   clk_r_REG3392_S7 : DFFR_X1 port map( D => n4855, CK => CLK, RN => RESET_BAR,
                           Q => n10059, QN => n_2813);
   clk_r_REG3414_S7 : DFFR_X1 port map( D => n4883, CK => CLK, RN => RESET_BAR,
                           Q => n10058, QN => n_2814);
   clk_r_REG3412_S7 : DFFR_X1 port map( D => n4920, CK => CLK, RN => RESET_BAR,
                           Q => n10057, QN => n_2815);
   clk_r_REG3410_S7 : DFFR_X1 port map( D => n4876, CK => CLK, RN => RESET_BAR,
                           Q => n10056, QN => n_2816);
   clk_r_REG3408_S7 : DFFR_X1 port map( D => n4804, CK => CLK, RN => RESET_BAR,
                           Q => n10055, QN => n_2817);
   clk_r_REG3384_S7 : DFFR_X1 port map( D => n5699, CK => CLK, RN => RESET_BAR,
                           Q => n10054, QN => n_2818);
   clk_r_REG3374_S7 : DFFR_X1 port map( D => n5599, CK => CLK, RN => RESET_BAR,
                           Q => n10053, QN => n_2819);
   clk_r_REG3382_S7 : DFFR_X1 port map( D => n5700, CK => CLK, RN => RESET_BAR,
                           Q => n10052, QN => n_2820);
   clk_r_REG3378_S7 : DFFR_X1 port map( D => n5688, CK => CLK, RN => RESET_BAR,
                           Q => n10051, QN => n_2821);
   clk_r_REG3346_S7 : DFFR_X1 port map( D => n5654, CK => CLK, RN => RESET_BAR,
                           Q => n10050, QN => n_2822);
   clk_r_REG3340_S7 : DFFR_X1 port map( D => n5697, CK => CLK, RN => RESET_BAR,
                           Q => n10049, QN => n_2823);
   clk_r_REG3365_S7 : DFFR_X1 port map( D => n5686, CK => CLK, RN => RESET_BAR,
                           Q => n10048, QN => n_2824);
   clk_r_REG3376_S7 : DFFR_X1 port map( D => n5645, CK => CLK, RN => RESET_BAR,
                           Q => n10047, QN => n_2825);
   clk_r_REG3372_S7 : DFFR_X1 port map( D => n5648, CK => CLK, RN => RESET_BAR,
                           Q => n10046, QN => n_2826);
   clk_r_REG3338_S7 : DFFR_X1 port map( D => n5624, CK => CLK, RN => RESET_BAR,
                           Q => n10045, QN => n_2827);
   clk_r_REG3361_S7 : DFFR_X1 port map( D => n5594, CK => CLK, RN => RESET_BAR,
                           Q => n10044, QN => n_2828);
   clk_r_REG3359_S7 : DFFR_X1 port map( D => n5696, CK => CLK, RN => RESET_BAR,
                           Q => n10043, QN => n_2829);
   clk_r_REG3352_S7 : DFFR_X1 port map( D => n5570, CK => CLK, RN => RESET_BAR,
                           Q => n10042, QN => n_2830);
   clk_r_REG3363_S7 : DFFR_X1 port map( D => n5694, CK => CLK, RN => RESET_BAR,
                           Q => n10041, QN => n_2831);
   clk_r_REG3344_S7 : DFFR_X1 port map( D => n5655, CK => CLK, RN => RESET_BAR,
                           Q => n10040, QN => n_2832);
   clk_r_REG3350_S7 : DFFR_X1 port map( D => n5625, CK => CLK, RN => RESET_BAR,
                           Q => n10039, QN => n_2833);
   clk_r_REG2167_S1 : DFF_X1 port map( D => n2557, CK => CLK, Q => n_2834, QN 
                           => n10038);
   clk_r_REG2242_S1 : DFF_X1 port map( D => n2590, CK => CLK, Q => n_2835, QN 
                           => n10037);
   clk_r_REG2318_S1 : DFF_X1 port map( D => n2622, CK => CLK, Q => n_2836, QN 
                           => n10036);
   clk_r_REG2394_S1 : DFF_X1 port map( D => n2654, CK => CLK, Q => n_2837, QN 
                           => n10035);
   clk_r_REG2475_S1 : DFF_X1 port map( D => n2686, CK => CLK, Q => n_2838, QN 
                           => n10034);
   clk_r_REG2553_S1 : DFF_X1 port map( D => n2718, CK => CLK, Q => n_2839, QN 
                           => n10033);
   clk_r_REG2633_S1 : DFF_X1 port map( D => n2750, CK => CLK, Q => n_2840, QN 
                           => n10032);
   clk_r_REG2709_S1 : DFF_X1 port map( D => n2782, CK => CLK, Q => n_2841, QN 
                           => n10031);
   clk_r_REG1865_S1 : DFF_X1 port map( D => n2812, CK => CLK, Q => n_2842, QN 
                           => n10030);
   clk_r_REG1939_S1 : DFF_X1 port map( D => n2844, CK => CLK, Q => n_2843, QN 
                           => n10029);
   clk_r_REG2014_S1 : DFF_X1 port map( D => n2876, CK => CLK, Q => n_2844, QN 
                           => n10028);
   clk_r_REG2788_S1 : DFF_X1 port map( D => n2908, CK => CLK, Q => n_2845, QN 
                           => n10027);
   clk_r_REG2863_S1 : DFF_X1 port map( D => n2940, CK => CLK, Q => n_2846, QN 
                           => n10026);
   clk_r_REG2935_S1 : DFF_X1 port map( D => n2972, CK => CLK, Q => n_2847, QN 
                           => n10025);
   clk_r_REG2071_S1 : DFF_X1 port map( D => n3004, CK => CLK, Q => n_2848, QN 
                           => n10024);
   clk_r_REG3012_S1 : DFF_X1 port map( D => n3036, CK => CLK, Q => n_2849, QN 
                           => n10023);
   clk_r_REG1631_S1 : DFF_X1 port map( D => n3068, CK => CLK, Q => n_2850, QN 
                           => n10022);
   clk_r_REG1708_S1 : DFF_X1 port map( D => n3100, CK => CLK, Q => n_2851, QN 
                           => n10021);
   clk_r_REG1455_S1 : DFF_X1 port map( D => n3132, CK => CLK, Q => n_2852, QN 
                           => n10020);
   clk_r_REG1792_S1 : DFF_X1 port map( D => n3164, CK => CLK, Q => n_2853, QN 
                           => n10019);
   clk_r_REG1071_S1 : DFF_X1 port map( D => n3196, CK => CLK, Q => n_2854, QN 
                           => n10018);
   clk_r_REG1146_S1 : DFF_X1 port map( D => n3228, CK => CLK, Q => n_2855, QN 
                           => n10017);
   clk_r_REG820_S1 : DFF_X1 port map( D => n3260, CK => CLK, Q => n_2856, QN =>
                           n10016);
   clk_r_REG897_S1 : DFF_X1 port map( D => n3292, CK => CLK, Q => n_2857, QN =>
                           n10015);
   clk_r_REG1210_S1 : DFF_X1 port map( D => n3324, CK => CLK, Q => n_2858, QN 
                           => n10014);
   clk_r_REG1276_S1 : DFF_X1 port map( D => n3356, CK => CLK, Q => n_2859, QN 
                           => n10013);
   clk_r_REG723_S1 : DFF_X1 port map( D => n3388, CK => CLK, Q => n_2860, QN =>
                           n10012);
   clk_r_REG996_S1 : DFF_X1 port map( D => n3420, CK => CLK, Q => n_2861, QN =>
                           n10011);
   clk_r_REG1377_S1 : DFF_X1 port map( D => n3452, CK => CLK, Q => n_2862, QN 
                           => n10010);
   clk_r_REG1539_S1 : DFF_X1 port map( D => n3484, CK => CLK, Q => n_2863, QN 
                           => n10009);
   clk_r_REG3104_S1 : DFF_X1 port map( D => n3516, CK => CLK, Q => n_2864, QN 
                           => n10008);
   clk_r_REG3176_S1 : DFF_X1 port map( D => n3548, CK => CLK, Q => n_2865, QN 
                           => n10007);
   clk_r_REG2165_S1 : DFF_X1 port map( D => n2558, CK => CLK, Q => n_2866, QN 
                           => n10006);
   clk_r_REG2240_S1 : DFF_X1 port map( D => n2589, CK => CLK, Q => n_2867, QN 
                           => n10005);
   clk_r_REG2316_S1 : DFF_X1 port map( D => n2621, CK => CLK, Q => n_2868, QN 
                           => n10004);
   clk_r_REG2392_S1 : DFF_X1 port map( D => n2653, CK => CLK, Q => n_2869, QN 
                           => n10003);
   clk_r_REG2473_S1 : DFF_X1 port map( D => n2685, CK => CLK, Q => n_2870, QN 
                           => n10002);
   clk_r_REG2551_S1 : DFF_X1 port map( D => n2717, CK => CLK, Q => n_2871, QN 
                           => n10001);
   clk_r_REG2631_S1 : DFF_X1 port map( D => n2749, CK => CLK, Q => n_2872, QN 
                           => n10000);
   clk_r_REG2707_S1 : DFF_X1 port map( D => n2781, CK => CLK, Q => n_2873, QN 
                           => n9999);
   clk_r_REG1863_S1 : DFF_X1 port map( D => n2811, CK => CLK, Q => n_2874, QN 
                           => n9998);
   clk_r_REG1937_S1 : DFF_X1 port map( D => n2843, CK => CLK, Q => n_2875, QN 
                           => n9997);
   clk_r_REG2012_S1 : DFF_X1 port map( D => n2875, CK => CLK, Q => n_2876, QN 
                           => n9996);
   clk_r_REG2786_S1 : DFF_X1 port map( D => n2907, CK => CLK, Q => n_2877, QN 
                           => n9995);
   clk_r_REG2861_S1 : DFF_X1 port map( D => n2939, CK => CLK, Q => n_2878, QN 
                           => n9994);
   clk_r_REG2933_S1 : DFF_X1 port map( D => n2971, CK => CLK, Q => n_2879, QN 
                           => n9993);
   clk_r_REG2073_S1 : DFF_X1 port map( D => n3003, CK => CLK, Q => n_2880, QN 
                           => n9992);
   clk_r_REG3010_S1 : DFF_X1 port map( D => n3035, CK => CLK, Q => n_2881, QN 
                           => n9991);
   clk_r_REG1629_S1 : DFF_X1 port map( D => n3067, CK => CLK, Q => n_2882, QN 
                           => n9990);
   clk_r_REG1706_S1 : DFF_X1 port map( D => n3099, CK => CLK, Q => n_2883, QN 
                           => n9989);
   clk_r_REG1453_S1 : DFF_X1 port map( D => n3131, CK => CLK, Q => n_2884, QN 
                           => n9988);
   clk_r_REG1790_S1 : DFF_X1 port map( D => n3163, CK => CLK, Q => n_2885, QN 
                           => n9987);
   clk_r_REG1069_S1 : DFF_X1 port map( D => n3195, CK => CLK, Q => n_2886, QN 
                           => n9986);
   clk_r_REG1144_S1 : DFF_X1 port map( D => n3227, CK => CLK, Q => n_2887, QN 
                           => n9985);
   clk_r_REG818_S1 : DFF_X1 port map( D => n3259, CK => CLK, Q => n_2888, QN =>
                           n9984);
   clk_r_REG895_S1 : DFF_X1 port map( D => n3291, CK => CLK, Q => n_2889, QN =>
                           n9983);
   clk_r_REG1208_S1 : DFF_X1 port map( D => n3323, CK => CLK, Q => n_2890, QN 
                           => n9982);
   clk_r_REG1278_S1 : DFF_X1 port map( D => n3355, CK => CLK, Q => n_2891, QN 
                           => n9981);
   clk_r_REG725_S1 : DFF_X1 port map( D => n3387, CK => CLK, Q => n_2892, QN =>
                           n9980);
   clk_r_REG994_S1 : DFF_X1 port map( D => n3419, CK => CLK, Q => n_2893, QN =>
                           n9979);
   clk_r_REG1375_S1 : DFF_X1 port map( D => n3451, CK => CLK, Q => n_2894, QN 
                           => n9978);
   clk_r_REG1541_S1 : DFF_X1 port map( D => n3483, CK => CLK, Q => n_2895, QN 
                           => n9977);
   clk_r_REG3102_S1 : DFF_X1 port map( D => n3515, CK => CLK, Q => n_2896, QN 
                           => n9976);
   clk_r_REG3174_S1 : DFF_X1 port map( D => n3547, CK => CLK, Q => n_2897, QN 
                           => n9975);
   clk_r_REG2163_S1 : DFF_X1 port map( D => n2559, CK => CLK, Q => n_2898, QN 
                           => n9974);
   clk_r_REG2238_S1 : DFF_X1 port map( D => n2588, CK => CLK, Q => n_2899, QN 
                           => n9973);
   clk_r_REG2314_S1 : DFF_X1 port map( D => n2620, CK => CLK, Q => n_2900, QN 
                           => n9972);
   clk_r_REG2390_S1 : DFF_X1 port map( D => n2652, CK => CLK, Q => n_2901, QN 
                           => n9971);
   clk_r_REG2471_S1 : DFF_X1 port map( D => n2684, CK => CLK, Q => n_2902, QN 
                           => n9970);
   clk_r_REG2549_S1 : DFF_X1 port map( D => n2716, CK => CLK, Q => n_2903, QN 
                           => n9969);
   clk_r_REG2629_S1 : DFF_X1 port map( D => n2748, CK => CLK, Q => n_2904, QN 
                           => n9968);
   clk_r_REG2705_S1 : DFF_X1 port map( D => n2780, CK => CLK, Q => n_2905, QN 
                           => n9967);
   clk_r_REG1861_S1 : DFF_X1 port map( D => n2810, CK => CLK, Q => n_2906, QN 
                           => n9966);
   clk_r_REG1935_S1 : DFF_X1 port map( D => n2842, CK => CLK, Q => n_2907, QN 
                           => n9965);
   clk_r_REG2010_S1 : DFF_X1 port map( D => n2874, CK => CLK, Q => n_2908, QN 
                           => n9964);
   clk_r_REG2784_S1 : DFF_X1 port map( D => n2906, CK => CLK, Q => n_2909, QN 
                           => n9963);
   clk_r_REG2859_S1 : DFF_X1 port map( D => n2938, CK => CLK, Q => n_2910, QN 
                           => n9962);
   clk_r_REG2931_S1 : DFF_X1 port map( D => n2970, CK => CLK, Q => n_2911, QN 
                           => n9961);
   clk_r_REG2075_S1 : DFF_X1 port map( D => n3002, CK => CLK, Q => n_2912, QN 
                           => n9960);
   clk_r_REG3008_S1 : DFF_X1 port map( D => n3034, CK => CLK, Q => n_2913, QN 
                           => n9959);
   clk_r_REG1627_S1 : DFF_X1 port map( D => n3066, CK => CLK, Q => n_2914, QN 
                           => n9958);
   clk_r_REG1704_S1 : DFF_X1 port map( D => n3098, CK => CLK, Q => n_2915, QN 
                           => n9957);
   clk_r_REG1451_S1 : DFF_X1 port map( D => n3130, CK => CLK, Q => n_2916, QN 
                           => n9956);
   clk_r_REG1788_S1 : DFF_X1 port map( D => n3162, CK => CLK, Q => n_2917, QN 
                           => n9955);
   clk_r_REG1067_S1 : DFF_X1 port map( D => n3194, CK => CLK, Q => n_2918, QN 
                           => n9954);
   clk_r_REG1142_S1 : DFF_X1 port map( D => n3226, CK => CLK, Q => n_2919, QN 
                           => n9953);
   clk_r_REG816_S1 : DFF_X1 port map( D => n3258, CK => CLK, Q => n_2920, QN =>
                           n9952);
   clk_r_REG893_S1 : DFF_X1 port map( D => n3290, CK => CLK, Q => n_2921, QN =>
                           n9951);
   clk_r_REG1206_S1 : DFF_X1 port map( D => n3322, CK => CLK, Q => n_2922, QN 
                           => n9950);
   clk_r_REG1280_S1 : DFF_X1 port map( D => n3354, CK => CLK, Q => n_2923, QN 
                           => n9949);
   clk_r_REG727_S1 : DFF_X1 port map( D => n3386, CK => CLK, Q => n_2924, QN =>
                           n9948);
   clk_r_REG992_S1 : DFF_X1 port map( D => n3418, CK => CLK, Q => n_2925, QN =>
                           n9947);
   clk_r_REG1373_S1 : DFF_X1 port map( D => n3450, CK => CLK, Q => n_2926, QN 
                           => n9946);
   clk_r_REG1543_S1 : DFF_X1 port map( D => n3482, CK => CLK, Q => n_2927, QN 
                           => n9945);
   clk_r_REG3100_S1 : DFF_X1 port map( D => n3514, CK => CLK, Q => n_2928, QN 
                           => n9944);
   clk_r_REG3172_S1 : DFF_X1 port map( D => n3546, CK => CLK, Q => n_2929, QN 
                           => n9943);
   clk_r_REG2161_S1 : DFF_X1 port map( D => n2560, CK => CLK, Q => n_2930, QN 
                           => n9942);
   clk_r_REG2236_S1 : DFF_X1 port map( D => n2587, CK => CLK, Q => n_2931, QN 
                           => n9941);
   clk_r_REG2312_S1 : DFF_X1 port map( D => n2619, CK => CLK, Q => n_2932, QN 
                           => n9940);
   clk_r_REG2388_S1 : DFF_X1 port map( D => n2651, CK => CLK, Q => n_2933, QN 
                           => n9939);
   clk_r_REG2469_S1 : DFF_X1 port map( D => n2683, CK => CLK, Q => n_2934, QN 
                           => n9938);
   clk_r_REG2547_S1 : DFF_X1 port map( D => n2715, CK => CLK, Q => n_2935, QN 
                           => n9937);
   clk_r_REG2627_S1 : DFF_X1 port map( D => n2747, CK => CLK, Q => n_2936, QN 
                           => n9936);
   clk_r_REG2703_S1 : DFF_X1 port map( D => n2779, CK => CLK, Q => n_2937, QN 
                           => n9935);
   clk_r_REG1859_S1 : DFF_X1 port map( D => n2809, CK => CLK, Q => n_2938, QN 
                           => n9934);
   clk_r_REG1933_S1 : DFF_X1 port map( D => n2841, CK => CLK, Q => n_2939, QN 
                           => n9933);
   clk_r_REG2008_S1 : DFF_X1 port map( D => n2873, CK => CLK, Q => n_2940, QN 
                           => n9932);
   clk_r_REG2782_S1 : DFF_X1 port map( D => n2905, CK => CLK, Q => n_2941, QN 
                           => n9931);
   clk_r_REG2857_S1 : DFF_X1 port map( D => n2937, CK => CLK, Q => n_2942, QN 
                           => n9930);
   clk_r_REG2929_S1 : DFF_X1 port map( D => n2969, CK => CLK, Q => n_2943, QN 
                           => n9929);
   clk_r_REG2077_S1 : DFF_X1 port map( D => n3001, CK => CLK, Q => n_2944, QN 
                           => n9928);
   clk_r_REG3006_S1 : DFF_X1 port map( D => n3033, CK => CLK, Q => n_2945, QN 
                           => n9927);
   clk_r_REG1625_S1 : DFF_X1 port map( D => n3065, CK => CLK, Q => n_2946, QN 
                           => n9926);
   clk_r_REG1702_S1 : DFF_X1 port map( D => n3097, CK => CLK, Q => n_2947, QN 
                           => n9925);
   clk_r_REG1449_S1 : DFF_X1 port map( D => n3129, CK => CLK, Q => n_2948, QN 
                           => n9924);
   clk_r_REG1786_S1 : DFF_X1 port map( D => n3161, CK => CLK, Q => n_2949, QN 
                           => n9923);
   clk_r_REG1065_S1 : DFF_X1 port map( D => n3193, CK => CLK, Q => n_2950, QN 
                           => n9922);
   clk_r_REG1140_S1 : DFF_X1 port map( D => n3225, CK => CLK, Q => n_2951, QN 
                           => n9921);
   clk_r_REG814_S1 : DFF_X1 port map( D => n3257, CK => CLK, Q => n_2952, QN =>
                           n9920);
   clk_r_REG891_S1 : DFF_X1 port map( D => n3289, CK => CLK, Q => n_2953, QN =>
                           n9919);
   clk_r_REG1204_S1 : DFF_X1 port map( D => n3321, CK => CLK, Q => n_2954, QN 
                           => n9918);
   clk_r_REG1282_S1 : DFF_X1 port map( D => n3353, CK => CLK, Q => n_2955, QN 
                           => n9917);
   clk_r_REG729_S1 : DFF_X1 port map( D => n3385, CK => CLK, Q => n_2956, QN =>
                           n9916);
   clk_r_REG990_S1 : DFF_X1 port map( D => n3417, CK => CLK, Q => n_2957, QN =>
                           n9915);
   clk_r_REG1371_S1 : DFF_X1 port map( D => n3449, CK => CLK, Q => n_2958, QN 
                           => n9914);
   clk_r_REG1545_S1 : DFF_X1 port map( D => n3481, CK => CLK, Q => n_2959, QN 
                           => n9913);
   clk_r_REG3098_S1 : DFF_X1 port map( D => n3513, CK => CLK, Q => n_2960, QN 
                           => n9912);
   clk_r_REG3170_S1 : DFF_X1 port map( D => n3545, CK => CLK, Q => n_2961, QN 
                           => n9911);
   clk_r_REG2159_S1 : DFF_X1 port map( D => n2561, CK => CLK, Q => n_2962, QN 
                           => n9910);
   clk_r_REG2234_S1 : DFF_X1 port map( D => n2586, CK => CLK, Q => n_2963, QN 
                           => n9909);
   clk_r_REG2310_S1 : DFF_X1 port map( D => n2618, CK => CLK, Q => n_2964, QN 
                           => n9908);
   clk_r_REG2386_S1 : DFF_X1 port map( D => n2650, CK => CLK, Q => n_2965, QN 
                           => n9907);
   clk_r_REG2467_S1 : DFF_X1 port map( D => n2682, CK => CLK, Q => n_2966, QN 
                           => n9906);
   clk_r_REG2545_S1 : DFF_X1 port map( D => n2714, CK => CLK, Q => n_2967, QN 
                           => n9905);
   clk_r_REG2625_S1 : DFF_X1 port map( D => n2746, CK => CLK, Q => n_2968, QN 
                           => n9904);
   clk_r_REG2701_S1 : DFF_X1 port map( D => n2778, CK => CLK, Q => n_2969, QN 
                           => n9903);
   clk_r_REG1857_S1 : DFF_X1 port map( D => n2808, CK => CLK, Q => n_2970, QN 
                           => n9902);
   clk_r_REG1931_S1 : DFF_X1 port map( D => n2840, CK => CLK, Q => n_2971, QN 
                           => n9901);
   clk_r_REG2006_S1 : DFF_X1 port map( D => n2872, CK => CLK, Q => n_2972, QN 
                           => n9900);
   clk_r_REG2780_S1 : DFF_X1 port map( D => n2904, CK => CLK, Q => n_2973, QN 
                           => n9899);
   clk_r_REG2855_S1 : DFF_X1 port map( D => n2936, CK => CLK, Q => n_2974, QN 
                           => n9898);
   clk_r_REG2927_S1 : DFF_X1 port map( D => n2968, CK => CLK, Q => n_2975, QN 
                           => n9897);
   clk_r_REG2079_S1 : DFF_X1 port map( D => n3000, CK => CLK, Q => n_2976, QN 
                           => n9896);
   clk_r_REG3004_S1 : DFF_X1 port map( D => n3032, CK => CLK, Q => n_2977, QN 
                           => n9895);
   clk_r_REG1623_S1 : DFF_X1 port map( D => n3064, CK => CLK, Q => n_2978, QN 
                           => n9894);
   clk_r_REG1700_S1 : DFF_X1 port map( D => n3096, CK => CLK, Q => n_2979, QN 
                           => n9893);
   clk_r_REG1447_S1 : DFF_X1 port map( D => n3128, CK => CLK, Q => n_2980, QN 
                           => n9892);
   clk_r_REG1784_S1 : DFF_X1 port map( D => n3160, CK => CLK, Q => n_2981, QN 
                           => n9891);
   clk_r_REG1063_S1 : DFF_X1 port map( D => n3192, CK => CLK, Q => n_2982, QN 
                           => n9890);
   clk_r_REG1138_S1 : DFF_X1 port map( D => n3224, CK => CLK, Q => n_2983, QN 
                           => n9889);
   clk_r_REG812_S1 : DFF_X1 port map( D => n3256, CK => CLK, Q => n_2984, QN =>
                           n9888);
   clk_r_REG889_S1 : DFF_X1 port map( D => n3288, CK => CLK, Q => n_2985, QN =>
                           n9887);
   clk_r_REG1202_S1 : DFF_X1 port map( D => n3320, CK => CLK, Q => n_2986, QN 
                           => n9886);
   clk_r_REG1284_S1 : DFF_X1 port map( D => n3352, CK => CLK, Q => n_2987, QN 
                           => n9885);
   clk_r_REG731_S1 : DFF_X1 port map( D => n3384, CK => CLK, Q => n_2988, QN =>
                           n9884);
   clk_r_REG988_S1 : DFF_X1 port map( D => n3416, CK => CLK, Q => n_2989, QN =>
                           n9883);
   clk_r_REG1369_S1 : DFF_X1 port map( D => n3448, CK => CLK, Q => n_2990, QN 
                           => n9882);
   clk_r_REG1547_S1 : DFF_X1 port map( D => n3480, CK => CLK, Q => n_2991, QN 
                           => n9881);
   clk_r_REG3096_S1 : DFF_X1 port map( D => n3512, CK => CLK, Q => n_2992, QN 
                           => n9880);
   clk_r_REG3168_S1 : DFF_X1 port map( D => n3544, CK => CLK, Q => n_2993, QN 
                           => n9879);
   clk_r_REG2157_S1 : DFF_X1 port map( D => n2562, CK => CLK, Q => n_2994, QN 
                           => n9878);
   clk_r_REG2232_S1 : DFF_X1 port map( D => n2585, CK => CLK, Q => n_2995, QN 
                           => n9877);
   clk_r_REG2308_S1 : DFF_X1 port map( D => n2617, CK => CLK, Q => n_2996, QN 
                           => n9876);
   clk_r_REG2384_S1 : DFF_X1 port map( D => n2649, CK => CLK, Q => n_2997, QN 
                           => n9875);
   clk_r_REG2465_S1 : DFF_X1 port map( D => n2681, CK => CLK, Q => n_2998, QN 
                           => n9874);
   clk_r_REG2543_S1 : DFF_X1 port map( D => n2713, CK => CLK, Q => n_2999, QN 
                           => n9873);
   clk_r_REG2623_S1 : DFF_X1 port map( D => n2745, CK => CLK, Q => n_3000, QN 
                           => n9872);
   clk_r_REG2699_S1 : DFF_X1 port map( D => n2777, CK => CLK, Q => n_3001, QN 
                           => n9871);
   clk_r_REG1855_S1 : DFF_X1 port map( D => n2807, CK => CLK, Q => n_3002, QN 
                           => n9870);
   clk_r_REG1929_S1 : DFF_X1 port map( D => n2839, CK => CLK, Q => n_3003, QN 
                           => n9869);
   clk_r_REG2004_S1 : DFF_X1 port map( D => n2871, CK => CLK, Q => n_3004, QN 
                           => n9868);
   clk_r_REG2778_S1 : DFF_X1 port map( D => n2903, CK => CLK, Q => n_3005, QN 
                           => n9867);
   clk_r_REG2853_S1 : DFF_X1 port map( D => n2935, CK => CLK, Q => n_3006, QN 
                           => n9866);
   clk_r_REG2925_S1 : DFF_X1 port map( D => n2967, CK => CLK, Q => n_3007, QN 
                           => n9865);
   clk_r_REG2081_S1 : DFF_X1 port map( D => n2999, CK => CLK, Q => n_3008, QN 
                           => n9864);
   clk_r_REG3002_S1 : DFF_X1 port map( D => n3031, CK => CLK, Q => n_3009, QN 
                           => n9863);
   clk_r_REG1621_S1 : DFF_X1 port map( D => n3063, CK => CLK, Q => n_3010, QN 
                           => n9862);
   clk_r_REG1698_S1 : DFF_X1 port map( D => n3095, CK => CLK, Q => n_3011, QN 
                           => n9861);
   clk_r_REG1445_S1 : DFF_X1 port map( D => n3127, CK => CLK, Q => n_3012, QN 
                           => n9860);
   clk_r_REG1782_S1 : DFF_X1 port map( D => n3159, CK => CLK, Q => n_3013, QN 
                           => n9859);
   clk_r_REG1061_S1 : DFF_X1 port map( D => n3191, CK => CLK, Q => n_3014, QN 
                           => n9858);
   clk_r_REG1136_S1 : DFF_X1 port map( D => n3223, CK => CLK, Q => n_3015, QN 
                           => n9857);
   clk_r_REG810_S1 : DFF_X1 port map( D => n3255, CK => CLK, Q => n_3016, QN =>
                           n9856);
   clk_r_REG887_S1 : DFF_X1 port map( D => n3287, CK => CLK, Q => n_3017, QN =>
                           n9855);
   clk_r_REG1200_S1 : DFF_X1 port map( D => n3319, CK => CLK, Q => n_3018, QN 
                           => n9854);
   clk_r_REG1286_S1 : DFF_X1 port map( D => n3351, CK => CLK, Q => n_3019, QN 
                           => n9853);
   clk_r_REG733_S1 : DFF_X1 port map( D => n3383, CK => CLK, Q => n_3020, QN =>
                           n9852);
   clk_r_REG986_S1 : DFF_X1 port map( D => n3415, CK => CLK, Q => n_3021, QN =>
                           n9851);
   clk_r_REG1367_S1 : DFF_X1 port map( D => n3447, CK => CLK, Q => n_3022, QN 
                           => n9850);
   clk_r_REG1549_S1 : DFF_X1 port map( D => n3479, CK => CLK, Q => n_3023, QN 
                           => n9849);
   clk_r_REG3094_S1 : DFF_X1 port map( D => n3511, CK => CLK, Q => n_3024, QN 
                           => n9848);
   clk_r_REG3166_S1 : DFF_X1 port map( D => n3543, CK => CLK, Q => n_3025, QN 
                           => n9847);
   clk_r_REG2155_S1 : DFF_X1 port map( D => n2563, CK => CLK, Q => n_3026, QN 
                           => n9846);
   clk_r_REG2230_S1 : DFF_X1 port map( D => n2584, CK => CLK, Q => n_3027, QN 
                           => n9845);
   clk_r_REG2306_S1 : DFF_X1 port map( D => n2616, CK => CLK, Q => n_3028, QN 
                           => n9844);
   clk_r_REG2382_S1 : DFF_X1 port map( D => n2648, CK => CLK, Q => n_3029, QN 
                           => n9843);
   clk_r_REG2463_S1 : DFF_X1 port map( D => n2680, CK => CLK, Q => n_3030, QN 
                           => n9842);
   clk_r_REG2541_S1 : DFF_X1 port map( D => n2712, CK => CLK, Q => n_3031, QN 
                           => n9841);
   clk_r_REG2621_S1 : DFF_X1 port map( D => n2744, CK => CLK, Q => n_3032, QN 
                           => n9840);
   clk_r_REG2697_S1 : DFF_X1 port map( D => n2776, CK => CLK, Q => n_3033, QN 
                           => n9839);
   clk_r_REG1853_S1 : DFF_X1 port map( D => n2806, CK => CLK, Q => n_3034, QN 
                           => n9838);
   clk_r_REG1927_S1 : DFF_X1 port map( D => n2838, CK => CLK, Q => n_3035, QN 
                           => n9837);
   clk_r_REG2002_S1 : DFF_X1 port map( D => n2870, CK => CLK, Q => n_3036, QN 
                           => n9836);
   clk_r_REG2776_S1 : DFF_X1 port map( D => n2902, CK => CLK, Q => n_3037, QN 
                           => n9835);
   clk_r_REG2851_S1 : DFF_X1 port map( D => n2934, CK => CLK, Q => n_3038, QN 
                           => n9834);
   clk_r_REG2923_S1 : DFF_X1 port map( D => n2966, CK => CLK, Q => n_3039, QN 
                           => n9833);
   clk_r_REG2083_S1 : DFF_X1 port map( D => n2998, CK => CLK, Q => n_3040, QN 
                           => n9832);
   clk_r_REG3000_S1 : DFF_X1 port map( D => n3030, CK => CLK, Q => n_3041, QN 
                           => n9831);
   clk_r_REG1619_S1 : DFF_X1 port map( D => n3062, CK => CLK, Q => n_3042, QN 
                           => n9830);
   clk_r_REG1696_S1 : DFF_X1 port map( D => n3094, CK => CLK, Q => n_3043, QN 
                           => n9829);
   clk_r_REG1443_S1 : DFF_X1 port map( D => n3126, CK => CLK, Q => n_3044, QN 
                           => n9828);
   clk_r_REG1780_S1 : DFF_X1 port map( D => n3158, CK => CLK, Q => n_3045, QN 
                           => n9827);
   clk_r_REG1059_S1 : DFF_X1 port map( D => n3190, CK => CLK, Q => n_3046, QN 
                           => n9826);
   clk_r_REG1134_S1 : DFF_X1 port map( D => n3222, CK => CLK, Q => n_3047, QN 
                           => n9825);
   clk_r_REG808_S1 : DFF_X1 port map( D => n3254, CK => CLK, Q => n_3048, QN =>
                           n9824);
   clk_r_REG885_S1 : DFF_X1 port map( D => n3286, CK => CLK, Q => n_3049, QN =>
                           n9823);
   clk_r_REG1198_S1 : DFF_X1 port map( D => n3318, CK => CLK, Q => n_3050, QN 
                           => n9822);
   clk_r_REG1288_S1 : DFF_X1 port map( D => n3350, CK => CLK, Q => n_3051, QN 
                           => n9821);
   clk_r_REG735_S1 : DFF_X1 port map( D => n3382, CK => CLK, Q => n_3052, QN =>
                           n9820);
   clk_r_REG984_S1 : DFF_X1 port map( D => n3414, CK => CLK, Q => n_3053, QN =>
                           n9819);
   clk_r_REG1365_S1 : DFF_X1 port map( D => n3446, CK => CLK, Q => n_3054, QN 
                           => n9818);
   clk_r_REG1551_S1 : DFF_X1 port map( D => n3478, CK => CLK, Q => n_3055, QN 
                           => n9817);
   clk_r_REG3092_S1 : DFF_X1 port map( D => n3510, CK => CLK, Q => n_3056, QN 
                           => n9816);
   clk_r_REG3164_S1 : DFF_X1 port map( D => n3542, CK => CLK, Q => n_3057, QN 
                           => n9815);
   clk_r_REG2153_S1 : DFF_X1 port map( D => n2564, CK => CLK, Q => n_3058, QN 
                           => n9814);
   clk_r_REG2228_S1 : DFF_X1 port map( D => n2583, CK => CLK, Q => n_3059, QN 
                           => n9813);
   clk_r_REG2304_S1 : DFF_X1 port map( D => n2615, CK => CLK, Q => n_3060, QN 
                           => n9812);
   clk_r_REG2380_S1 : DFF_X1 port map( D => n2647, CK => CLK, Q => n_3061, QN 
                           => n9811);
   clk_r_REG2461_S1 : DFF_X1 port map( D => n2679, CK => CLK, Q => n_3062, QN 
                           => n9810);
   clk_r_REG2539_S1 : DFF_X1 port map( D => n2711, CK => CLK, Q => n_3063, QN 
                           => n9809);
   clk_r_REG2619_S1 : DFF_X1 port map( D => n2743, CK => CLK, Q => n_3064, QN 
                           => n9808);
   clk_r_REG2695_S1 : DFF_X1 port map( D => n2775, CK => CLK, Q => n_3065, QN 
                           => n9807);
   clk_r_REG1851_S1 : DFF_X1 port map( D => n2805, CK => CLK, Q => n_3066, QN 
                           => n9806);
   clk_r_REG1925_S1 : DFF_X1 port map( D => n2837, CK => CLK, Q => n_3067, QN 
                           => n9805);
   clk_r_REG2000_S1 : DFF_X1 port map( D => n2869, CK => CLK, Q => n_3068, QN 
                           => n9804);
   clk_r_REG2774_S1 : DFF_X1 port map( D => n2901, CK => CLK, Q => n_3069, QN 
                           => n9803);
   clk_r_REG2849_S1 : DFF_X1 port map( D => n2933, CK => CLK, Q => n_3070, QN 
                           => n9802);
   clk_r_REG2921_S1 : DFF_X1 port map( D => n2965, CK => CLK, Q => n_3071, QN 
                           => n9801);
   clk_r_REG2085_S1 : DFF_X1 port map( D => n2997, CK => CLK, Q => n_3072, QN 
                           => n9800);
   clk_r_REG2998_S1 : DFF_X1 port map( D => n3029, CK => CLK, Q => n_3073, QN 
                           => n9799);
   clk_r_REG1617_S1 : DFF_X1 port map( D => n3061, CK => CLK, Q => n_3074, QN 
                           => n9798);
   clk_r_REG1694_S1 : DFF_X1 port map( D => n3093, CK => CLK, Q => n_3075, QN 
                           => n9797);
   clk_r_REG1441_S1 : DFF_X1 port map( D => n3125, CK => CLK, Q => n_3076, QN 
                           => n9796);
   clk_r_REG1778_S1 : DFF_X1 port map( D => n3157, CK => CLK, Q => n_3077, QN 
                           => n9795);
   clk_r_REG1057_S1 : DFF_X1 port map( D => n3189, CK => CLK, Q => n_3078, QN 
                           => n9794);
   clk_r_REG1132_S1 : DFF_X1 port map( D => n3221, CK => CLK, Q => n_3079, QN 
                           => n9793);
   clk_r_REG806_S1 : DFF_X1 port map( D => n3253, CK => CLK, Q => n_3080, QN =>
                           n9792);
   clk_r_REG883_S1 : DFF_X1 port map( D => n3285, CK => CLK, Q => n_3081, QN =>
                           n9791);
   clk_r_REG1196_S1 : DFF_X1 port map( D => n3317, CK => CLK, Q => n_3082, QN 
                           => n9790);
   clk_r_REG1290_S1 : DFF_X1 port map( D => n3349, CK => CLK, Q => n_3083, QN 
                           => n9789);
   clk_r_REG737_S1 : DFF_X1 port map( D => n3381, CK => CLK, Q => n_3084, QN =>
                           n9788);
   clk_r_REG982_S1 : DFF_X1 port map( D => n3413, CK => CLK, Q => n_3085, QN =>
                           n9787);
   clk_r_REG1363_S1 : DFF_X1 port map( D => n3445, CK => CLK, Q => n_3086, QN 
                           => n9786);
   clk_r_REG1553_S1 : DFF_X1 port map( D => n3477, CK => CLK, Q => n_3087, QN 
                           => n9785);
   clk_r_REG3090_S1 : DFF_X1 port map( D => n3509, CK => CLK, Q => n_3088, QN 
                           => n9784);
   clk_r_REG3162_S1 : DFF_X1 port map( D => n3541, CK => CLK, Q => n_3089, QN 
                           => n9783);
   clk_r_REG2151_S1 : DFF_X1 port map( D => n2565, CK => CLK, Q => n_3090, QN 
                           => n9782);
   clk_r_REG2222_S1 : DFF_X1 port map( D => n2591, CK => CLK, Q => n_3091, QN 
                           => n9781);
   clk_r_REG2298_S1 : DFF_X1 port map( D => n2623, CK => CLK, Q => n_3092, QN 
                           => n9780);
   clk_r_REG2374_S1 : DFF_X1 port map( D => n2655, CK => CLK, Q => n_3093, QN 
                           => n9779);
   clk_r_REG2455_S1 : DFF_X1 port map( D => n2687, CK => CLK, Q => n_3094, QN 
                           => n9778);
   clk_r_REG2533_S1 : DFF_X1 port map( D => n2719, CK => CLK, Q => n_3095, QN 
                           => n9777);
   clk_r_REG2613_S1 : DFF_X1 port map( D => n2751, CK => CLK, Q => n_3096, QN 
                           => n9776);
   clk_r_REG2689_S1 : DFF_X1 port map( D => n2783, CK => CLK, Q => n_3097, QN 
                           => n9775);
   clk_r_REG1849_S1 : DFF_X1 port map( D => n2813, CK => CLK, Q => n_3098, QN 
                           => n9774);
   clk_r_REG1923_S1 : DFF_X1 port map( D => n2845, CK => CLK, Q => n_3099, QN 
                           => n9773);
   clk_r_REG1998_S1 : DFF_X1 port map( D => n2877, CK => CLK, Q => n_3100, QN 
                           => n9772);
   clk_r_REG2772_S1 : DFF_X1 port map( D => n2909, CK => CLK, Q => n_3101, QN 
                           => n9771);
   clk_r_REG2847_S1 : DFF_X1 port map( D => n2941, CK => CLK, Q => n_3102, QN 
                           => n9770);
   clk_r_REG2919_S1 : DFF_X1 port map( D => n2973, CK => CLK, Q => n_3103, QN 
                           => n9769);
   clk_r_REG2069_S1 : DFF_X1 port map( D => n3005, CK => CLK, Q => n_3104, QN 
                           => n9768);
   clk_r_REG2996_S1 : DFF_X1 port map( D => n3037, CK => CLK, Q => n_3105, QN 
                           => n9767);
   clk_r_REG1615_S1 : DFF_X1 port map( D => n3069, CK => CLK, Q => n_3106, QN 
                           => n9766);
   clk_r_REG1692_S1 : DFF_X1 port map( D => n3101, CK => CLK, Q => n_3107, QN 
                           => n9765);
   clk_r_REG1439_S1 : DFF_X1 port map( D => n3133, CK => CLK, Q => n_3108, QN 
                           => n9764);
   clk_r_REG1776_S1 : DFF_X1 port map( D => n3165, CK => CLK, Q => n_3109, QN 
                           => n9763);
   clk_r_REG1055_S1 : DFF_X1 port map( D => n3197, CK => CLK, Q => n_3110, QN 
                           => n9762);
   clk_r_REG1130_S1 : DFF_X1 port map( D => n3229, CK => CLK, Q => n_3111, QN 
                           => n9761);
   clk_r_REG804_S1 : DFF_X1 port map( D => n3261, CK => CLK, Q => n_3112, QN =>
                           n9760);
   clk_r_REG881_S1 : DFF_X1 port map( D => n3293, CK => CLK, Q => n_3113, QN =>
                           n9759);
   clk_r_REG1194_S1 : DFF_X1 port map( D => n3325, CK => CLK, Q => n_3114, QN 
                           => n9758);
   clk_r_REG1274_S1 : DFF_X1 port map( D => n3357, CK => CLK, Q => n_3115, QN 
                           => n9757);
   clk_r_REG721_S1 : DFF_X1 port map( D => n3389, CK => CLK, Q => n_3116, QN =>
                           n9756);
   clk_r_REG980_S1 : DFF_X1 port map( D => n3421, CK => CLK, Q => n_3117, QN =>
                           n9755);
   clk_r_REG1361_S1 : DFF_X1 port map( D => n3453, CK => CLK, Q => n_3118, QN 
                           => n9754);
   clk_r_REG1537_S1 : DFF_X1 port map( D => n3485, CK => CLK, Q => n_3119, QN 
                           => n9753);
   clk_r_REG3088_S1 : DFF_X1 port map( D => n3517, CK => CLK, Q => n_3120, QN 
                           => n9752);
   clk_r_REG3160_S1 : DFF_X1 port map( D => n3549, CK => CLK, Q => n_3121, QN 
                           => n9751);
   clk_r_REG2149_S1 : DFF_X1 port map( D => n2566, CK => CLK, Q => n_3122, QN 
                           => n9750);
   clk_r_REG2220_S1 : DFF_X1 port map( D => n2592, CK => CLK, Q => n_3123, QN 
                           => n9749);
   clk_r_REG2296_S1 : DFF_X1 port map( D => n2624, CK => CLK, Q => n_3124, QN 
                           => n9748);
   clk_r_REG2372_S1 : DFF_X1 port map( D => n2656, CK => CLK, Q => n_3125, QN 
                           => n9747);
   clk_r_REG2453_S1 : DFF_X1 port map( D => n2688, CK => CLK, Q => n_3126, QN 
                           => n9746);
   clk_r_REG2531_S1 : DFF_X1 port map( D => n2720, CK => CLK, Q => n_3127, QN 
                           => n9745);
   clk_r_REG2611_S1 : DFF_X1 port map( D => n2752, CK => CLK, Q => n_3128, QN 
                           => n9744);
   clk_r_REG2687_S1 : DFF_X1 port map( D => n2784, CK => CLK, Q => n_3129, QN 
                           => n9743);
   clk_r_REG1847_S1 : DFF_X1 port map( D => n2814, CK => CLK, Q => n_3130, QN 
                           => n9742);
   clk_r_REG1921_S1 : DFF_X1 port map( D => n2846, CK => CLK, Q => n_3131, QN 
                           => n9741);
   clk_r_REG1996_S1 : DFF_X1 port map( D => n2878, CK => CLK, Q => n_3132, QN 
                           => n9740);
   clk_r_REG2770_S1 : DFF_X1 port map( D => n2910, CK => CLK, Q => n_3133, QN 
                           => n9739);
   clk_r_REG2845_S1 : DFF_X1 port map( D => n2942, CK => CLK, Q => n_3134, QN 
                           => n9738);
   clk_r_REG2917_S1 : DFF_X1 port map( D => n2974, CK => CLK, Q => n_3135, QN 
                           => n9737);
   clk_r_REG2067_S1 : DFF_X1 port map( D => n3006, CK => CLK, Q => n_3136, QN 
                           => n9736);
   clk_r_REG2994_S1 : DFF_X1 port map( D => n3038, CK => CLK, Q => n_3137, QN 
                           => n9735);
   clk_r_REG1613_S1 : DFF_X1 port map( D => n3070, CK => CLK, Q => n_3138, QN 
                           => n9734);
   clk_r_REG1690_S1 : DFF_X1 port map( D => n3102, CK => CLK, Q => n_3139, QN 
                           => n9733);
   clk_r_REG1437_S1 : DFF_X1 port map( D => n3134, CK => CLK, Q => n_3140, QN 
                           => n9732);
   clk_r_REG1774_S1 : DFF_X1 port map( D => n3166, CK => CLK, Q => n_3141, QN 
                           => n9731);
   clk_r_REG1053_S1 : DFF_X1 port map( D => n3198, CK => CLK, Q => n_3142, QN 
                           => n9730);
   clk_r_REG1128_S1 : DFF_X1 port map( D => n3230, CK => CLK, Q => n_3143, QN 
                           => n9729);
   clk_r_REG802_S1 : DFF_X1 port map( D => n3262, CK => CLK, Q => n_3144, QN =>
                           n9728);
   clk_r_REG879_S1 : DFF_X1 port map( D => n3294, CK => CLK, Q => n_3145, QN =>
                           n9727);
   clk_r_REG1192_S1 : DFF_X1 port map( D => n3326, CK => CLK, Q => n_3146, QN 
                           => n9726);
   clk_r_REG1272_S1 : DFF_X1 port map( D => n3358, CK => CLK, Q => n_3147, QN 
                           => n9725);
   clk_r_REG719_S1 : DFF_X1 port map( D => n3390, CK => CLK, Q => n_3148, QN =>
                           n9724);
   clk_r_REG978_S1 : DFF_X1 port map( D => n3422, CK => CLK, Q => n_3149, QN =>
                           n9723);
   clk_r_REG1359_S1 : DFF_X1 port map( D => n3454, CK => CLK, Q => n_3150, QN 
                           => n9722);
   clk_r_REG1535_S1 : DFF_X1 port map( D => n3486, CK => CLK, Q => n_3151, QN 
                           => n9721);
   clk_r_REG3086_S1 : DFF_X1 port map( D => n3518, CK => CLK, Q => n_3152, QN 
                           => n9720);
   clk_r_REG3158_S1 : DFF_X1 port map( D => n3550, CK => CLK, Q => n_3153, QN 
                           => n9719);
   clk_r_REG2147_S1 : DFF_X1 port map( D => n2567, CK => CLK, Q => n_3154, QN 
                           => n9718);
   clk_r_REG2218_S1 : DFF_X1 port map( D => n2593, CK => CLK, Q => n_3155, QN 
                           => n9717);
   clk_r_REG2294_S1 : DFF_X1 port map( D => n2625, CK => CLK, Q => n_3156, QN 
                           => n9716);
   clk_r_REG2370_S1 : DFF_X1 port map( D => n2657, CK => CLK, Q => n_3157, QN 
                           => n9715);
   clk_r_REG2451_S1 : DFF_X1 port map( D => n2689, CK => CLK, Q => n_3158, QN 
                           => n9714);
   clk_r_REG2529_S1 : DFF_X1 port map( D => n2721, CK => CLK, Q => n_3159, QN 
                           => n9713);
   clk_r_REG2609_S1 : DFF_X1 port map( D => n2753, CK => CLK, Q => n_3160, QN 
                           => n9712);
   clk_r_REG2685_S1 : DFF_X1 port map( D => n2785, CK => CLK, Q => n_3161, QN 
                           => n9711);
   clk_r_REG1845_S1 : DFF_X1 port map( D => n2815, CK => CLK, Q => n_3162, QN 
                           => n9710);
   clk_r_REG1919_S1 : DFF_X1 port map( D => n2847, CK => CLK, Q => n_3163, QN 
                           => n9709);
   clk_r_REG1994_S1 : DFF_X1 port map( D => n2879, CK => CLK, Q => n_3164, QN 
                           => n9708);
   clk_r_REG2768_S1 : DFF_X1 port map( D => n2911, CK => CLK, Q => n_3165, QN 
                           => n9707);
   clk_r_REG2843_S1 : DFF_X1 port map( D => n2943, CK => CLK, Q => n_3166, QN 
                           => n9706);
   clk_r_REG2915_S1 : DFF_X1 port map( D => n2975, CK => CLK, Q => n_3167, QN 
                           => n9705);
   clk_r_REG2065_S1 : DFF_X1 port map( D => n3007, CK => CLK, Q => n_3168, QN 
                           => n9704);
   clk_r_REG2992_S1 : DFF_X1 port map( D => n3039, CK => CLK, Q => n_3169, QN 
                           => n9703);
   clk_r_REG1611_S1 : DFF_X1 port map( D => n3071, CK => CLK, Q => n_3170, QN 
                           => n9702);
   clk_r_REG1688_S1 : DFF_X1 port map( D => n3103, CK => CLK, Q => n_3171, QN 
                           => n9701);
   clk_r_REG1435_S1 : DFF_X1 port map( D => n3135, CK => CLK, Q => n_3172, QN 
                           => n9700);
   clk_r_REG1772_S1 : DFF_X1 port map( D => n3167, CK => CLK, Q => n_3173, QN 
                           => n9699);
   clk_r_REG1051_S1 : DFF_X1 port map( D => n3199, CK => CLK, Q => n_3174, QN 
                           => n9698);
   clk_r_REG1126_S1 : DFF_X1 port map( D => n3231, CK => CLK, Q => n_3175, QN 
                           => n9697);
   clk_r_REG800_S1 : DFF_X1 port map( D => n3263, CK => CLK, Q => n_3176, QN =>
                           n9696);
   clk_r_REG877_S1 : DFF_X1 port map( D => n3295, CK => CLK, Q => n_3177, QN =>
                           n9695);
   clk_r_REG1190_S1 : DFF_X1 port map( D => n3327, CK => CLK, Q => n_3178, QN 
                           => n9694);
   clk_r_REG1270_S1 : DFF_X1 port map( D => n3359, CK => CLK, Q => n_3179, QN 
                           => n9693);
   clk_r_REG717_S1 : DFF_X1 port map( D => n3391, CK => CLK, Q => n_3180, QN =>
                           n9692);
   clk_r_REG976_S1 : DFF_X1 port map( D => n3423, CK => CLK, Q => n_3181, QN =>
                           n9691);
   clk_r_REG1357_S1 : DFF_X1 port map( D => n3455, CK => CLK, Q => n_3182, QN 
                           => n9690);
   clk_r_REG1533_S1 : DFF_X1 port map( D => n3487, CK => CLK, Q => n_3183, QN 
                           => n9689);
   clk_r_REG3084_S1 : DFF_X1 port map( D => n3519, CK => CLK, Q => n_3184, QN 
                           => n9688);
   clk_r_REG3156_S1 : DFF_X1 port map( D => n3551, CK => CLK, Q => n_3185, QN 
                           => n9687);
   clk_r_REG2145_S1 : DFF_X1 port map( D => n2568, CK => CLK, Q => n_3186, QN 
                           => n9686);
   clk_r_REG2216_S1 : DFF_X1 port map( D => n2594, CK => CLK, Q => n_3187, QN 
                           => n9685);
   clk_r_REG2292_S1 : DFF_X1 port map( D => n2626, CK => CLK, Q => n_3188, QN 
                           => n9684);
   clk_r_REG2368_S1 : DFF_X1 port map( D => n2658, CK => CLK, Q => n_3189, QN 
                           => n9683);
   clk_r_REG2449_S1 : DFF_X1 port map( D => n2690, CK => CLK, Q => n_3190, QN 
                           => n9682);
   clk_r_REG2527_S1 : DFF_X1 port map( D => n2722, CK => CLK, Q => n_3191, QN 
                           => n9681);
   clk_r_REG2607_S1 : DFF_X1 port map( D => n2754, CK => CLK, Q => n_3192, QN 
                           => n9680);
   clk_r_REG2683_S1 : DFF_X1 port map( D => n2786, CK => CLK, Q => n_3193, QN 
                           => n9679);
   clk_r_REG1843_S1 : DFF_X1 port map( D => n2816, CK => CLK, Q => n_3194, QN 
                           => n9678);
   clk_r_REG1917_S1 : DFF_X1 port map( D => n2848, CK => CLK, Q => n_3195, QN 
                           => n9677);
   clk_r_REG1992_S1 : DFF_X1 port map( D => n2880, CK => CLK, Q => n_3196, QN 
                           => n9676);
   clk_r_REG2766_S1 : DFF_X1 port map( D => n2912, CK => CLK, Q => n_3197, QN 
                           => n9675);
   clk_r_REG2841_S1 : DFF_X1 port map( D => n2944, CK => CLK, Q => n_3198, QN 
                           => n9674);
   clk_r_REG2913_S1 : DFF_X1 port map( D => n2976, CK => CLK, Q => n_3199, QN 
                           => n9673);
   clk_r_REG2063_S1 : DFF_X1 port map( D => n3008, CK => CLK, Q => n_3200, QN 
                           => n9672);
   clk_r_REG2990_S1 : DFF_X1 port map( D => n3040, CK => CLK, Q => n_3201, QN 
                           => n9671);
   clk_r_REG1609_S1 : DFF_X1 port map( D => n3072, CK => CLK, Q => n_3202, QN 
                           => n9670);
   clk_r_REG1686_S1 : DFF_X1 port map( D => n3104, CK => CLK, Q => n_3203, QN 
                           => n9669);
   clk_r_REG1433_S1 : DFF_X1 port map( D => n3136, CK => CLK, Q => n_3204, QN 
                           => n9668);
   clk_r_REG1770_S1 : DFF_X1 port map( D => n3168, CK => CLK, Q => n_3205, QN 
                           => n9667);
   clk_r_REG1049_S1 : DFF_X1 port map( D => n3200, CK => CLK, Q => n_3206, QN 
                           => n9666);
   clk_r_REG1124_S1 : DFF_X1 port map( D => n3232, CK => CLK, Q => n_3207, QN 
                           => n9665);
   clk_r_REG798_S1 : DFF_X1 port map( D => n3264, CK => CLK, Q => n_3208, QN =>
                           n9664);
   clk_r_REG875_S1 : DFF_X1 port map( D => n3296, CK => CLK, Q => n_3209, QN =>
                           n9663);
   clk_r_REG1188_S1 : DFF_X1 port map( D => n3328, CK => CLK, Q => n_3210, QN 
                           => n9662);
   clk_r_REG1268_S1 : DFF_X1 port map( D => n3360, CK => CLK, Q => n_3211, QN 
                           => n9661);
   clk_r_REG715_S1 : DFF_X1 port map( D => n3392, CK => CLK, Q => n_3212, QN =>
                           n9660);
   clk_r_REG974_S1 : DFF_X1 port map( D => n3424, CK => CLK, Q => n_3213, QN =>
                           n9659);
   clk_r_REG1355_S1 : DFF_X1 port map( D => n3456, CK => CLK, Q => n_3214, QN 
                           => n9658);
   clk_r_REG1531_S1 : DFF_X1 port map( D => n3488, CK => CLK, Q => n_3215, QN 
                           => n9657);
   clk_r_REG3082_S1 : DFF_X1 port map( D => n3520, CK => CLK, Q => n_3216, QN 
                           => n9656);
   clk_r_REG3154_S1 : DFF_X1 port map( D => n3552, CK => CLK, Q => n_3217, QN 
                           => n9655);
   clk_r_REG2143_S1 : DFF_X1 port map( D => n2569, CK => CLK, Q => n_3218, QN 
                           => n9654);
   clk_r_REG2214_S1 : DFF_X1 port map( D => n2595, CK => CLK, Q => n_3219, QN 
                           => n9653);
   clk_r_REG2290_S1 : DFF_X1 port map( D => n2627, CK => CLK, Q => n_3220, QN 
                           => n9652);
   clk_r_REG2366_S1 : DFF_X1 port map( D => n2659, CK => CLK, Q => n_3221, QN 
                           => n9651);
   clk_r_REG2447_S1 : DFF_X1 port map( D => n2691, CK => CLK, Q => n_3222, QN 
                           => n9650);
   clk_r_REG2525_S1 : DFF_X1 port map( D => n2723, CK => CLK, Q => n_3223, QN 
                           => n9649);
   clk_r_REG2605_S1 : DFF_X1 port map( D => n2755, CK => CLK, Q => n_3224, QN 
                           => n9648);
   clk_r_REG2681_S1 : DFF_X1 port map( D => n2787, CK => CLK, Q => n_3225, QN 
                           => n9647);
   clk_r_REG1841_S1 : DFF_X1 port map( D => n2817, CK => CLK, Q => n_3226, QN 
                           => n9646);
   clk_r_REG1915_S1 : DFF_X1 port map( D => n2849, CK => CLK, Q => n_3227, QN 
                           => n9645);
   clk_r_REG1990_S1 : DFF_X1 port map( D => n2881, CK => CLK, Q => n_3228, QN 
                           => n9644);
   clk_r_REG2764_S1 : DFF_X1 port map( D => n2913, CK => CLK, Q => n_3229, QN 
                           => n9643);
   clk_r_REG2839_S1 : DFF_X1 port map( D => n2945, CK => CLK, Q => n_3230, QN 
                           => n9642);
   clk_r_REG2911_S1 : DFF_X1 port map( D => n2977, CK => CLK, Q => n_3231, QN 
                           => n9641);
   clk_r_REG2061_S1 : DFF_X1 port map( D => n3009, CK => CLK, Q => n_3232, QN 
                           => n9640);
   clk_r_REG2988_S1 : DFF_X1 port map( D => n3041, CK => CLK, Q => n_3233, QN 
                           => n9639);
   clk_r_REG1607_S1 : DFF_X1 port map( D => n3073, CK => CLK, Q => n_3234, QN 
                           => n9638);
   clk_r_REG1684_S1 : DFF_X1 port map( D => n3105, CK => CLK, Q => n_3235, QN 
                           => n9637);
   clk_r_REG1431_S1 : DFF_X1 port map( D => n3137, CK => CLK, Q => n_3236, QN 
                           => n9636);
   clk_r_REG1768_S1 : DFF_X1 port map( D => n3169, CK => CLK, Q => n_3237, QN 
                           => n9635);
   clk_r_REG1047_S1 : DFF_X1 port map( D => n3201, CK => CLK, Q => n_3238, QN 
                           => n9634);
   clk_r_REG1122_S1 : DFF_X1 port map( D => n3233, CK => CLK, Q => n_3239, QN 
                           => n9633);
   clk_r_REG796_S1 : DFF_X1 port map( D => n3265, CK => CLK, Q => n_3240, QN =>
                           n9632);
   clk_r_REG873_S1 : DFF_X1 port map( D => n3297, CK => CLK, Q => n_3241, QN =>
                           n9631);
   clk_r_REG1186_S1 : DFF_X1 port map( D => n3329, CK => CLK, Q => n_3242, QN 
                           => n9630);
   clk_r_REG1266_S1 : DFF_X1 port map( D => n3361, CK => CLK, Q => n_3243, QN 
                           => n9629);
   clk_r_REG713_S1 : DFF_X1 port map( D => n3393, CK => CLK, Q => n_3244, QN =>
                           n9628);
   clk_r_REG972_S1 : DFF_X1 port map( D => n3425, CK => CLK, Q => n_3245, QN =>
                           n9627);
   clk_r_REG1353_S1 : DFF_X1 port map( D => n3457, CK => CLK, Q => n_3246, QN 
                           => n9626);
   clk_r_REG1529_S1 : DFF_X1 port map( D => n3489, CK => CLK, Q => n_3247, QN 
                           => n9625);
   clk_r_REG3080_S1 : DFF_X1 port map( D => n3521, CK => CLK, Q => n_3248, QN 
                           => n9624);
   clk_r_REG3152_S1 : DFF_X1 port map( D => n3553, CK => CLK, Q => n_3249, QN 
                           => n9623);
   clk_r_REG2141_S1 : DFF_X1 port map( D => n2570, CK => CLK, Q => n_3250, QN 
                           => n9622);
   clk_r_REG2226_S1 : DFF_X1 port map( D => n2582, CK => CLK, Q => n_3251, QN 
                           => n9621);
   clk_r_REG2302_S1 : DFF_X1 port map( D => n2614, CK => CLK, Q => n_3252, QN 
                           => n9620);
   clk_r_REG2378_S1 : DFF_X1 port map( D => n2646, CK => CLK, Q => n_3253, QN 
                           => n9619);
   clk_r_REG2459_S1 : DFF_X1 port map( D => n2678, CK => CLK, Q => n_3254, QN 
                           => n9618);
   clk_r_REG2537_S1 : DFF_X1 port map( D => n2710, CK => CLK, Q => n_3255, QN 
                           => n9617);
   clk_r_REG2617_S1 : DFF_X1 port map( D => n2742, CK => CLK, Q => n_3256, QN 
                           => n9616);
   clk_r_REG2693_S1 : DFF_X1 port map( D => n2774, CK => CLK, Q => n_3257, QN 
                           => n9615);
   clk_r_REG1839_S1 : DFF_X1 port map( D => n2818, CK => CLK, Q => n_3258, QN 
                           => n9614);
   clk_r_REG1913_S1 : DFF_X1 port map( D => n2850, CK => CLK, Q => n_3259, QN 
                           => n9613);
   clk_r_REG1988_S1 : DFF_X1 port map( D => n2882, CK => CLK, Q => n_3260, QN 
                           => n9612);
   clk_r_REG2762_S1 : DFF_X1 port map( D => n2914, CK => CLK, Q => n_3261, QN 
                           => n9611);
   clk_r_REG2837_S1 : DFF_X1 port map( D => n2946, CK => CLK, Q => n_3262, QN 
                           => n9610);
   clk_r_REG2909_S1 : DFF_X1 port map( D => n2978, CK => CLK, Q => n_3263, QN 
                           => n9609);
   clk_r_REG2059_S1 : DFF_X1 port map( D => n3010, CK => CLK, Q => n_3264, QN 
                           => n9608);
   clk_r_REG2986_S1 : DFF_X1 port map( D => n3042, CK => CLK, Q => n_3265, QN 
                           => n9607);
   clk_r_REG1605_S1 : DFF_X1 port map( D => n3074, CK => CLK, Q => n_3266, QN 
                           => n9606);
   clk_r_REG1682_S1 : DFF_X1 port map( D => n3106, CK => CLK, Q => n_3267, QN 
                           => n9605);
   clk_r_REG1429_S1 : DFF_X1 port map( D => n3138, CK => CLK, Q => n_3268, QN 
                           => n9604);
   clk_r_REG1766_S1 : DFF_X1 port map( D => n3170, CK => CLK, Q => n_3269, QN 
                           => n9603);
   clk_r_REG1045_S1 : DFF_X1 port map( D => n3202, CK => CLK, Q => n_3270, QN 
                           => n9602);
   clk_r_REG1120_S1 : DFF_X1 port map( D => n3234, CK => CLK, Q => n_3271, QN 
                           => n9601);
   clk_r_REG794_S1 : DFF_X1 port map( D => n3266, CK => CLK, Q => n_3272, QN =>
                           n9600);
   clk_r_REG871_S1 : DFF_X1 port map( D => n3298, CK => CLK, Q => n_3273, QN =>
                           n9599);
   clk_r_REG1184_S1 : DFF_X1 port map( D => n3330, CK => CLK, Q => n_3274, QN 
                           => n9598);
   clk_r_REG1264_S1 : DFF_X1 port map( D => n3362, CK => CLK, Q => n_3275, QN 
                           => n9597);
   clk_r_REG711_S1 : DFF_X1 port map( D => n3394, CK => CLK, Q => n_3276, QN =>
                           n9596);
   clk_r_REG970_S1 : DFF_X1 port map( D => n3426, CK => CLK, Q => n_3277, QN =>
                           n9595);
   clk_r_REG1351_S1 : DFF_X1 port map( D => n3458, CK => CLK, Q => n_3278, QN 
                           => n9594);
   clk_r_REG1527_S1 : DFF_X1 port map( D => n3490, CK => CLK, Q => n_3279, QN 
                           => n9593);
   clk_r_REG3078_S1 : DFF_X1 port map( D => n3522, CK => CLK, Q => n_3280, QN 
                           => n9592);
   clk_r_REG3150_S1 : DFF_X1 port map( D => n3554, CK => CLK, Q => n_3281, QN 
                           => n9591);
   clk_r_REG2139_S1 : DFF_X1 port map( D => n2571, CK => CLK, Q => n_3282, QN 
                           => n9590);
   clk_r_REG2212_S1 : DFF_X1 port map( D => n2596, CK => CLK, Q => n_3283, QN 
                           => n9589);
   clk_r_REG2288_S1 : DFF_X1 port map( D => n2628, CK => CLK, Q => n_3284, QN 
                           => n9588);
   clk_r_REG2364_S1 : DFF_X1 port map( D => n2660, CK => CLK, Q => n_3285, QN 
                           => n9587);
   clk_r_REG2445_S1 : DFF_X1 port map( D => n2692, CK => CLK, Q => n_3286, QN 
                           => n9586);
   clk_r_REG2523_S1 : DFF_X1 port map( D => n2724, CK => CLK, Q => n_3287, QN 
                           => n9585);
   clk_r_REG2603_S1 : DFF_X1 port map( D => n2756, CK => CLK, Q => n_3288, QN 
                           => n9584);
   clk_r_REG2679_S1 : DFF_X1 port map( D => n2788, CK => CLK, Q => n_3289, QN 
                           => n9583);
   clk_r_REG1837_S1 : DFF_X1 port map( D => n2819, CK => CLK, Q => n_3290, QN 
                           => n9582);
   clk_r_REG1911_S1 : DFF_X1 port map( D => n2851, CK => CLK, Q => n_3291, QN 
                           => n9581);
   clk_r_REG1986_S1 : DFF_X1 port map( D => n2883, CK => CLK, Q => n_3292, QN 
                           => n9580);
   clk_r_REG2760_S1 : DFF_X1 port map( D => n2915, CK => CLK, Q => n_3293, QN 
                           => n9579);
   clk_r_REG2835_S1 : DFF_X1 port map( D => n2947, CK => CLK, Q => n_3294, QN 
                           => n9578);
   clk_r_REG2907_S1 : DFF_X1 port map( D => n2979, CK => CLK, Q => n_3295, QN 
                           => n9577);
   clk_r_REG2057_S1 : DFF_X1 port map( D => n3011, CK => CLK, Q => n_3296, QN 
                           => n9576);
   clk_r_REG2984_S1 : DFF_X1 port map( D => n3043, CK => CLK, Q => n_3297, QN 
                           => n9575);
   clk_r_REG1603_S1 : DFF_X1 port map( D => n3075, CK => CLK, Q => n_3298, QN 
                           => n9574);
   clk_r_REG1680_S1 : DFF_X1 port map( D => n3107, CK => CLK, Q => n_3299, QN 
                           => n9573);
   clk_r_REG1427_S1 : DFF_X1 port map( D => n3139, CK => CLK, Q => n_3300, QN 
                           => n9572);
   clk_r_REG1764_S1 : DFF_X1 port map( D => n3171, CK => CLK, Q => n_3301, QN 
                           => n9571);
   clk_r_REG1043_S1 : DFF_X1 port map( D => n3203, CK => CLK, Q => n_3302, QN 
                           => n9570);
   clk_r_REG1118_S1 : DFF_X1 port map( D => n3235, CK => CLK, Q => n_3303, QN 
                           => n9569);
   clk_r_REG792_S1 : DFF_X1 port map( D => n3267, CK => CLK, Q => n_3304, QN =>
                           n9568);
   clk_r_REG869_S1 : DFF_X1 port map( D => n3299, CK => CLK, Q => n_3305, QN =>
                           n9567);
   clk_r_REG1182_S1 : DFF_X1 port map( D => n3331, CK => CLK, Q => n_3306, QN 
                           => n9566);
   clk_r_REG1262_S1 : DFF_X1 port map( D => n3363, CK => CLK, Q => n_3307, QN 
                           => n9565);
   clk_r_REG709_S1 : DFF_X1 port map( D => n3395, CK => CLK, Q => n_3308, QN =>
                           n9564);
   clk_r_REG968_S1 : DFF_X1 port map( D => n3427, CK => CLK, Q => n_3309, QN =>
                           n9563);
   clk_r_REG1349_S1 : DFF_X1 port map( D => n3459, CK => CLK, Q => n_3310, QN 
                           => n9562);
   clk_r_REG1525_S1 : DFF_X1 port map( D => n3491, CK => CLK, Q => n_3311, QN 
                           => n9561);
   clk_r_REG3076_S1 : DFF_X1 port map( D => n3523, CK => CLK, Q => n_3312, QN 
                           => n9560);
   clk_r_REG3148_S1 : DFF_X1 port map( D => n3555, CK => CLK, Q => n_3313, QN 
                           => n9559);
   clk_r_REG2137_S1 : DFF_X1 port map( D => n2572, CK => CLK, Q => n_3314, QN 
                           => n9558);
   clk_r_REG2210_S1 : DFF_X1 port map( D => n2597, CK => CLK, Q => n_3315, QN 
                           => n9557);
   clk_r_REG2286_S1 : DFF_X1 port map( D => n2629, CK => CLK, Q => n_3316, QN 
                           => n9556);
   clk_r_REG2362_S1 : DFF_X1 port map( D => n2661, CK => CLK, Q => n_3317, QN 
                           => n9555);
   clk_r_REG2443_S1 : DFF_X1 port map( D => n2693, CK => CLK, Q => n_3318, QN 
                           => n9554);
   clk_r_REG2521_S1 : DFF_X1 port map( D => n2725, CK => CLK, Q => n_3319, QN 
                           => n9553);
   clk_r_REG2601_S1 : DFF_X1 port map( D => n2757, CK => CLK, Q => n_3320, QN 
                           => n9552);
   clk_r_REG2677_S1 : DFF_X1 port map( D => n2789, CK => CLK, Q => n_3321, QN 
                           => n9551);
   clk_r_REG1835_S1 : DFF_X1 port map( D => n2820, CK => CLK, Q => n_3322, QN 
                           => n9550);
   clk_r_REG1909_S1 : DFF_X1 port map( D => n2852, CK => CLK, Q => n_3323, QN 
                           => n9549);
   clk_r_REG1984_S1 : DFF_X1 port map( D => n2884, CK => CLK, Q => n_3324, QN 
                           => n9548);
   clk_r_REG2758_S1 : DFF_X1 port map( D => n2916, CK => CLK, Q => n_3325, QN 
                           => n9547);
   clk_r_REG2833_S1 : DFF_X1 port map( D => n2948, CK => CLK, Q => n_3326, QN 
                           => n9546);
   clk_r_REG2905_S1 : DFF_X1 port map( D => n2980, CK => CLK, Q => n_3327, QN 
                           => n9545);
   clk_r_REG2055_S1 : DFF_X1 port map( D => n3012, CK => CLK, Q => n_3328, QN 
                           => n9544);
   clk_r_REG2982_S1 : DFF_X1 port map( D => n3044, CK => CLK, Q => n_3329, QN 
                           => n9543);
   clk_r_REG1601_S1 : DFF_X1 port map( D => n3076, CK => CLK, Q => n_3330, QN 
                           => n9542);
   clk_r_REG1678_S1 : DFF_X1 port map( D => n3108, CK => CLK, Q => n_3331, QN 
                           => n9541);
   clk_r_REG1425_S1 : DFF_X1 port map( D => n3140, CK => CLK, Q => n_3332, QN 
                           => n9540);
   clk_r_REG1762_S1 : DFF_X1 port map( D => n3172, CK => CLK, Q => n_3333, QN 
                           => n9539);
   clk_r_REG1041_S1 : DFF_X1 port map( D => n3204, CK => CLK, Q => n_3334, QN 
                           => n9538);
   clk_r_REG1116_S1 : DFF_X1 port map( D => n3236, CK => CLK, Q => n_3335, QN 
                           => n9537);
   clk_r_REG790_S1 : DFF_X1 port map( D => n3268, CK => CLK, Q => n_3336, QN =>
                           n9536);
   clk_r_REG867_S1 : DFF_X1 port map( D => n3300, CK => CLK, Q => n_3337, QN =>
                           n9535);
   clk_r_REG1180_S1 : DFF_X1 port map( D => n3332, CK => CLK, Q => n_3338, QN 
                           => n9534);
   clk_r_REG1260_S1 : DFF_X1 port map( D => n3364, CK => CLK, Q => n_3339, QN 
                           => n9533);
   clk_r_REG707_S1 : DFF_X1 port map( D => n3396, CK => CLK, Q => n_3340, QN =>
                           n9532);
   clk_r_REG966_S1 : DFF_X1 port map( D => n3428, CK => CLK, Q => n_3341, QN =>
                           n9531);
   clk_r_REG1347_S1 : DFF_X1 port map( D => n3460, CK => CLK, Q => n_3342, QN 
                           => n9530);
   clk_r_REG1523_S1 : DFF_X1 port map( D => n3492, CK => CLK, Q => n_3343, QN 
                           => n9529);
   clk_r_REG3074_S1 : DFF_X1 port map( D => n3524, CK => CLK, Q => n_3344, QN 
                           => n9528);
   clk_r_REG3146_S1 : DFF_X1 port map( D => n3556, CK => CLK, Q => n_3345, QN 
                           => n9527);
   clk_r_REG2135_S1 : DFF_X1 port map( D => n2573, CK => CLK, Q => n_3346, QN 
                           => n9526);
   clk_r_REG2208_S1 : DFF_X1 port map( D => n2598, CK => CLK, Q => n_3347, QN 
                           => n9525);
   clk_r_REG2284_S1 : DFF_X1 port map( D => n2630, CK => CLK, Q => n_3348, QN 
                           => n9524);
   clk_r_REG2360_S1 : DFF_X1 port map( D => n2662, CK => CLK, Q => n_3349, QN 
                           => n9523);
   clk_r_REG2441_S1 : DFF_X1 port map( D => n2694, CK => CLK, Q => n_3350, QN 
                           => n9522);
   clk_r_REG2519_S1 : DFF_X1 port map( D => n2726, CK => CLK, Q => n_3351, QN 
                           => n9521);
   clk_r_REG2599_S1 : DFF_X1 port map( D => n2758, CK => CLK, Q => n_3352, QN 
                           => n9520);
   clk_r_REG2675_S1 : DFF_X1 port map( D => n2790, CK => CLK, Q => n_3353, QN 
                           => n9519);
   clk_r_REG1833_S1 : DFF_X1 port map( D => n2821, CK => CLK, Q => n_3354, QN 
                           => n9518);
   clk_r_REG1907_S1 : DFF_X1 port map( D => n2853, CK => CLK, Q => n_3355, QN 
                           => n9517);
   clk_r_REG1982_S1 : DFF_X1 port map( D => n2885, CK => CLK, Q => n_3356, QN 
                           => n9516);
   clk_r_REG2756_S1 : DFF_X1 port map( D => n2917, CK => CLK, Q => n_3357, QN 
                           => n9515);
   clk_r_REG2831_S1 : DFF_X1 port map( D => n2949, CK => CLK, Q => n_3358, QN 
                           => n9514);
   clk_r_REG2903_S1 : DFF_X1 port map( D => n2981, CK => CLK, Q => n_3359, QN 
                           => n9513);
   clk_r_REG2053_S1 : DFF_X1 port map( D => n3013, CK => CLK, Q => n_3360, QN 
                           => n9512);
   clk_r_REG2980_S1 : DFF_X1 port map( D => n3045, CK => CLK, Q => n_3361, QN 
                           => n9511);
   clk_r_REG1599_S1 : DFF_X1 port map( D => n3077, CK => CLK, Q => n_3362, QN 
                           => n9510);
   clk_r_REG1676_S1 : DFF_X1 port map( D => n3109, CK => CLK, Q => n_3363, QN 
                           => n9509);
   clk_r_REG1423_S1 : DFF_X1 port map( D => n3141, CK => CLK, Q => n_3364, QN 
                           => n9508);
   clk_r_REG1760_S1 : DFF_X1 port map( D => n3173, CK => CLK, Q => n_3365, QN 
                           => n9507);
   clk_r_REG1039_S1 : DFF_X1 port map( D => n3205, CK => CLK, Q => n_3366, QN 
                           => n9506);
   clk_r_REG1114_S1 : DFF_X1 port map( D => n3237, CK => CLK, Q => n_3367, QN 
                           => n9505);
   clk_r_REG788_S1 : DFF_X1 port map( D => n3269, CK => CLK, Q => n_3368, QN =>
                           n9504);
   clk_r_REG865_S1 : DFF_X1 port map( D => n3301, CK => CLK, Q => n_3369, QN =>
                           n9503);
   clk_r_REG1178_S1 : DFF_X1 port map( D => n3333, CK => CLK, Q => n_3370, QN 
                           => n9502);
   clk_r_REG1258_S1 : DFF_X1 port map( D => n3365, CK => CLK, Q => n_3371, QN 
                           => n9501);
   clk_r_REG705_S1 : DFF_X1 port map( D => n3397, CK => CLK, Q => n_3372, QN =>
                           n9500);
   clk_r_REG964_S1 : DFF_X1 port map( D => n3429, CK => CLK, Q => n_3373, QN =>
                           n9499);
   clk_r_REG1345_S1 : DFF_X1 port map( D => n3461, CK => CLK, Q => n_3374, QN 
                           => n9498);
   clk_r_REG1521_S1 : DFF_X1 port map( D => n3493, CK => CLK, Q => n_3375, QN 
                           => n9497);
   clk_r_REG3072_S1 : DFF_X1 port map( D => n3525, CK => CLK, Q => n_3376, QN 
                           => n9496);
   clk_r_REG3144_S1 : DFF_X1 port map( D => n3557, CK => CLK, Q => n_3377, QN 
                           => n9495);
   clk_r_REG2133_S1 : DFF_X1 port map( D => n2574, CK => CLK, Q => n_3378, QN 
                           => n9494);
   clk_r_REG2206_S1 : DFF_X1 port map( D => n2599, CK => CLK, Q => n_3379, QN 
                           => n9493);
   clk_r_REG2282_S1 : DFF_X1 port map( D => n2631, CK => CLK, Q => n_3380, QN 
                           => n9492);
   clk_r_REG2358_S1 : DFF_X1 port map( D => n2663, CK => CLK, Q => n_3381, QN 
                           => n9491);
   clk_r_REG2439_S1 : DFF_X1 port map( D => n2695, CK => CLK, Q => n_3382, QN 
                           => n9490);
   clk_r_REG2517_S1 : DFF_X1 port map( D => n2727, CK => CLK, Q => n_3383, QN 
                           => n9489);
   clk_r_REG2597_S1 : DFF_X1 port map( D => n2759, CK => CLK, Q => n_3384, QN 
                           => n9488);
   clk_r_REG2673_S1 : DFF_X1 port map( D => n2791, CK => CLK, Q => n_3385, QN 
                           => n9487);
   clk_r_REG1831_S1 : DFF_X1 port map( D => n2822, CK => CLK, Q => n_3386, QN 
                           => n9486);
   clk_r_REG1905_S1 : DFF_X1 port map( D => n2854, CK => CLK, Q => n_3387, QN 
                           => n9485);
   clk_r_REG1980_S1 : DFF_X1 port map( D => n2886, CK => CLK, Q => n_3388, QN 
                           => n9484);
   clk_r_REG2754_S1 : DFF_X1 port map( D => n2918, CK => CLK, Q => n_3389, QN 
                           => n9483);
   clk_r_REG2829_S1 : DFF_X1 port map( D => n2950, CK => CLK, Q => n_3390, QN 
                           => n9482);
   clk_r_REG2901_S1 : DFF_X1 port map( D => n2982, CK => CLK, Q => n_3391, QN 
                           => n9481);
   clk_r_REG2051_S1 : DFF_X1 port map( D => n3014, CK => CLK, Q => n_3392, QN 
                           => n9480);
   clk_r_REG2978_S1 : DFF_X1 port map( D => n3046, CK => CLK, Q => n_3393, QN 
                           => n9479);
   clk_r_REG1597_S1 : DFF_X1 port map( D => n3078, CK => CLK, Q => n_3394, QN 
                           => n9478);
   clk_r_REG1674_S1 : DFF_X1 port map( D => n3110, CK => CLK, Q => n_3395, QN 
                           => n9477);
   clk_r_REG1421_S1 : DFF_X1 port map( D => n3142, CK => CLK, Q => n_3396, QN 
                           => n9476);
   clk_r_REG1758_S1 : DFF_X1 port map( D => n3174, CK => CLK, Q => n_3397, QN 
                           => n9475);
   clk_r_REG1037_S1 : DFF_X1 port map( D => n3206, CK => CLK, Q => n_3398, QN 
                           => n9474);
   clk_r_REG1112_S1 : DFF_X1 port map( D => n3238, CK => CLK, Q => n_3399, QN 
                           => n9473);
   clk_r_REG786_S1 : DFF_X1 port map( D => n3270, CK => CLK, Q => n_3400, QN =>
                           n9472);
   clk_r_REG863_S1 : DFF_X1 port map( D => n3302, CK => CLK, Q => n_3401, QN =>
                           n9471);
   clk_r_REG1176_S1 : DFF_X1 port map( D => n3334, CK => CLK, Q => n_3402, QN 
                           => n9470);
   clk_r_REG1256_S1 : DFF_X1 port map( D => n3366, CK => CLK, Q => n_3403, QN 
                           => n9469);
   clk_r_REG703_S1 : DFF_X1 port map( D => n3398, CK => CLK, Q => n_3404, QN =>
                           n9468);
   clk_r_REG962_S1 : DFF_X1 port map( D => n3430, CK => CLK, Q => n_3405, QN =>
                           n9467);
   clk_r_REG1343_S1 : DFF_X1 port map( D => n3462, CK => CLK, Q => n_3406, QN 
                           => n9466);
   clk_r_REG1519_S1 : DFF_X1 port map( D => n3494, CK => CLK, Q => n_3407, QN 
                           => n9465);
   clk_r_REG3070_S1 : DFF_X1 port map( D => n3526, CK => CLK, Q => n_3408, QN 
                           => n9464);
   clk_r_REG3142_S1 : DFF_X1 port map( D => n3558, CK => CLK, Q => n_3409, QN 
                           => n9463);
   clk_r_REG2131_S1 : DFF_X1 port map( D => n2575, CK => CLK, Q => n_3410, QN 
                           => n9462);
   clk_r_REG2204_S1 : DFF_X1 port map( D => n2600, CK => CLK, Q => n_3411, QN 
                           => n9461);
   clk_r_REG2280_S1 : DFF_X1 port map( D => n2632, CK => CLK, Q => n_3412, QN 
                           => n9460);
   clk_r_REG2356_S1 : DFF_X1 port map( D => n2664, CK => CLK, Q => n_3413, QN 
                           => n9459);
   clk_r_REG2437_S1 : DFF_X1 port map( D => n2696, CK => CLK, Q => n_3414, QN 
                           => n9458);
   clk_r_REG2515_S1 : DFF_X1 port map( D => n2728, CK => CLK, Q => n_3415, QN 
                           => n9457);
   clk_r_REG2595_S1 : DFF_X1 port map( D => n2760, CK => CLK, Q => n_3416, QN 
                           => n9456);
   clk_r_REG2671_S1 : DFF_X1 port map( D => n2792, CK => CLK, Q => n_3417, QN 
                           => n9455);
   clk_r_REG1829_S1 : DFF_X1 port map( D => n2823, CK => CLK, Q => n_3418, QN 
                           => n9454);
   clk_r_REG1903_S1 : DFF_X1 port map( D => n2855, CK => CLK, Q => n_3419, QN 
                           => n9453);
   clk_r_REG1978_S1 : DFF_X1 port map( D => n2887, CK => CLK, Q => n_3420, QN 
                           => n9452);
   clk_r_REG2752_S1 : DFF_X1 port map( D => n2919, CK => CLK, Q => n_3421, QN 
                           => n9451);
   clk_r_REG2827_S1 : DFF_X1 port map( D => n2951, CK => CLK, Q => n_3422, QN 
                           => n9450);
   clk_r_REG2899_S1 : DFF_X1 port map( D => n2983, CK => CLK, Q => n_3423, QN 
                           => n9449);
   clk_r_REG2049_S1 : DFF_X1 port map( D => n3015, CK => CLK, Q => n_3424, QN 
                           => n9448);
   clk_r_REG2976_S1 : DFF_X1 port map( D => n3047, CK => CLK, Q => n_3425, QN 
                           => n9447);
   clk_r_REG1595_S1 : DFF_X1 port map( D => n3079, CK => CLK, Q => n_3426, QN 
                           => n9446);
   clk_r_REG1672_S1 : DFF_X1 port map( D => n3111, CK => CLK, Q => n_3427, QN 
                           => n9445);
   clk_r_REG1419_S1 : DFF_X1 port map( D => n3143, CK => CLK, Q => n_3428, QN 
                           => n9444);
   clk_r_REG1756_S1 : DFF_X1 port map( D => n3175, CK => CLK, Q => n_3429, QN 
                           => n9443);
   clk_r_REG1035_S1 : DFF_X1 port map( D => n3207, CK => CLK, Q => n_3430, QN 
                           => n9442);
   clk_r_REG1110_S1 : DFF_X1 port map( D => n3239, CK => CLK, Q => n_3431, QN 
                           => n9441);
   clk_r_REG784_S1 : DFF_X1 port map( D => n3271, CK => CLK, Q => n_3432, QN =>
                           n9440);
   clk_r_REG861_S1 : DFF_X1 port map( D => n3303, CK => CLK, Q => n_3433, QN =>
                           n9439);
   clk_r_REG1174_S1 : DFF_X1 port map( D => n3335, CK => CLK, Q => n_3434, QN 
                           => n9438);
   clk_r_REG1254_S1 : DFF_X1 port map( D => n3367, CK => CLK, Q => n_3435, QN 
                           => n9437);
   clk_r_REG701_S1 : DFF_X1 port map( D => n3399, CK => CLK, Q => n_3436, QN =>
                           n9436);
   clk_r_REG960_S1 : DFF_X1 port map( D => n3431, CK => CLK, Q => n_3437, QN =>
                           n9435);
   clk_r_REG1341_S1 : DFF_X1 port map( D => n3463, CK => CLK, Q => n_3438, QN 
                           => n9434);
   clk_r_REG1517_S1 : DFF_X1 port map( D => n3495, CK => CLK, Q => n_3439, QN 
                           => n9433);
   clk_r_REG3068_S1 : DFF_X1 port map( D => n3527, CK => CLK, Q => n_3440, QN 
                           => n9432);
   clk_r_REG3140_S1 : DFF_X1 port map( D => n3559, CK => CLK, Q => n_3441, QN 
                           => n9431);
   clk_r_REG2129_S1 : DFF_X1 port map( D => n2576, CK => CLK, Q => n_3442, QN 
                           => n9430);
   clk_r_REG2202_S1 : DFF_X1 port map( D => n2601, CK => CLK, Q => n_3443, QN 
                           => n9429);
   clk_r_REG2278_S1 : DFF_X1 port map( D => n2633, CK => CLK, Q => n_3444, QN 
                           => n9428);
   clk_r_REG2354_S1 : DFF_X1 port map( D => n2665, CK => CLK, Q => n_3445, QN 
                           => n9427);
   clk_r_REG2435_S1 : DFF_X1 port map( D => n2697, CK => CLK, Q => n_3446, QN 
                           => n9426);
   clk_r_REG2513_S1 : DFF_X1 port map( D => n2729, CK => CLK, Q => n_3447, QN 
                           => n9425);
   clk_r_REG2593_S1 : DFF_X1 port map( D => n2761, CK => CLK, Q => n_3448, QN 
                           => n9424);
   clk_r_REG2669_S1 : DFF_X1 port map( D => n2793, CK => CLK, Q => n_3449, QN 
                           => n9423);
   clk_r_REG1827_S1 : DFF_X1 port map( D => n2824, CK => CLK, Q => n_3450, QN 
                           => n9422);
   clk_r_REG1901_S1 : DFF_X1 port map( D => n2856, CK => CLK, Q => n_3451, QN 
                           => n9421);
   clk_r_REG1976_S1 : DFF_X1 port map( D => n2888, CK => CLK, Q => n_3452, QN 
                           => n9420);
   clk_r_REG2750_S1 : DFF_X1 port map( D => n2920, CK => CLK, Q => n_3453, QN 
                           => n9419);
   clk_r_REG2825_S1 : DFF_X1 port map( D => n2952, CK => CLK, Q => n_3454, QN 
                           => n9418);
   clk_r_REG2897_S1 : DFF_X1 port map( D => n2984, CK => CLK, Q => n_3455, QN 
                           => n9417);
   clk_r_REG2047_S1 : DFF_X1 port map( D => n3016, CK => CLK, Q => n_3456, QN 
                           => n9416);
   clk_r_REG2974_S1 : DFF_X1 port map( D => n3048, CK => CLK, Q => n_3457, QN 
                           => n9415);
   clk_r_REG1593_S1 : DFF_X1 port map( D => n3080, CK => CLK, Q => n_3458, QN 
                           => n9414);
   clk_r_REG1670_S1 : DFF_X1 port map( D => n3112, CK => CLK, Q => n_3459, QN 
                           => n9413);
   clk_r_REG1417_S1 : DFF_X1 port map( D => n3144, CK => CLK, Q => n_3460, QN 
                           => n9412);
   clk_r_REG1754_S1 : DFF_X1 port map( D => n3176, CK => CLK, Q => n_3461, QN 
                           => n9411);
   clk_r_REG1033_S1 : DFF_X1 port map( D => n3208, CK => CLK, Q => n_3462, QN 
                           => n9410);
   clk_r_REG1108_S1 : DFF_X1 port map( D => n3240, CK => CLK, Q => n_3463, QN 
                           => n9409);
   clk_r_REG782_S1 : DFF_X1 port map( D => n3272, CK => CLK, Q => n_3464, QN =>
                           n9408);
   clk_r_REG859_S1 : DFF_X1 port map( D => n3304, CK => CLK, Q => n_3465, QN =>
                           n9407);
   clk_r_REG1172_S1 : DFF_X1 port map( D => n3336, CK => CLK, Q => n_3466, QN 
                           => n9406);
   clk_r_REG1252_S1 : DFF_X1 port map( D => n3368, CK => CLK, Q => n_3467, QN 
                           => n9405);
   clk_r_REG699_S1 : DFF_X1 port map( D => n3400, CK => CLK, Q => n_3468, QN =>
                           n9404);
   clk_r_REG958_S1 : DFF_X1 port map( D => n3432, CK => CLK, Q => n_3469, QN =>
                           n9403);
   clk_r_REG1339_S1 : DFF_X1 port map( D => n3464, CK => CLK, Q => n_3470, QN 
                           => n9402);
   clk_r_REG1515_S1 : DFF_X1 port map( D => n3496, CK => CLK, Q => n_3471, QN 
                           => n9401);
   clk_r_REG3066_S1 : DFF_X1 port map( D => n3528, CK => CLK, Q => n_3472, QN 
                           => n9400);
   clk_r_REG3138_S1 : DFF_X1 port map( D => n3560, CK => CLK, Q => n_3473, QN 
                           => n9399);
   clk_r_REG2127_S1 : DFF_X1 port map( D => n2577, CK => CLK, Q => n_3474, QN 
                           => n9398);
   clk_r_REG2224_S1 : DFF_X1 port map( D => n2581, CK => CLK, Q => n_3475, QN 
                           => n9397);
   clk_r_REG2300_S1 : DFF_X1 port map( D => n2613, CK => CLK, Q => n_3476, QN 
                           => n9396);
   clk_r_REG2376_S1 : DFF_X1 port map( D => n2645, CK => CLK, Q => n_3477, QN 
                           => n9395);
   clk_r_REG2457_S1 : DFF_X1 port map( D => n2677, CK => CLK, Q => n_3478, QN 
                           => n9394);
   clk_r_REG2535_S1 : DFF_X1 port map( D => n2709, CK => CLK, Q => n_3479, QN 
                           => n9393);
   clk_r_REG2615_S1 : DFF_X1 port map( D => n2741, CK => CLK, Q => n_3480, QN 
                           => n9392);
   clk_r_REG2691_S1 : DFF_X1 port map( D => n2773, CK => CLK, Q => n_3481, QN 
                           => n9391);
   clk_r_REG1825_S1 : DFF_X1 port map( D => n2825, CK => CLK, Q => n_3482, QN 
                           => n9390);
   clk_r_REG1899_S1 : DFF_X1 port map( D => n2857, CK => CLK, Q => n_3483, QN 
                           => n9389);
   clk_r_REG1974_S1 : DFF_X1 port map( D => n2889, CK => CLK, Q => n_3484, QN 
                           => n9388);
   clk_r_REG2748_S1 : DFF_X1 port map( D => n2921, CK => CLK, Q => n_3485, QN 
                           => n9387);
   clk_r_REG2823_S1 : DFF_X1 port map( D => n2953, CK => CLK, Q => n_3486, QN 
                           => n9386);
   clk_r_REG2895_S1 : DFF_X1 port map( D => n2985, CK => CLK, Q => n_3487, QN 
                           => n9385);
   clk_r_REG2045_S1 : DFF_X1 port map( D => n3017, CK => CLK, Q => n_3488, QN 
                           => n9384);
   clk_r_REG2972_S1 : DFF_X1 port map( D => n3049, CK => CLK, Q => n_3489, QN 
                           => n9383);
   clk_r_REG1591_S1 : DFF_X1 port map( D => n3081, CK => CLK, Q => n_3490, QN 
                           => n9382);
   clk_r_REG1668_S1 : DFF_X1 port map( D => n3113, CK => CLK, Q => n_3491, QN 
                           => n9381);
   clk_r_REG1415_S1 : DFF_X1 port map( D => n3145, CK => CLK, Q => n_3492, QN 
                           => n9380);
   clk_r_REG1752_S1 : DFF_X1 port map( D => n3177, CK => CLK, Q => n_3493, QN 
                           => n9379);
   clk_r_REG1031_S1 : DFF_X1 port map( D => n3209, CK => CLK, Q => n_3494, QN 
                           => n9378);
   clk_r_REG1106_S1 : DFF_X1 port map( D => n3241, CK => CLK, Q => n_3495, QN 
                           => n9377);
   clk_r_REG780_S1 : DFF_X1 port map( D => n3273, CK => CLK, Q => n_3496, QN =>
                           n9376);
   clk_r_REG857_S1 : DFF_X1 port map( D => n3305, CK => CLK, Q => n_3497, QN =>
                           n9375);
   clk_r_REG1170_S1 : DFF_X1 port map( D => n3337, CK => CLK, Q => n_3498, QN 
                           => n9374);
   clk_r_REG1250_S1 : DFF_X1 port map( D => n3369, CK => CLK, Q => n_3499, QN 
                           => n9373);
   clk_r_REG697_S1 : DFF_X1 port map( D => n3401, CK => CLK, Q => n_3500, QN =>
                           n9372);
   clk_r_REG956_S1 : DFF_X1 port map( D => n3433, CK => CLK, Q => n_3501, QN =>
                           n9371);
   clk_r_REG1337_S1 : DFF_X1 port map( D => n3465, CK => CLK, Q => n_3502, QN 
                           => n9370);
   clk_r_REG1513_S1 : DFF_X1 port map( D => n3497, CK => CLK, Q => n_3503, QN 
                           => n9369);
   clk_r_REG3064_S1 : DFF_X1 port map( D => n3529, CK => CLK, Q => n_3504, QN 
                           => n9368);
   clk_r_REG3136_S1 : DFF_X1 port map( D => n3561, CK => CLK, Q => n_3505, QN 
                           => n9367);
   clk_r_REG2125_S1 : DFF_X1 port map( D => n2578, CK => CLK, Q => n_3506, QN 
                           => n9366);
   clk_r_REG2200_S1 : DFF_X1 port map( D => n2602, CK => CLK, Q => n_3507, QN 
                           => n9365);
   clk_r_REG2276_S1 : DFF_X1 port map( D => n2634, CK => CLK, Q => n_3508, QN 
                           => n9364);
   clk_r_REG2352_S1 : DFF_X1 port map( D => n2666, CK => CLK, Q => n_3509, QN 
                           => n9363);
   clk_r_REG2433_S1 : DFF_X1 port map( D => n2698, CK => CLK, Q => n_3510, QN 
                           => n9362);
   clk_r_REG2511_S1 : DFF_X1 port map( D => n2730, CK => CLK, Q => n_3511, QN 
                           => n9361);
   clk_r_REG2591_S1 : DFF_X1 port map( D => n2762, CK => CLK, Q => n_3512, QN 
                           => n9360);
   clk_r_REG2667_S1 : DFF_X1 port map( D => n2794, CK => CLK, Q => n_3513, QN 
                           => n9359);
   clk_r_REG1823_S1 : DFF_X1 port map( D => n2826, CK => CLK, Q => n_3514, QN 
                           => n9358);
   clk_r_REG1897_S1 : DFF_X1 port map( D => n2858, CK => CLK, Q => n_3515, QN 
                           => n9357);
   clk_r_REG1972_S1 : DFF_X1 port map( D => n2890, CK => CLK, Q => n_3516, QN 
                           => n9356);
   clk_r_REG2746_S1 : DFF_X1 port map( D => n2922, CK => CLK, Q => n_3517, QN 
                           => n9355);
   clk_r_REG2821_S1 : DFF_X1 port map( D => n2954, CK => CLK, Q => n_3518, QN 
                           => n9354);
   clk_r_REG2893_S1 : DFF_X1 port map( D => n2986, CK => CLK, Q => n_3519, QN 
                           => n9353);
   clk_r_REG2043_S1 : DFF_X1 port map( D => n3018, CK => CLK, Q => n_3520, QN 
                           => n9352);
   clk_r_REG2970_S1 : DFF_X1 port map( D => n3050, CK => CLK, Q => n_3521, QN 
                           => n9351);
   clk_r_REG1589_S1 : DFF_X1 port map( D => n3082, CK => CLK, Q => n_3522, QN 
                           => n9350);
   clk_r_REG1666_S1 : DFF_X1 port map( D => n3114, CK => CLK, Q => n_3523, QN 
                           => n9349);
   clk_r_REG1413_S1 : DFF_X1 port map( D => n3146, CK => CLK, Q => n_3524, QN 
                           => n9348);
   clk_r_REG1750_S1 : DFF_X1 port map( D => n3178, CK => CLK, Q => n_3525, QN 
                           => n9347);
   clk_r_REG1029_S1 : DFF_X1 port map( D => n3210, CK => CLK, Q => n_3526, QN 
                           => n9346);
   clk_r_REG1104_S1 : DFF_X1 port map( D => n3242, CK => CLK, Q => n_3527, QN 
                           => n9345);
   clk_r_REG778_S1 : DFF_X1 port map( D => n3274, CK => CLK, Q => n_3528, QN =>
                           n9344);
   clk_r_REG855_S1 : DFF_X1 port map( D => n3306, CK => CLK, Q => n_3529, QN =>
                           n9343);
   clk_r_REG1168_S1 : DFF_X1 port map( D => n3338, CK => CLK, Q => n_3530, QN 
                           => n9342);
   clk_r_REG1248_S1 : DFF_X1 port map( D => n3370, CK => CLK, Q => n_3531, QN 
                           => n9341);
   clk_r_REG695_S1 : DFF_X1 port map( D => n3402, CK => CLK, Q => n_3532, QN =>
                           n9340);
   clk_r_REG954_S1 : DFF_X1 port map( D => n3434, CK => CLK, Q => n_3533, QN =>
                           n9339);
   clk_r_REG1335_S1 : DFF_X1 port map( D => n3466, CK => CLK, Q => n_3534, QN 
                           => n9338);
   clk_r_REG1511_S1 : DFF_X1 port map( D => n3498, CK => CLK, Q => n_3535, QN 
                           => n9337);
   clk_r_REG3062_S1 : DFF_X1 port map( D => n3530, CK => CLK, Q => n_3536, QN 
                           => n9336);
   clk_r_REG3134_S1 : DFF_X1 port map( D => n3562, CK => CLK, Q => n_3537, QN 
                           => n9335);
   clk_r_REG2123_S1 : DFF_X1 port map( D => n2579, CK => CLK, Q => n_3538, QN 
                           => n9334);
   clk_r_REG2198_S1 : DFF_X1 port map( D => n2603, CK => CLK, Q => n_3539, QN 
                           => n9333);
   clk_r_REG2274_S1 : DFF_X1 port map( D => n2635, CK => CLK, Q => n_3540, QN 
                           => n9332);
   clk_r_REG2350_S1 : DFF_X1 port map( D => n2667, CK => CLK, Q => n_3541, QN 
                           => n9331);
   clk_r_REG2431_S1 : DFF_X1 port map( D => n2699, CK => CLK, Q => n_3542, QN 
                           => n9330);
   clk_r_REG2509_S1 : DFF_X1 port map( D => n2731, CK => CLK, Q => n_3543, QN 
                           => n9329);
   clk_r_REG2589_S1 : DFF_X1 port map( D => n2763, CK => CLK, Q => n_3544, QN 
                           => n9328);
   clk_r_REG2665_S1 : DFF_X1 port map( D => n2795, CK => CLK, Q => n_3545, QN 
                           => n9327);
   clk_r_REG1821_S1 : DFF_X1 port map( D => n2827, CK => CLK, Q => n_3546, QN 
                           => n9326);
   clk_r_REG1895_S1 : DFF_X1 port map( D => n2859, CK => CLK, Q => n_3547, QN 
                           => n9325);
   clk_r_REG1970_S1 : DFF_X1 port map( D => n2891, CK => CLK, Q => n_3548, QN 
                           => n9324);
   clk_r_REG2744_S1 : DFF_X1 port map( D => n2923, CK => CLK, Q => n_3549, QN 
                           => n9323);
   clk_r_REG2819_S1 : DFF_X1 port map( D => n2955, CK => CLK, Q => n_3550, QN 
                           => n9322);
   clk_r_REG2891_S1 : DFF_X1 port map( D => n2987, CK => CLK, Q => n_3551, QN 
                           => n9321);
   clk_r_REG2041_S1 : DFF_X1 port map( D => n3019, CK => CLK, Q => n_3552, QN 
                           => n9320);
   clk_r_REG2968_S1 : DFF_X1 port map( D => n3051, CK => CLK, Q => n_3553, QN 
                           => n9319);
   clk_r_REG1587_S1 : DFF_X1 port map( D => n3083, CK => CLK, Q => n_3554, QN 
                           => n9318);
   clk_r_REG1664_S1 : DFF_X1 port map( D => n3115, CK => CLK, Q => n_3555, QN 
                           => n9317);
   clk_r_REG1411_S1 : DFF_X1 port map( D => n3147, CK => CLK, Q => n_3556, QN 
                           => n9316);
   clk_r_REG1748_S1 : DFF_X1 port map( D => n3179, CK => CLK, Q => n_3557, QN 
                           => n9315);
   clk_r_REG1027_S1 : DFF_X1 port map( D => n3211, CK => CLK, Q => n_3558, QN 
                           => n9314);
   clk_r_REG1102_S1 : DFF_X1 port map( D => n3243, CK => CLK, Q => n_3559, QN 
                           => n9313);
   clk_r_REG776_S1 : DFF_X1 port map( D => n3275, CK => CLK, Q => n_3560, QN =>
                           n9312);
   clk_r_REG853_S1 : DFF_X1 port map( D => n3307, CK => CLK, Q => n_3561, QN =>
                           n9311);
   clk_r_REG1166_S1 : DFF_X1 port map( D => n3339, CK => CLK, Q => n_3562, QN 
                           => n9310);
   clk_r_REG1246_S1 : DFF_X1 port map( D => n3371, CK => CLK, Q => n_3563, QN 
                           => n9309);
   clk_r_REG693_S1 : DFF_X1 port map( D => n3403, CK => CLK, Q => n_3564, QN =>
                           n9308);
   clk_r_REG952_S1 : DFF_X1 port map( D => n3435, CK => CLK, Q => n_3565, QN =>
                           n9307);
   clk_r_REG1333_S1 : DFF_X1 port map( D => n3467, CK => CLK, Q => n_3566, QN 
                           => n9306);
   clk_r_REG1509_S1 : DFF_X1 port map( D => n3499, CK => CLK, Q => n_3567, QN 
                           => n9305);
   clk_r_REG3060_S1 : DFF_X1 port map( D => n3531, CK => CLK, Q => n_3568, QN 
                           => n9304);
   clk_r_REG3132_S1 : DFF_X1 port map( D => n3563, CK => CLK, Q => n_3569, QN 
                           => n9303);
   clk_r_REG2121_S1 : DFF_X1 port map( D => n2580, CK => CLK, Q => n_3570, QN 
                           => n9302);
   clk_r_REG2196_S1 : DFF_X1 port map( D => n2604, CK => CLK, Q => n_3571, QN 
                           => n9301);
   clk_r_REG2272_S1 : DFF_X1 port map( D => n2636, CK => CLK, Q => n_3572, QN 
                           => n9300);
   clk_r_REG2348_S1 : DFF_X1 port map( D => n2668, CK => CLK, Q => n_3573, QN 
                           => n9299);
   clk_r_REG2429_S1 : DFF_X1 port map( D => n2700, CK => CLK, Q => n_3574, QN 
                           => n9298);
   clk_r_REG2507_S1 : DFF_X1 port map( D => n2732, CK => CLK, Q => n_3575, QN 
                           => n9297);
   clk_r_REG2587_S1 : DFF_X1 port map( D => n2764, CK => CLK, Q => n_3576, QN 
                           => n9296);
   clk_r_REG2663_S1 : DFF_X1 port map( D => n2796, CK => CLK, Q => n_3577, QN 
                           => n9295);
   clk_r_REG1819_S1 : DFF_X1 port map( D => n2828, CK => CLK, Q => n_3578, QN 
                           => n9294);
   clk_r_REG1893_S1 : DFF_X1 port map( D => n2860, CK => CLK, Q => n_3579, QN 
                           => n9293);
   clk_r_REG1968_S1 : DFF_X1 port map( D => n2892, CK => CLK, Q => n_3580, QN 
                           => n9292);
   clk_r_REG2742_S1 : DFF_X1 port map( D => n2924, CK => CLK, Q => n_3581, QN 
                           => n9291);
   clk_r_REG2817_S1 : DFF_X1 port map( D => n2956, CK => CLK, Q => n_3582, QN 
                           => n9290);
   clk_r_REG2889_S1 : DFF_X1 port map( D => n2988, CK => CLK, Q => n_3583, QN 
                           => n9289);
   clk_r_REG2039_S1 : DFF_X1 port map( D => n3020, CK => CLK, Q => n_3584, QN 
                           => n9288);
   clk_r_REG2966_S1 : DFF_X1 port map( D => n3052, CK => CLK, Q => n_3585, QN 
                           => n9287);
   clk_r_REG1585_S1 : DFF_X1 port map( D => n3084, CK => CLK, Q => n_3586, QN 
                           => n9286);
   clk_r_REG1662_S1 : DFF_X1 port map( D => n3116, CK => CLK, Q => n_3587, QN 
                           => n9285);
   clk_r_REG1409_S1 : DFF_X1 port map( D => n3148, CK => CLK, Q => n_3588, QN 
                           => n9284);
   clk_r_REG1746_S1 : DFF_X1 port map( D => n3180, CK => CLK, Q => n_3589, QN 
                           => n9283);
   clk_r_REG1025_S1 : DFF_X1 port map( D => n3212, CK => CLK, Q => n_3590, QN 
                           => n9282);
   clk_r_REG1100_S1 : DFF_X1 port map( D => n3244, CK => CLK, Q => n_3591, QN 
                           => n9281);
   clk_r_REG774_S1 : DFF_X1 port map( D => n3276, CK => CLK, Q => n_3592, QN =>
                           n9280);
   clk_r_REG851_S1 : DFF_X1 port map( D => n3308, CK => CLK, Q => n_3593, QN =>
                           n9279);
   clk_r_REG1164_S1 : DFF_X1 port map( D => n3340, CK => CLK, Q => n_3594, QN 
                           => n9278);
   clk_r_REG1244_S1 : DFF_X1 port map( D => n3372, CK => CLK, Q => n_3595, QN 
                           => n9277);
   clk_r_REG691_S1 : DFF_X1 port map( D => n3404, CK => CLK, Q => n_3596, QN =>
                           n9276);
   clk_r_REG950_S1 : DFF_X1 port map( D => n3436, CK => CLK, Q => n_3597, QN =>
                           n9275);
   clk_r_REG1331_S1 : DFF_X1 port map( D => n3468, CK => CLK, Q => n_3598, QN 
                           => n9274);
   clk_r_REG1507_S1 : DFF_X1 port map( D => n3500, CK => CLK, Q => n_3599, QN 
                           => n9273);
   clk_r_REG3058_S1 : DFF_X1 port map( D => n3532, CK => CLK, Q => n_3600, QN 
                           => n9272);
   clk_r_REG3130_S1 : DFF_X1 port map( D => n3564, CK => CLK, Q => n_3601, QN 
                           => n9271);
   clk_r_REG2119_S1 : DFF_X1 port map( D => n2556, CK => CLK, Q => n_3602, QN 
                           => n9270);
   clk_r_REG2194_S1 : DFF_X1 port map( D => n2605, CK => CLK, Q => n_3603, QN 
                           => n9269);
   clk_r_REG2270_S1 : DFF_X1 port map( D => n2637, CK => CLK, Q => n_3604, QN 
                           => n9268);
   clk_r_REG2346_S1 : DFF_X1 port map( D => n2669, CK => CLK, Q => n_3605, QN 
                           => n9267);
   clk_r_REG2427_S1 : DFF_X1 port map( D => n2701, CK => CLK, Q => n_3606, QN 
                           => n9266);
   clk_r_REG2505_S1 : DFF_X1 port map( D => n2733, CK => CLK, Q => n_3607, QN 
                           => n9265);
   clk_r_REG2585_S1 : DFF_X1 port map( D => n2765, CK => CLK, Q => n_3608, QN 
                           => n9264);
   clk_r_REG2661_S1 : DFF_X1 port map( D => n2797, CK => CLK, Q => n_3609, QN 
                           => n9263);
   clk_r_REG1817_S1 : DFF_X1 port map( D => n2829, CK => CLK, Q => n_3610, QN 
                           => n9262);
   clk_r_REG1891_S1 : DFF_X1 port map( D => n2861, CK => CLK, Q => n_3611, QN 
                           => n9261);
   clk_r_REG1966_S1 : DFF_X1 port map( D => n2893, CK => CLK, Q => n_3612, QN 
                           => n9260);
   clk_r_REG2740_S1 : DFF_X1 port map( D => n2925, CK => CLK, Q => n_3613, QN 
                           => n9259);
   clk_r_REG2815_S1 : DFF_X1 port map( D => n2957, CK => CLK, Q => n_3614, QN 
                           => n9258);
   clk_r_REG2887_S1 : DFF_X1 port map( D => n2989, CK => CLK, Q => n_3615, QN 
                           => n9257);
   clk_r_REG2037_S1 : DFF_X1 port map( D => n3021, CK => CLK, Q => n_3616, QN 
                           => n9256);
   clk_r_REG2964_S1 : DFF_X1 port map( D => n3053, CK => CLK, Q => n_3617, QN 
                           => n9255);
   clk_r_REG1583_S1 : DFF_X1 port map( D => n3085, CK => CLK, Q => n_3618, QN 
                           => n9254);
   clk_r_REG1660_S1 : DFF_X1 port map( D => n3117, CK => CLK, Q => n_3619, QN 
                           => n9253);
   clk_r_REG1407_S1 : DFF_X1 port map( D => n3149, CK => CLK, Q => n_3620, QN 
                           => n9252);
   clk_r_REG1744_S1 : DFF_X1 port map( D => n3181, CK => CLK, Q => n_3621, QN 
                           => n9251);
   clk_r_REG1023_S1 : DFF_X1 port map( D => n3213, CK => CLK, Q => n_3622, QN 
                           => n9250);
   clk_r_REG1098_S1 : DFF_X1 port map( D => n3245, CK => CLK, Q => n_3623, QN 
                           => n9249);
   clk_r_REG772_S1 : DFF_X1 port map( D => n3277, CK => CLK, Q => n_3624, QN =>
                           n9248);
   clk_r_REG849_S1 : DFF_X1 port map( D => n3309, CK => CLK, Q => n_3625, QN =>
                           n9247);
   clk_r_REG1162_S1 : DFF_X1 port map( D => n3341, CK => CLK, Q => n_3626, QN 
                           => n9246);
   clk_r_REG1242_S1 : DFF_X1 port map( D => n3373, CK => CLK, Q => n_3627, QN 
                           => n9245);
   clk_r_REG689_S1 : DFF_X1 port map( D => n3405, CK => CLK, Q => n_3628, QN =>
                           n9244);
   clk_r_REG948_S1 : DFF_X1 port map( D => n3437, CK => CLK, Q => n_3629, QN =>
                           n9243);
   clk_r_REG1329_S1 : DFF_X1 port map( D => n3469, CK => CLK, Q => n_3630, QN 
                           => n9242);
   clk_r_REG1505_S1 : DFF_X1 port map( D => n3501, CK => CLK, Q => n_3631, QN 
                           => n9241);
   clk_r_REG3056_S1 : DFF_X1 port map( D => n3533, CK => CLK, Q => n_3632, QN 
                           => n9240);
   clk_r_REG3128_S1 : DFF_X1 port map( D => n3565, CK => CLK, Q => n_3633, QN 
                           => n9239);
   clk_r_REG2117_S1 : DFF_X1 port map( D => n2555, CK => CLK, Q => n_3634, QN 
                           => n9238);
   clk_r_REG2192_S1 : DFF_X1 port map( D => n2606, CK => CLK, Q => n_3635, QN 
                           => n9237);
   clk_r_REG2268_S1 : DFF_X1 port map( D => n2638, CK => CLK, Q => n_3636, QN 
                           => n9236);
   clk_r_REG2344_S1 : DFF_X1 port map( D => n2670, CK => CLK, Q => n_3637, QN 
                           => n9235);
   clk_r_REG2425_S1 : DFF_X1 port map( D => n2702, CK => CLK, Q => n_3638, QN 
                           => n9234);
   clk_r_REG2503_S1 : DFF_X1 port map( D => n2734, CK => CLK, Q => n_3639, QN 
                           => n9233);
   clk_r_REG2583_S1 : DFF_X1 port map( D => n2766, CK => CLK, Q => n_3640, QN 
                           => n9232);
   clk_r_REG2659_S1 : DFF_X1 port map( D => n2798, CK => CLK, Q => n_3641, QN 
                           => n9231);
   clk_r_REG1815_S1 : DFF_X1 port map( D => n2830, CK => CLK, Q => n_3642, QN 
                           => n9230);
   clk_r_REG1889_S1 : DFF_X1 port map( D => n2862, CK => CLK, Q => n_3643, QN 
                           => n9229);
   clk_r_REG1964_S1 : DFF_X1 port map( D => n2894, CK => CLK, Q => n_3644, QN 
                           => n9228);
   clk_r_REG2738_S1 : DFF_X1 port map( D => n2926, CK => CLK, Q => n_3645, QN 
                           => n9227);
   clk_r_REG2813_S1 : DFF_X1 port map( D => n2958, CK => CLK, Q => n_3646, QN 
                           => n9226);
   clk_r_REG2885_S1 : DFF_X1 port map( D => n2990, CK => CLK, Q => n_3647, QN 
                           => n9225);
   clk_r_REG2035_S1 : DFF_X1 port map( D => n3022, CK => CLK, Q => n_3648, QN 
                           => n9224);
   clk_r_REG2962_S1 : DFF_X1 port map( D => n3054, CK => CLK, Q => n_3649, QN 
                           => n9223);
   clk_r_REG1581_S1 : DFF_X1 port map( D => n3086, CK => CLK, Q => n_3650, QN 
                           => n9222);
   clk_r_REG1658_S1 : DFF_X1 port map( D => n3118, CK => CLK, Q => n_3651, QN 
                           => n9221);
   clk_r_REG1405_S1 : DFF_X1 port map( D => n3150, CK => CLK, Q => n_3652, QN 
                           => n9220);
   clk_r_REG1742_S1 : DFF_X1 port map( D => n3182, CK => CLK, Q => n_3653, QN 
                           => n9219);
   clk_r_REG1021_S1 : DFF_X1 port map( D => n3214, CK => CLK, Q => n_3654, QN 
                           => n9218);
   clk_r_REG1096_S1 : DFF_X1 port map( D => n3246, CK => CLK, Q => n_3655, QN 
                           => n9217);
   clk_r_REG770_S1 : DFF_X1 port map( D => n3278, CK => CLK, Q => n_3656, QN =>
                           n9216);
   clk_r_REG847_S1 : DFF_X1 port map( D => n3310, CK => CLK, Q => n_3657, QN =>
                           n9215);
   clk_r_REG1160_S1 : DFF_X1 port map( D => n3342, CK => CLK, Q => n_3658, QN 
                           => n9214);
   clk_r_REG1240_S1 : DFF_X1 port map( D => n3374, CK => CLK, Q => n_3659, QN 
                           => n9213);
   clk_r_REG687_S1 : DFF_X1 port map( D => n3406, CK => CLK, Q => n_3660, QN =>
                           n9212);
   clk_r_REG946_S1 : DFF_X1 port map( D => n3438, CK => CLK, Q => n_3661, QN =>
                           n9211);
   clk_r_REG1327_S1 : DFF_X1 port map( D => n3470, CK => CLK, Q => n_3662, QN 
                           => n9210);
   clk_r_REG1503_S1 : DFF_X1 port map( D => n3502, CK => CLK, Q => n_3663, QN 
                           => n9209);
   clk_r_REG3054_S1 : DFF_X1 port map( D => n3534, CK => CLK, Q => n_3664, QN 
                           => n9208);
   clk_r_REG3126_S1 : DFF_X1 port map( D => n3566, CK => CLK, Q => n_3665, QN 
                           => n9207);
   clk_r_REG2115_S1 : DFF_X1 port map( D => n2554, CK => CLK, Q => n_3666, QN 
                           => n9206);
   clk_r_REG2190_S1 : DFF_X1 port map( D => n2607, CK => CLK, Q => n_3667, QN 
                           => n9205);
   clk_r_REG2266_S1 : DFF_X1 port map( D => n2639, CK => CLK, Q => n_3668, QN 
                           => n9204);
   clk_r_REG2342_S1 : DFF_X1 port map( D => n2671, CK => CLK, Q => n_3669, QN 
                           => n9203);
   clk_r_REG2423_S1 : DFF_X1 port map( D => n2703, CK => CLK, Q => n_3670, QN 
                           => n9202);
   clk_r_REG2501_S1 : DFF_X1 port map( D => n2735, CK => CLK, Q => n_3671, QN 
                           => n9201);
   clk_r_REG2581_S1 : DFF_X1 port map( D => n2767, CK => CLK, Q => n_3672, QN 
                           => n9200);
   clk_r_REG2657_S1 : DFF_X1 port map( D => n2799, CK => CLK, Q => n_3673, QN 
                           => n9199);
   clk_r_REG1813_S1 : DFF_X1 port map( D => n2831, CK => CLK, Q => n_3674, QN 
                           => n9198);
   clk_r_REG1887_S1 : DFF_X1 port map( D => n2863, CK => CLK, Q => n_3675, QN 
                           => n9197);
   clk_r_REG1962_S1 : DFF_X1 port map( D => n2895, CK => CLK, Q => n_3676, QN 
                           => n9196);
   clk_r_REG2736_S1 : DFF_X1 port map( D => n2927, CK => CLK, Q => n_3677, QN 
                           => n9195);
   clk_r_REG2811_S1 : DFF_X1 port map( D => n2959, CK => CLK, Q => n_3678, QN 
                           => n9194);
   clk_r_REG2883_S1 : DFF_X1 port map( D => n2991, CK => CLK, Q => n_3679, QN 
                           => n9193);
   clk_r_REG2033_S1 : DFF_X1 port map( D => n3023, CK => CLK, Q => n_3680, QN 
                           => n9192);
   clk_r_REG2960_S1 : DFF_X1 port map( D => n3055, CK => CLK, Q => n_3681, QN 
                           => n9191);
   clk_r_REG1579_S1 : DFF_X1 port map( D => n3087, CK => CLK, Q => n_3682, QN 
                           => n9190);
   clk_r_REG1656_S1 : DFF_X1 port map( D => n3119, CK => CLK, Q => n_3683, QN 
                           => n9189);
   clk_r_REG1403_S1 : DFF_X1 port map( D => n3151, CK => CLK, Q => n_3684, QN 
                           => n9188);
   clk_r_REG1740_S1 : DFF_X1 port map( D => n3183, CK => CLK, Q => n_3685, QN 
                           => n9187);
   clk_r_REG1019_S1 : DFF_X1 port map( D => n3215, CK => CLK, Q => n_3686, QN 
                           => n9186);
   clk_r_REG1094_S1 : DFF_X1 port map( D => n3247, CK => CLK, Q => n_3687, QN 
                           => n9185);
   clk_r_REG768_S1 : DFF_X1 port map( D => n3279, CK => CLK, Q => n_3688, QN =>
                           n9184);
   clk_r_REG845_S1 : DFF_X1 port map( D => n3311, CK => CLK, Q => n_3689, QN =>
                           n9183);
   clk_r_REG1158_S1 : DFF_X1 port map( D => n3343, CK => CLK, Q => n_3690, QN 
                           => n9182);
   clk_r_REG1238_S1 : DFF_X1 port map( D => n3375, CK => CLK, Q => n_3691, QN 
                           => n9181);
   clk_r_REG685_S1 : DFF_X1 port map( D => n3407, CK => CLK, Q => n_3692, QN =>
                           n9180);
   clk_r_REG944_S1 : DFF_X1 port map( D => n3439, CK => CLK, Q => n_3693, QN =>
                           n9179);
   clk_r_REG1325_S1 : DFF_X1 port map( D => n3471, CK => CLK, Q => n_3694, QN 
                           => n9178);
   clk_r_REG1501_S1 : DFF_X1 port map( D => n3503, CK => CLK, Q => n_3695, QN 
                           => n9177);
   clk_r_REG3052_S1 : DFF_X1 port map( D => n3535, CK => CLK, Q => n_3696, QN 
                           => n9176);
   clk_r_REG3124_S1 : DFF_X1 port map( D => n3567, CK => CLK, Q => n_3697, QN 
                           => n9175);
   clk_r_REG2113_S1 : DFF_X1 port map( D => n2553, CK => CLK, Q => n_3698, QN 
                           => n9174);
   clk_r_REG2188_S1 : DFF_X1 port map( D => n2608, CK => CLK, Q => n_3699, QN 
                           => n9173);
   clk_r_REG2264_S1 : DFF_X1 port map( D => n2640, CK => CLK, Q => n_3700, QN 
                           => n9172);
   clk_r_REG2340_S1 : DFF_X1 port map( D => n2672, CK => CLK, Q => n_3701, QN 
                           => n9171);
   clk_r_REG2421_S1 : DFF_X1 port map( D => n2704, CK => CLK, Q => n_3702, QN 
                           => n9170);
   clk_r_REG2499_S1 : DFF_X1 port map( D => n2736, CK => CLK, Q => n_3703, QN 
                           => n9169);
   clk_r_REG2579_S1 : DFF_X1 port map( D => n2768, CK => CLK, Q => n_3704, QN 
                           => n9168);
   clk_r_REG2655_S1 : DFF_X1 port map( D => n2800, CK => CLK, Q => n_3705, QN 
                           => n9167);
   clk_r_REG1811_S1 : DFF_X1 port map( D => n2832, CK => CLK, Q => n_3706, QN 
                           => n9166);
   clk_r_REG1885_S1 : DFF_X1 port map( D => n2864, CK => CLK, Q => n_3707, QN 
                           => n9165);
   clk_r_REG1960_S1 : DFF_X1 port map( D => n2896, CK => CLK, Q => n_3708, QN 
                           => n9164);
   clk_r_REG2734_S1 : DFF_X1 port map( D => n2928, CK => CLK, Q => n_3709, QN 
                           => n9163);
   clk_r_REG2809_S1 : DFF_X1 port map( D => n2960, CK => CLK, Q => n_3710, QN 
                           => n9162);
   clk_r_REG2881_S1 : DFF_X1 port map( D => n2992, CK => CLK, Q => n_3711, QN 
                           => n9161);
   clk_r_REG2031_S1 : DFF_X1 port map( D => n3024, CK => CLK, Q => n_3712, QN 
                           => n9160);
   clk_r_REG2958_S1 : DFF_X1 port map( D => n3056, CK => CLK, Q => n_3713, QN 
                           => n9159);
   clk_r_REG1577_S1 : DFF_X1 port map( D => n3088, CK => CLK, Q => n_3714, QN 
                           => n9158);
   clk_r_REG1654_S1 : DFF_X1 port map( D => n3120, CK => CLK, Q => n_3715, QN 
                           => n9157);
   clk_r_REG1401_S1 : DFF_X1 port map( D => n3152, CK => CLK, Q => n_3716, QN 
                           => n9156);
   clk_r_REG1738_S1 : DFF_X1 port map( D => n3184, CK => CLK, Q => n_3717, QN 
                           => n9155);
   clk_r_REG1017_S1 : DFF_X1 port map( D => n3216, CK => CLK, Q => n_3718, QN 
                           => n9154);
   clk_r_REG1092_S1 : DFF_X1 port map( D => n3248, CK => CLK, Q => n_3719, QN 
                           => n9153);
   clk_r_REG766_S1 : DFF_X1 port map( D => n3280, CK => CLK, Q => n_3720, QN =>
                           n9152);
   clk_r_REG843_S1 : DFF_X1 port map( D => n3312, CK => CLK, Q => n_3721, QN =>
                           n9151);
   clk_r_REG1156_S1 : DFF_X1 port map( D => n3344, CK => CLK, Q => n_3722, QN 
                           => n9150);
   clk_r_REG1236_S1 : DFF_X1 port map( D => n3376, CK => CLK, Q => n_3723, QN 
                           => n9149);
   clk_r_REG683_S1 : DFF_X1 port map( D => n3408, CK => CLK, Q => n_3724, QN =>
                           n9148);
   clk_r_REG942_S1 : DFF_X1 port map( D => n3440, CK => CLK, Q => n_3725, QN =>
                           n9147);
   clk_r_REG1323_S1 : DFF_X1 port map( D => n3472, CK => CLK, Q => n_3726, QN 
                           => n9146);
   clk_r_REG1499_S1 : DFF_X1 port map( D => n3504, CK => CLK, Q => n_3727, QN 
                           => n9145);
   clk_r_REG3050_S1 : DFF_X1 port map( D => n3536, CK => CLK, Q => n_3728, QN 
                           => n9144);
   clk_r_REG3122_S1 : DFF_X1 port map( D => n3568, CK => CLK, Q => n_3729, QN 
                           => n9143);
   clk_r_REG2111_S1 : DFF_X1 port map( D => n2552, CK => CLK, Q => n_3730, QN 
                           => n9142);
   clk_r_REG2186_S1 : DFF_X1 port map( D => n2609, CK => CLK, Q => n_3731, QN 
                           => n9141);
   clk_r_REG2262_S1 : DFF_X1 port map( D => n2641, CK => CLK, Q => n_3732, QN 
                           => n9140);
   clk_r_REG2338_S1 : DFF_X1 port map( D => n2673, CK => CLK, Q => n_3733, QN 
                           => n9139);
   clk_r_REG2419_S1 : DFF_X1 port map( D => n2705, CK => CLK, Q => n_3734, QN 
                           => n9138);
   clk_r_REG2497_S1 : DFF_X1 port map( D => n2737, CK => CLK, Q => n_3735, QN 
                           => n9137);
   clk_r_REG2577_S1 : DFF_X1 port map( D => n2769, CK => CLK, Q => n_3736, QN 
                           => n9136);
   clk_r_REG2653_S1 : DFF_X1 port map( D => n2801, CK => CLK, Q => n_3737, QN 
                           => n9135);
   clk_r_REG1809_S1 : DFF_X1 port map( D => n2833, CK => CLK, Q => n_3738, QN 
                           => n9134);
   clk_r_REG1883_S1 : DFF_X1 port map( D => n2865, CK => CLK, Q => n_3739, QN 
                           => n9133);
   clk_r_REG1958_S1 : DFF_X1 port map( D => n2897, CK => CLK, Q => n_3740, QN 
                           => n9132);
   clk_r_REG2732_S1 : DFF_X1 port map( D => n2929, CK => CLK, Q => n_3741, QN 
                           => n9131);
   clk_r_REG2807_S1 : DFF_X1 port map( D => n2961, CK => CLK, Q => n_3742, QN 
                           => n9130);
   clk_r_REG2879_S1 : DFF_X1 port map( D => n2993, CK => CLK, Q => n_3743, QN 
                           => n9129);
   clk_r_REG2029_S1 : DFF_X1 port map( D => n3025, CK => CLK, Q => n_3744, QN 
                           => n9128);
   clk_r_REG2956_S1 : DFF_X1 port map( D => n3057, CK => CLK, Q => n_3745, QN 
                           => n9127);
   clk_r_REG1575_S1 : DFF_X1 port map( D => n3089, CK => CLK, Q => n_3746, QN 
                           => n9126);
   clk_r_REG1652_S1 : DFF_X1 port map( D => n3121, CK => CLK, Q => n_3747, QN 
                           => n9125);
   clk_r_REG1399_S1 : DFF_X1 port map( D => n3153, CK => CLK, Q => n_3748, QN 
                           => n9124);
   clk_r_REG1736_S1 : DFF_X1 port map( D => n3185, CK => CLK, Q => n_3749, QN 
                           => n9123);
   clk_r_REG1015_S1 : DFF_X1 port map( D => n3217, CK => CLK, Q => n_3750, QN 
                           => n9122);
   clk_r_REG1090_S1 : DFF_X1 port map( D => n3249, CK => CLK, Q => n_3751, QN 
                           => n9121);
   clk_r_REG764_S1 : DFF_X1 port map( D => n3281, CK => CLK, Q => n_3752, QN =>
                           n9120);
   clk_r_REG841_S1 : DFF_X1 port map( D => n3313, CK => CLK, Q => n_3753, QN =>
                           n9119);
   clk_r_REG1154_S1 : DFF_X1 port map( D => n3345, CK => CLK, Q => n_3754, QN 
                           => n9118);
   clk_r_REG1234_S1 : DFF_X1 port map( D => n3377, CK => CLK, Q => n_3755, QN 
                           => n9117);
   clk_r_REG681_S1 : DFF_X1 port map( D => n3409, CK => CLK, Q => n_3756, QN =>
                           n9116);
   clk_r_REG940_S1 : DFF_X1 port map( D => n3441, CK => CLK, Q => n_3757, QN =>
                           n9115);
   clk_r_REG1321_S1 : DFF_X1 port map( D => n3473, CK => CLK, Q => n_3758, QN 
                           => n9114);
   clk_r_REG1497_S1 : DFF_X1 port map( D => n3505, CK => CLK, Q => n_3759, QN 
                           => n9113);
   clk_r_REG3048_S1 : DFF_X1 port map( D => n3537, CK => CLK, Q => n_3760, QN 
                           => n9112);
   clk_r_REG3120_S1 : DFF_X1 port map( D => n3569, CK => CLK, Q => n_3761, QN 
                           => n9111);
   clk_r_REG2109_S1 : DFF_X1 port map( D => n2551, CK => CLK, Q => n_3762, QN 
                           => n9110);
   clk_r_REG2184_S1 : DFF_X1 port map( D => n2610, CK => CLK, Q => n_3763, QN 
                           => n9109);
   clk_r_REG2260_S1 : DFF_X1 port map( D => n2642, CK => CLK, Q => n_3764, QN 
                           => n9108);
   clk_r_REG2336_S1 : DFF_X1 port map( D => n2674, CK => CLK, Q => n_3765, QN 
                           => n9107);
   clk_r_REG2417_S1 : DFF_X1 port map( D => n2706, CK => CLK, Q => n_3766, QN 
                           => n9106);
   clk_r_REG2495_S1 : DFF_X1 port map( D => n2738, CK => CLK, Q => n_3767, QN 
                           => n9105);
   clk_r_REG2575_S1 : DFF_X1 port map( D => n2770, CK => CLK, Q => n_3768, QN 
                           => n9104);
   clk_r_REG2651_S1 : DFF_X1 port map( D => n2802, CK => CLK, Q => n_3769, QN 
                           => n9103);
   clk_r_REG1807_S1 : DFF_X1 port map( D => n2834, CK => CLK, Q => n_3770, QN 
                           => n9102);
   clk_r_REG1881_S1 : DFF_X1 port map( D => n2866, CK => CLK, Q => n_3771, QN 
                           => n9101);
   clk_r_REG1956_S1 : DFF_X1 port map( D => n2898, CK => CLK, Q => n_3772, QN 
                           => n9100);
   clk_r_REG2730_S1 : DFF_X1 port map( D => n2930, CK => CLK, Q => n_3773, QN 
                           => n9099);
   clk_r_REG2805_S1 : DFF_X1 port map( D => n2962, CK => CLK, Q => n_3774, QN 
                           => n9098);
   clk_r_REG2877_S1 : DFF_X1 port map( D => n2994, CK => CLK, Q => n_3775, QN 
                           => n9097);
   clk_r_REG2027_S1 : DFF_X1 port map( D => n3026, CK => CLK, Q => n_3776, QN 
                           => n9096);
   clk_r_REG2954_S1 : DFF_X1 port map( D => n3058, CK => CLK, Q => n_3777, QN 
                           => n9095);
   clk_r_REG1573_S1 : DFF_X1 port map( D => n3090, CK => CLK, Q => n_3778, QN 
                           => n9094);
   clk_r_REG1650_S1 : DFF_X1 port map( D => n3122, CK => CLK, Q => n_3779, QN 
                           => n9093);
   clk_r_REG1397_S1 : DFF_X1 port map( D => n3154, CK => CLK, Q => n_3780, QN 
                           => n9092);
   clk_r_REG1734_S1 : DFF_X1 port map( D => n3186, CK => CLK, Q => n_3781, QN 
                           => n9091);
   clk_r_REG1013_S1 : DFF_X1 port map( D => n3218, CK => CLK, Q => n_3782, QN 
                           => n9090);
   clk_r_REG1088_S1 : DFF_X1 port map( D => n3250, CK => CLK, Q => n_3783, QN 
                           => n9089);
   clk_r_REG762_S1 : DFF_X1 port map( D => n3282, CK => CLK, Q => n_3784, QN =>
                           n9088);
   clk_r_REG839_S1 : DFF_X1 port map( D => n3314, CK => CLK, Q => n_3785, QN =>
                           n9087);
   clk_r_REG1152_S1 : DFF_X1 port map( D => n3346, CK => CLK, Q => n_3786, QN 
                           => n9086);
   clk_r_REG1232_S1 : DFF_X1 port map( D => n3378, CK => CLK, Q => n_3787, QN 
                           => n9085);
   clk_r_REG679_S1 : DFF_X1 port map( D => n3410, CK => CLK, Q => n_3788, QN =>
                           n9084);
   clk_r_REG938_S1 : DFF_X1 port map( D => n3442, CK => CLK, Q => n_3789, QN =>
                           n9083);
   clk_r_REG1319_S1 : DFF_X1 port map( D => n3474, CK => CLK, Q => n_3790, QN 
                           => n9082);
   clk_r_REG1495_S1 : DFF_X1 port map( D => n3506, CK => CLK, Q => n_3791, QN 
                           => n9081);
   clk_r_REG3046_S1 : DFF_X1 port map( D => n3538, CK => CLK, Q => n_3792, QN 
                           => n9080);
   clk_r_REG3118_S1 : DFF_X1 port map( D => n3570, CK => CLK, Q => n_3793, QN 
                           => n9079);
   clk_r_REG2107_S1 : DFF_X1 port map( D => n2550, CK => CLK, Q => n_3794, QN 
                           => n9078);
   clk_r_REG2182_S1 : DFF_X1 port map( D => n2611, CK => CLK, Q => n_3795, QN 
                           => n9077);
   clk_r_REG2258_S1 : DFF_X1 port map( D => n2643, CK => CLK, Q => n_3796, QN 
                           => n9076);
   clk_r_REG2334_S1 : DFF_X1 port map( D => n2675, CK => CLK, Q => n_3797, QN 
                           => n9075);
   clk_r_REG2415_S1 : DFF_X1 port map( D => n2707, CK => CLK, Q => n_3798, QN 
                           => n9074);
   clk_r_REG2493_S1 : DFF_X1 port map( D => n2739, CK => CLK, Q => n_3799, QN 
                           => n9073);
   clk_r_REG2573_S1 : DFF_X1 port map( D => n2771, CK => CLK, Q => n_3800, QN 
                           => n9072);
   clk_r_REG2649_S1 : DFF_X1 port map( D => n2803, CK => CLK, Q => n_3801, QN 
                           => n9071);
   clk_r_REG1805_S1 : DFF_X1 port map( D => n2835, CK => CLK, Q => n_3802, QN 
                           => n9070);
   clk_r_REG1879_S1 : DFF_X1 port map( D => n2867, CK => CLK, Q => n_3803, QN 
                           => n9069);
   clk_r_REG1954_S1 : DFF_X1 port map( D => n2899, CK => CLK, Q => n_3804, QN 
                           => n9068);
   clk_r_REG2728_S1 : DFF_X1 port map( D => n2931, CK => CLK, Q => n_3805, QN 
                           => n9067);
   clk_r_REG2803_S1 : DFF_X1 port map( D => n2963, CK => CLK, Q => n_3806, QN 
                           => n9066);
   clk_r_REG2875_S1 : DFF_X1 port map( D => n2995, CK => CLK, Q => n_3807, QN 
                           => n9065);
   clk_r_REG2025_S1 : DFF_X1 port map( D => n3027, CK => CLK, Q => n_3808, QN 
                           => n9064);
   clk_r_REG2952_S1 : DFF_X1 port map( D => n3059, CK => CLK, Q => n_3809, QN 
                           => n9063);
   clk_r_REG1571_S1 : DFF_X1 port map( D => n3091, CK => CLK, Q => n_3810, QN 
                           => n9062);
   clk_r_REG1648_S1 : DFF_X1 port map( D => n3123, CK => CLK, Q => n_3811, QN 
                           => n9061);
   clk_r_REG1395_S1 : DFF_X1 port map( D => n3155, CK => CLK, Q => n_3812, QN 
                           => n9060);
   clk_r_REG1732_S1 : DFF_X1 port map( D => n3187, CK => CLK, Q => n_3813, QN 
                           => n9059);
   clk_r_REG1011_S1 : DFF_X1 port map( D => n3219, CK => CLK, Q => n_3814, QN 
                           => n9058);
   clk_r_REG1086_S1 : DFF_X1 port map( D => n3251, CK => CLK, Q => n_3815, QN 
                           => n9057);
   clk_r_REG760_S1 : DFF_X1 port map( D => n3283, CK => CLK, Q => n_3816, QN =>
                           n9056);
   clk_r_REG837_S1 : DFF_X1 port map( D => n3315, CK => CLK, Q => n_3817, QN =>
                           n9055);
   clk_r_REG1150_S1 : DFF_X1 port map( D => n3347, CK => CLK, Q => n_3818, QN 
                           => n9054);
   clk_r_REG1230_S1 : DFF_X1 port map( D => n3379, CK => CLK, Q => n_3819, QN 
                           => n9053);
   clk_r_REG677_S1 : DFF_X1 port map( D => n3411, CK => CLK, Q => n_3820, QN =>
                           n9052);
   clk_r_REG936_S1 : DFF_X1 port map( D => n3443, CK => CLK, Q => n_3821, QN =>
                           n9051);
   clk_r_REG1317_S1 : DFF_X1 port map( D => n3475, CK => CLK, Q => n_3822, QN 
                           => n9050);
   clk_r_REG1493_S1 : DFF_X1 port map( D => n3507, CK => CLK, Q => n_3823, QN 
                           => n9049);
   clk_r_REG3044_S1 : DFF_X1 port map( D => n3539, CK => CLK, Q => n_3824, QN 
                           => n9048);
   clk_r_REG3116_S1 : DFF_X1 port map( D => n3571, CK => CLK, Q => n_3825, QN 
                           => n9047);
   clk_r_REG121_S1 : DFF_X1 port map( D => n2549, CK => CLK, Q => n_3826, QN =>
                           n9046);
   clk_r_REG2171_S1 : DFF_X1 port map( D => n2612, CK => CLK, Q => n_3827, QN 
                           => n9045);
   clk_r_REG2248_S1 : DFF_X1 port map( D => n2644, CK => CLK, Q => n_3828, QN 
                           => n9044);
   clk_r_REG2322_S1 : DFF_X1 port map( D => n2676, CK => CLK, Q => n_3829, QN 
                           => n9043);
   clk_r_REG2402_S1 : DFF_X1 port map( D => n2708, CK => CLK, Q => n_3830, QN 
                           => n9042);
   clk_r_REG2479_S1 : DFF_X1 port map( D => n2740, CK => CLK, Q => n_3831, QN 
                           => n9041);
   clk_r_REG2560_S1 : DFF_X1 port map( D => n2772, CK => CLK, Q => n_3832, QN 
                           => n9040);
   clk_r_REG2637_S1 : DFF_X1 port map( D => n2804, CK => CLK, Q => n_3833, QN 
                           => n9039);
   clk_r_REG1797_S1 : DFF_X1 port map( D => n2836, CK => CLK, Q => n_3834, QN 
                           => n9038);
   clk_r_REG1869_S1 : DFF_X1 port map( D => n2868, CK => CLK, Q => n_3835, QN 
                           => n9037);
   clk_r_REG1946_S1 : DFF_X1 port map( D => n2900, CK => CLK, Q => n_3836, QN 
                           => n9036);
   clk_r_REG2718_S1 : DFF_X1 port map( D => n2932, CK => CLK, Q => n_3837, QN 
                           => n9035);
   clk_r_REG2794_S1 : DFF_X1 port map( D => n2964, CK => CLK, Q => n_3838, QN 
                           => n9034);
   clk_r_REG2867_S1 : DFF_X1 port map( D => n2996, CK => CLK, Q => n_3839, QN 
                           => n9033);
   clk_r_REG2018_S1 : DFF_X1 port map( D => n3028, CK => CLK, Q => n_3840, QN 
                           => n9032);
   clk_r_REG2944_S1 : DFF_X1 port map( D => n3060, CK => CLK, Q => n_3841, QN 
                           => n9031);
   clk_r_REG1559_S1 : DFF_X1 port map( D => n3092, CK => CLK, Q => n_3842, QN 
                           => n9030);
   clk_r_REG1635_S1 : DFF_X1 port map( D => n3124, CK => CLK, Q => n_3843, QN 
                           => n9029);
   clk_r_REG1381_S1 : DFF_X1 port map( D => n3156, CK => CLK, Q => n_3844, QN 
                           => n9028);
   clk_r_REG1721_S1 : DFF_X1 port map( D => n3188, CK => CLK, Q => n_3845, QN 
                           => n9027);
   clk_r_REG1000_S1 : DFF_X1 port map( D => n3220, CK => CLK, Q => n_3846, QN 
                           => n9026);
   clk_r_REG1075_S1 : DFF_X1 port map( D => n3252, CK => CLK, Q => n_3847, QN 
                           => n9025);
   clk_r_REG746_S1 : DFF_X1 port map( D => n3284, CK => CLK, Q => n_3848, QN =>
                           n9024);
   clk_r_REG824_S1 : DFF_X1 port map( D => n3316, CK => CLK, Q => n_3849, QN =>
                           n9023);
   clk_r_REG385_S1 : DFF_X1 port map( D => n3348, CK => CLK, Q => n_3850, QN =>
                           n9022);
   clk_r_REG1222_S1 : DFF_X1 port map( D => n3380, CK => CLK, Q => n_3851, QN 
                           => n9021);
   clk_r_REG521_S1 : DFF_X1 port map( D => n3412, CK => CLK, Q => n_3852, QN =>
                           n9020);
   clk_r_REG905_S1 : DFF_X1 port map( D => n3444, CK => CLK, Q => n_3853, QN =>
                           n9019);
   clk_r_REG358_S1 : DFF_X1 port map( D => n3476, CK => CLK, Q => n_3854, QN =>
                           n9018);
   clk_r_REG1486_S1 : DFF_X1 port map( D => n3508, CK => CLK, Q => n_3855, QN 
                           => n9017);
   clk_r_REG3038_S1 : DFF_X1 port map( D => n3540, CK => CLK, Q => n_3856, QN 
                           => n9016);
   clk_r_REG3113_S1 : DFF_X1 port map( D => n3572, CK => CLK, Q => n_3857, QN 
                           => n9015);
   clk_r_REG3354_S7 : DFFR_X1 port map( D => n3575, CK => CLK, RN => RESET_BAR,
                           Q => n11228, QN => n_3858);
   clk_r_REG3342_S7 : DFFR_X1 port map( D => n3582, CK => CLK, RN => RESET_BAR,
                           Q => n11225, QN => n_3859);
   clk_r_REG3380_S7 : DFFR_X1 port map( D => n3580, CK => CLK, RN => RESET_BAR,
                           Q => n11230, QN => n_3860);
   clk_r_REG3434_S7 : DFFS_X1 port map( D => n3589, CK => CLK, SN => RESET_BAR,
                           Q => n11227, QN => n_3861);
   clk_r_REG3367_S7 : DFFR_X1 port map( D => n3577, CK => CLK, RN => RESET_BAR,
                           Q => n11232, QN => n_3862);
   clk_r_REG3386_S7 : DFFS_X1 port map( D => n3579, CK => CLK, SN => RESET_BAR,
                           Q => n11231, QN => n_3863);
   clk_r_REG3348_S7 : DFFR_X1 port map( D => n3581, CK => CLK, RN => RESET_BAR,
                           Q => n11229, QN => n_3864);
   clk_r_REG3436_S7 : DFFR_X1 port map( D => n3588, CK => CLK, RN => RESET_BAR,
                           Q => n11226, QN => n_3865);
   clk_r_REG3202_S2 : DFFS_X1 port map( D => n4097, CK => CLK, SN => RESET_BAR,
                           Q => n11224, QN => n_3866);
   clk_r_REG3216_S2 : DFFS_X1 port map( D => n4063, CK => CLK, SN => RESET_BAR,
                           Q => n11223, QN => n_3867);
   clk_r_REG3236_S2 : DFFS_X1 port map( D => n4005, CK => CLK, SN => RESET_BAR,
                           Q => n11222, QN => n_3868);
   clk_r_REG3244_S2 : DFFS_X1 port map( D => n3991, CK => CLK, SN => RESET_BAR,
                           Q => n11220, QN => n_3869);
   clk_r_REG3242_S2 : DFFS_X1 port map( D => n3994, CK => CLK, SN => RESET_BAR,
                           Q => n11219, QN => n_3870);
   clk_r_REG3240_S2 : DFFS_X1 port map( D => n3997, CK => CLK, SN => RESET_BAR,
                           Q => n11218, QN => n_3871);
   clk_r_REG3238_S2 : DFFS_X1 port map( D => n4000, CK => CLK, SN => RESET_BAR,
                           Q => n11217, QN => n_3872);
   clk_r_REG3234_S2 : DFFS_X1 port map( D => n4009, CK => CLK, SN => RESET_BAR,
                           Q => n11216, QN => n_3873);
   clk_r_REG3232_S2 : DFFS_X1 port map( D => n4034, CK => CLK, SN => RESET_BAR,
                           Q => n11215, QN => n_3874);
   clk_r_REG3230_S2 : DFFS_X1 port map( D => n4039, CK => CLK, SN => RESET_BAR,
                           Q => n11214, QN => n_3875);
   clk_r_REG3228_S2 : DFFS_X1 port map( D => n4043, CK => CLK, SN => RESET_BAR,
                           Q => n11213, QN => n_3876);
   clk_r_REG3226_S2 : DFFS_X1 port map( D => n4046, CK => CLK, SN => RESET_BAR,
                           Q => n11212, QN => n_3877);
   clk_r_REG3224_S2 : DFFS_X1 port map( D => n4049, CK => CLK, SN => RESET_BAR,
                           Q => n11211, QN => n_3878);
   clk_r_REG3222_S2 : DFFS_X1 port map( D => n4052, CK => CLK, SN => RESET_BAR,
                           Q => n11210, QN => n_3879);
   clk_r_REG3220_S2 : DFFS_X1 port map( D => n4055, CK => CLK, SN => RESET_BAR,
                           Q => n11209, QN => n_3880);
   clk_r_REG3218_S2 : DFFS_X1 port map( D => n4059, CK => CLK, SN => RESET_BAR,
                           Q => n11208, QN => n_3881);
   clk_r_REG3214_S2 : DFFS_X1 port map( D => n4067, CK => CLK, SN => RESET_BAR,
                           Q => n11207, QN => n_3882);
   clk_r_REG3212_S2 : DFFS_X1 port map( D => n4071, CK => CLK, SN => RESET_BAR,
                           Q => n11206, QN => n_3883);
   clk_r_REG3210_S2 : DFFS_X1 port map( D => n4075, CK => CLK, SN => RESET_BAR,
                           Q => n11205, QN => n_3884);
   clk_r_REG3208_S2 : DFFS_X1 port map( D => n4079, CK => CLK, SN => RESET_BAR,
                           Q => n11204, QN => n_3885);
   clk_r_REG3206_S2 : DFFS_X1 port map( D => n4090, CK => CLK, SN => RESET_BAR,
                           Q => n11203, QN => n_3886);
   clk_r_REG3204_S2 : DFFS_X1 port map( D => n4094, CK => CLK, SN => RESET_BAR,
                           Q => n11202, QN => n_3887);
   clk_r_REG3200_S2 : DFFS_X1 port map( D => n4102, CK => CLK, SN => RESET_BAR,
                           Q => n11201, QN => n_3888);
   clk_r_REG3198_S2 : DFFS_X1 port map( D => n4110, CK => CLK, SN => RESET_BAR,
                           Q => n11200, QN => n_3889);
   clk_r_REG3196_S2 : DFFS_X1 port map( D => n4115, CK => CLK, SN => RESET_BAR,
                           Q => n11199, QN => n_3890);
   clk_r_REG3194_S2 : DFFS_X1 port map( D => n4120, CK => CLK, SN => RESET_BAR,
                           Q => n11198, QN => n_3891);
   clk_r_REG3192_S2 : DFFS_X1 port map( D => n4125, CK => CLK, SN => RESET_BAR,
                           Q => n11197, QN => n_3892);
   clk_r_REG3190_S2 : DFFS_X1 port map( D => n4130, CK => CLK, SN => RESET_BAR,
                           Q => n11196, QN => n_3893);
   clk_r_REG3188_S2 : DFFS_X1 port map( D => n4135, CK => CLK, SN => RESET_BAR,
                           Q => n11195, QN => n_3894);
   clk_r_REG3186_S2 : DFFS_X1 port map( D => n4140, CK => CLK, SN => RESET_BAR,
                           Q => n11194, QN => n_3895);
   clk_r_REG3184_S2 : DFFS_X1 port map( D => n4177, CK => CLK, SN => RESET_BAR,
                           Q => n11193, QN => n_3896);
   clk_r_REG3243_S2 : DFFS_X1 port map( D => n3991, CK => CLK, SN => RESET_BAR,
                           Q => n10101, QN => n_3897);
   clk_r_REG3241_S2 : DFFS_X1 port map( D => n3994, CK => CLK, SN => RESET_BAR,
                           Q => n10100, QN => n_3898);
   clk_r_REG3239_S2 : DFFS_X1 port map( D => n3997, CK => CLK, SN => RESET_BAR,
                           Q => n10099, QN => n_3899);
   clk_r_REG3237_S2 : DFFS_X1 port map( D => n4000, CK => CLK, SN => RESET_BAR,
                           Q => n10098, QN => n_3900);
   clk_r_REG3235_S2 : DFFS_X1 port map( D => n4005, CK => CLK, SN => RESET_BAR,
                           Q => n10097, QN => n_3901);
   clk_r_REG3233_S2 : DFFS_X1 port map( D => n4009, CK => CLK, SN => RESET_BAR,
                           Q => n10096, QN => n_3902);
   clk_r_REG3231_S2 : DFFS_X1 port map( D => n4034, CK => CLK, SN => RESET_BAR,
                           Q => n10095, QN => n_3903);
   clk_r_REG3229_S2 : DFFS_X1 port map( D => n4039, CK => CLK, SN => RESET_BAR,
                           Q => n10094, QN => n_3904);
   clk_r_REG3227_S2 : DFFS_X1 port map( D => n4043, CK => CLK, SN => RESET_BAR,
                           Q => n10093, QN => n_3905);
   clk_r_REG3225_S2 : DFFS_X1 port map( D => n4046, CK => CLK, SN => RESET_BAR,
                           Q => n10092, QN => n_3906);
   clk_r_REG3223_S2 : DFFS_X1 port map( D => n4049, CK => CLK, SN => RESET_BAR,
                           Q => n10091, QN => n_3907);
   clk_r_REG3221_S2 : DFFS_X1 port map( D => n4052, CK => CLK, SN => RESET_BAR,
                           Q => n10090, QN => n_3908);
   clk_r_REG3219_S2 : DFFS_X1 port map( D => n4055, CK => CLK, SN => RESET_BAR,
                           Q => n10089, QN => n_3909);
   clk_r_REG3217_S2 : DFFS_X1 port map( D => n4059, CK => CLK, SN => RESET_BAR,
                           Q => n10088, QN => n_3910);
   clk_r_REG3215_S2 : DFFS_X1 port map( D => n4063, CK => CLK, SN => RESET_BAR,
                           Q => n10087, QN => n_3911);
   clk_r_REG3213_S2 : DFFS_X1 port map( D => n4067, CK => CLK, SN => RESET_BAR,
                           Q => n10086, QN => n_3912);
   clk_r_REG3211_S2 : DFFS_X1 port map( D => n4071, CK => CLK, SN => RESET_BAR,
                           Q => n10085, QN => n_3913);
   clk_r_REG3209_S2 : DFFS_X1 port map( D => n4075, CK => CLK, SN => RESET_BAR,
                           Q => n10084, QN => n_3914);
   clk_r_REG3207_S2 : DFFS_X1 port map( D => n4079, CK => CLK, SN => RESET_BAR,
                           Q => n10083, QN => n_3915);
   clk_r_REG3205_S2 : DFFS_X1 port map( D => n4090, CK => CLK, SN => RESET_BAR,
                           Q => n10082, QN => n_3916);
   clk_r_REG3203_S2 : DFFS_X1 port map( D => n4094, CK => CLK, SN => RESET_BAR,
                           Q => n10081, QN => n_3917);
   clk_r_REG3201_S2 : DFFS_X1 port map( D => n4097, CK => CLK, SN => RESET_BAR,
                           Q => n10080, QN => n_3918);
   clk_r_REG3199_S2 : DFFS_X1 port map( D => n4102, CK => CLK, SN => RESET_BAR,
                           Q => n10079, QN => n_3919);
   clk_r_REG3197_S2 : DFFS_X1 port map( D => n4110, CK => CLK, SN => RESET_BAR,
                           Q => n10078, QN => n_3920);
   clk_r_REG3195_S2 : DFFS_X1 port map( D => n4115, CK => CLK, SN => RESET_BAR,
                           Q => n10077, QN => n_3921);
   clk_r_REG3193_S2 : DFFS_X1 port map( D => n4120, CK => CLK, SN => RESET_BAR,
                           Q => n10076, QN => n_3922);
   clk_r_REG3191_S2 : DFFS_X1 port map( D => n4125, CK => CLK, SN => RESET_BAR,
                           Q => n10075, QN => n_3923);
   clk_r_REG3189_S2 : DFFS_X1 port map( D => n4130, CK => CLK, SN => RESET_BAR,
                           Q => n10074, QN => n_3924);
   clk_r_REG3187_S2 : DFFS_X1 port map( D => n4135, CK => CLK, SN => RESET_BAR,
                           Q => n10073, QN => n_3925);
   clk_r_REG3185_S2 : DFFS_X1 port map( D => n4140, CK => CLK, SN => RESET_BAR,
                           Q => n10072, QN => n_3926);
   clk_r_REG3183_S2 : DFFS_X1 port map( D => n4177, CK => CLK, SN => RESET_BAR,
                           Q => n10071, QN => n_3927);
   clk_r_REG3245_S2 : DFFS_X1 port map( D => n3987, CK => CLK, SN => RESET_BAR,
                           Q => n10102, QN => n_3928);
   U3 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n11272, A3 => n11269, ZN => 
                           n15363);
   U4 : CLKBUF_X1 port map( A => n15363, Z => n15182);
   U5 : NAND3_X1 port map( A1 => RESET_BAR, A2 => n11272, A3 => n11270, ZN => 
                           n16090);
   U6 : CLKBUF_X1 port map( A => n16090, Z => n15905);
   U7 : INV_X1 port map( A => ADD_RD1(1), ZN => n13464);
   U8 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), ZN => n13461);
   U9 : NOR2_X1 port map( A1 => n13464, A2 => n13461, ZN => n3582);
   U10 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => n13461, ZN => n3581);
   U11 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => ADD_RD1(0)
                           , ZN => n3579);
   U12 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), A3 => ADD_RD2(0)
                           , ZN => n3589);
   U13 : NAND2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), ZN => n13462);
   U14 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => n13462, ZN => n3590);
   U15 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(0), A3 => n13464, ZN
                           => n3580);
   U16 : INV_X1 port map( A => ADD_RD2(2), ZN => n13468);
   U17 : NOR2_X1 port map( A1 => n13468, A2 => n13462, ZN => n3585);
   U18 : INV_X1 port map( A => ADD_RD1(2), ZN => n13465);
   U19 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => n13465, ZN
                           => n3578);
   U20 : INV_X1 port map( A => ADD_RD2(1), ZN => n13467);
   U21 : NOR3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => n13467, ZN
                           => n3588);
   U22 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n13465, ZN => n13463);
   U23 : NOR2_X1 port map( A1 => n13464, A2 => n13463, ZN => n3577);
   U24 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => n13463, ZN => n3575);
   U25 : INV_X1 port map( A => ADD_RD1(3), ZN => n3574);
   U26 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => n13465, A3 => n13464, ZN => 
                           n3576);
   U27 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n13467, ZN => n13466);
   U28 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => n13466, ZN => n3591);
   U29 : NOR2_X1 port map( A1 => n13468, A2 => n13466, ZN => n3584);
   U30 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => n13467, A3 => n13468, ZN => 
                           n3586);
   U31 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), A3 => n13468, ZN
                           => n3587);
   U32 : INV_X1 port map( A => ADD_RD2(3), ZN => n3583);
   U33 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11264, ZN => n14163);
   U34 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11222, ZN => n14408);
   U35 : OAI22_X1 port map( A1 => n11222, A2 => n14163, B1 => n10122, B2 => 
                           n14408, ZN => n13469);
   U36 : INV_X1 port map( A => n13469, ZN => n2562);
   U37 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11217, ZN => n14404);
   U38 : OAI22_X1 port map( A1 => n11217, A2 => n14163, B1 => n10121, B2 => 
                           n14404, ZN => n13470);
   U39 : INV_X1 port map( A => n13470, ZN => n2561);
   U40 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11215, ZN => n14410);
   U41 : OAI22_X1 port map( A1 => n11215, A2 => n14163, B1 => n10124, B2 => 
                           n14410, ZN => n13471);
   U42 : INV_X1 port map( A => n13471, ZN => n2564);
   U43 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11257, ZN => n14267);
   U44 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11220, ZN => n14365);
   U45 : OAI22_X1 port map( A1 => n11220, A2 => n14267, B1 => n10353, B2 => 
                           n14365, ZN => n13472);
   U46 : INV_X1 port map( A => n13472, ZN => n2781);
   U47 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11259, ZN => n14241);
   U48 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11221, ZN => n14358);
   U49 : OAI22_X1 port map( A1 => n11221, A2 => n14241, B1 => n10323, B2 => 
                           n14358, ZN => n13473);
   U50 : INV_X1 port map( A => n13473, ZN => n2718);
   U51 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11262, ZN => n14261);
   U52 : OAI22_X1 port map( A1 => n11220, A2 => n14261, B1 => n10202, B2 => 
                           n14365, ZN => n13474);
   U53 : INV_X1 port map( A => n13474, ZN => n2621);
   U54 : OAI22_X1 port map( A1 => n11221, A2 => n14261, B1 => n10201, B2 => 
                           n14358, ZN => n13475);
   U55 : INV_X1 port map( A => n13475, ZN => n2622);
   U56 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11219, ZN => n14406);
   U57 : OAI22_X1 port map( A1 => n11219, A2 => n14163, B1 => n10139, B2 => 
                           n14406, ZN => n13476);
   U58 : INV_X1 port map( A => n13476, ZN => n2559);
   U59 : OAI22_X1 port map( A1 => n11220, A2 => n14163, B1 => n10138, B2 => 
                           n14365, ZN => n13477);
   U60 : INV_X1 port map( A => n13477, ZN => n2558);
   U61 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11216, ZN => n14419);
   U62 : OAI22_X1 port map( A1 => n11216, A2 => n14163, B1 => n10123, B2 => 
                           n14419, ZN => n13478);
   U63 : INV_X1 port map( A => n13478, ZN => n2563);
   U64 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11218, ZN => n14422);
   U65 : OAI22_X1 port map( A1 => n11218, A2 => n14163, B1 => n10140, B2 => 
                           n14422, ZN => n13479);
   U66 : INV_X1 port map( A => n13479, ZN => n2560);
   U67 : OAI22_X1 port map( A1 => n11221, A2 => n14267, B1 => n10352, B2 => 
                           n14358, ZN => n13480);
   U68 : INV_X1 port map( A => n13480, ZN => n2782);
   U69 : OAI22_X1 port map( A1 => n11220, A2 => n14241, B1 => n10324, B2 => 
                           n14365, ZN => n13481);
   U70 : INV_X1 port map( A => n13481, ZN => n2717);
   U71 : OAI22_X1 port map( A1 => n11221, A2 => n14163, B1 => n10137, B2 => 
                           n14358, ZN => n13482);
   U72 : INV_X1 port map( A => n13482, ZN => n2557);
   U73 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11248, ZN => n14484);
   U74 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11193, ZN => n13921);
   U75 : OAI22_X1 port map( A1 => n10071, A2 => n14484, B1 => n10798, B2 => 
                           n13921, ZN => n13483);
   U76 : INV_X1 port map( A => n13483, ZN => n3092);
   U77 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11250, ZN => n14490);
   U78 : OAI22_X1 port map( A1 => n10071, A2 => n14490, B1 => n10416, B2 => 
                           n13921, ZN => n13484);
   U79 : INV_X1 port map( A => n13484, ZN => n3028);
   U80 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11197, ZN => n13900);
   U81 : OAI22_X1 port map( A1 => n11197, A2 => n14267, B1 => n10461, B2 => 
                           n13900, ZN => n13485);
   U82 : INV_X1 port map( A => n13485, ZN => n2800);
   U83 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11251, ZN => n14276);
   U84 : OAI22_X1 port map( A1 => n10071, A2 => n14276, B1 => n10526, B2 => 
                           n13921, ZN => n13486);
   U85 : INV_X1 port map( A => n13486, ZN => n2996);
   U86 : OAI22_X1 port map( A1 => n11197, A2 => n14241, B1 => n10307, B2 => 
                           n13900, ZN => n13487);
   U87 : INV_X1 port map( A => n13487, ZN => n2736);
   U88 : OAI22_X1 port map( A1 => n11197, A2 => n14261, B1 => n10166, B2 => 
                           n13900, ZN => n13488);
   U89 : INV_X1 port map( A => n13488, ZN => n2640);
   U90 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11252, ZN => n14274);
   U91 : OAI22_X1 port map( A1 => n10071, A2 => n14274, B1 => n10618, B2 => 
                           n13921, ZN => n13489);
   U92 : INV_X1 port map( A => n13489, ZN => n2964);
   U93 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11247, ZN => n14282);
   U94 : OAI22_X1 port map( A1 => n10071, A2 => n14282, B1 => n10767, B2 => 
                           n13921, ZN => n13490);
   U95 : INV_X1 port map( A => n13490, ZN => n3124);
   U96 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11254, ZN => n14271);
   U97 : OAI22_X1 port map( A1 => n11193, A2 => n14271, B1 => n10382, B2 => 
                           n13921, ZN => n13491);
   U98 : INV_X1 port map( A => n13491, ZN => n2900);
   U99 : OAI22_X1 port map( A1 => n11193, A2 => n14267, B1 => n10446, B2 => 
                           n13921, ZN => n13492);
   U100 : INV_X1 port map( A => n13492, ZN => n2804);
   U101 : OAI22_X1 port map( A1 => n11193, A2 => n14241, B1 => n10291, B2 => 
                           n13921, ZN => n13493);
   U102 : INV_X1 port map( A => n13493, ZN => n2740);
   U103 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11241, ZN => n14220);
   U104 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11198, ZN => n14414);
   U105 : OAI22_X1 port map( A1 => n10076, A2 => n14220, B1 => n10992, B2 => 
                           n14414, ZN => n13494);
   U106 : INV_X1 port map( A => n13494, ZN => n3311);
   U107 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11242, ZN => n14218);
   U108 : OAI22_X1 port map( A1 => n11198, A2 => n14218, B1 => n10962, B2 => 
                           n14414, ZN => n13495);
   U109 : INV_X1 port map( A => n13495, ZN => n3279);
   U110 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11244, ZN => n14210);
   U111 : OAI22_X1 port map( A1 => n11198, A2 => n14210, B1 => n10902, B2 => 
                           n14414, ZN => n13496);
   U112 : INV_X1 port map( A => n13496, ZN => n3215);
   U113 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11245, ZN => n14287);
   U114 : OAI22_X1 port map( A1 => n10076, A2 => n14287, B1 => n10872, B2 => 
                           n14414, ZN => n13497);
   U115 : INV_X1 port map( A => n13497, ZN => n3183);
   U116 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11246, ZN => n14280);
   U117 : OAI22_X1 port map( A1 => n10076, A2 => n14280, B1 => n10842, B2 => 
                           n14414, ZN => n13498);
   U118 : INV_X1 port map( A => n13498, ZN => n3151);
   U119 : OAI22_X1 port map( A1 => n10076, A2 => n14282, B1 => n10762, B2 => 
                           n14414, ZN => n13499);
   U120 : INV_X1 port map( A => n13499, ZN => n3119);
   U121 : OAI22_X1 port map( A1 => n11193, A2 => n14261, B1 => n10170, B2 => 
                           n13921, ZN => n13500);
   U122 : INV_X1 port map( A => n13500, ZN => n2644);
   U123 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11249, ZN => n14285);
   U124 : OAI22_X1 port map( A1 => n10075, A2 => n14285, B1 => n10491, B2 => 
                           n13900, ZN => n13501);
   U125 : INV_X1 port map( A => n13501, ZN => n3056);
   U126 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11195, ZN => n13918);
   U127 : OAI22_X1 port map( A1 => n10073, A2 => n14490, B1 => n10414, B2 => 
                           n13918, ZN => n13502);
   U128 : INV_X1 port map( A => n13502, ZN => n3026);
   U129 : OAI22_X1 port map( A1 => n10076, A2 => n14484, B1 => n10793, B2 => 
                           n14414, ZN => n13503);
   U130 : INV_X1 port map( A => n13503, ZN => n3087);
   U131 : OAI22_X1 port map( A1 => n10076, A2 => n14285, B1 => n10490, B2 => 
                           n14414, ZN => n13504);
   U132 : INV_X1 port map( A => n13504, ZN => n3055);
   U133 : OAI22_X1 port map( A1 => n10076, A2 => n14490, B1 => n10431, B2 => 
                           n14414, ZN => n13505);
   U134 : INV_X1 port map( A => n13505, ZN => n3023);
   U135 : OAI22_X1 port map( A1 => n10076, A2 => n14276, B1 => n10521, B2 => 
                           n14414, ZN => n13506);
   U136 : INV_X1 port map( A => n13506, ZN => n2991);
   U137 : OAI22_X1 port map( A1 => n10076, A2 => n14274, B1 => n10613, B2 => 
                           n14414, ZN => n13507);
   U138 : INV_X1 port map( A => n13507, ZN => n2959);
   U139 : OAI22_X1 port map( A1 => n10075, A2 => n14484, B1 => n10794, B2 => 
                           n13900, ZN => n13508);
   U140 : INV_X1 port map( A => n13508, ZN => n3088);
   U141 : OAI22_X1 port map( A1 => n10075, A2 => n14490, B1 => n10432, B2 => 
                           n13900, ZN => n13509);
   U142 : INV_X1 port map( A => n13509, ZN => n3024);
   U143 : OAI22_X1 port map( A1 => n10075, A2 => n14282, B1 => n10763, B2 => 
                           n13900, ZN => n13510);
   U144 : INV_X1 port map( A => n13510, ZN => n3120);
   U145 : OAI22_X1 port map( A1 => n11198, A2 => n14271, B1 => n10398, B2 => 
                           n14414, ZN => n13511);
   U146 : INV_X1 port map( A => n13511, ZN => n2895);
   U147 : OAI22_X1 port map( A1 => n10075, A2 => n14280, B1 => n10823, B2 => 
                           n13900, ZN => n13512);
   U148 : INV_X1 port map( A => n13512, ZN => n3152);
   U149 : OAI22_X1 port map( A1 => n10075, A2 => n14287, B1 => n10873, B2 => 
                           n13900, ZN => n13513);
   U150 : INV_X1 port map( A => n13513, ZN => n3184);
   U151 : OAI22_X1 port map( A1 => n11197, A2 => n14210, B1 => n10903, B2 => 
                           n13900, ZN => n13514);
   U152 : INV_X1 port map( A => n13514, ZN => n3216);
   U153 : OAI22_X1 port map( A1 => n10075, A2 => n14276, B1 => n10522, B2 => 
                           n13900, ZN => n13515);
   U154 : INV_X1 port map( A => n13515, ZN => n2992);
   U155 : OAI22_X1 port map( A1 => n11197, A2 => n14218, B1 => n10963, B2 => 
                           n13900, ZN => n13516);
   U156 : INV_X1 port map( A => n13516, ZN => n3280);
   U157 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11194, ZN => n13916);
   U158 : OAI22_X1 port map( A1 => n10072, A2 => n14220, B1 => n10996, B2 => 
                           n13916, ZN => n13517);
   U159 : INV_X1 port map( A => n13517, ZN => n3315);
   U160 : OAI22_X1 port map( A1 => n11194, A2 => n14218, B1 => n10966, B2 => 
                           n13916, ZN => n13518);
   U161 : INV_X1 port map( A => n13518, ZN => n3283);
   U162 : OAI22_X1 port map( A1 => n10075, A2 => n14274, B1 => n10614, B2 => 
                           n13900, ZN => n13519);
   U163 : INV_X1 port map( A => n13519, ZN => n2960);
   U164 : OAI22_X1 port map( A1 => n11194, A2 => n14210, B1 => n10886, B2 => 
                           n13916, ZN => n13520);
   U165 : INV_X1 port map( A => n13520, ZN => n3219);
   U166 : OAI22_X1 port map( A1 => n10072, A2 => n14287, B1 => n10856, B2 => 
                           n13916, ZN => n13521);
   U167 : INV_X1 port map( A => n13521, ZN => n3187);
   U168 : OAI22_X1 port map( A1 => n11197, A2 => n14271, B1 => n10399, B2 => 
                           n13900, ZN => n13522);
   U169 : INV_X1 port map( A => n13522, ZN => n2896);
   U170 : OAI22_X1 port map( A1 => n10072, A2 => n14280, B1 => n10826, B2 => 
                           n13916, ZN => n13523);
   U171 : INV_X1 port map( A => n13523, ZN => n3155);
   U172 : OAI22_X1 port map( A1 => n10072, A2 => n14282, B1 => n10766, B2 => 
                           n13916, ZN => n13524);
   U173 : INV_X1 port map( A => n13524, ZN => n3123);
   U174 : OAI22_X1 port map( A1 => n10075, A2 => n14220, B1 => n10993, B2 => 
                           n13900, ZN => n13525);
   U175 : INV_X1 port map( A => n13525, ZN => n3312);
   U176 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11196, ZN => n13912);
   U177 : OAI22_X1 port map( A1 => n11196, A2 => n14261, B1 => n10167, B2 => 
                           n13912, ZN => n13526);
   U178 : INV_X1 port map( A => n13526, ZN => n2641);
   U179 : OAI22_X1 port map( A1 => n11196, A2 => n14241, B1 => n10288, B2 => 
                           n13912, ZN => n13527);
   U180 : INV_X1 port map( A => n13527, ZN => n2737);
   U181 : OAI22_X1 port map( A1 => n11196, A2 => n14267, B1 => n10462, B2 => 
                           n13912, ZN => n13528);
   U182 : INV_X1 port map( A => n13528, ZN => n2801);
   U183 : OAI22_X1 port map( A1 => n11196, A2 => n14271, B1 => n10400, B2 => 
                           n13912, ZN => n13529);
   U184 : INV_X1 port map( A => n13529, ZN => n2897);
   U185 : OAI22_X1 port map( A1 => n10074, A2 => n14274, B1 => n10615, B2 => 
                           n13912, ZN => n13530);
   U186 : INV_X1 port map( A => n13530, ZN => n2961);
   U187 : OAI22_X1 port map( A1 => n10074, A2 => n14276, B1 => n10523, B2 => 
                           n13912, ZN => n13531);
   U188 : INV_X1 port map( A => n13531, ZN => n2993);
   U189 : OAI22_X1 port map( A1 => n10072, A2 => n14484, B1 => n10797, B2 => 
                           n13916, ZN => n13532);
   U190 : INV_X1 port map( A => n13532, ZN => n3091);
   U191 : OAI22_X1 port map( A1 => n10072, A2 => n14285, B1 => n10494, B2 => 
                           n13916, ZN => n13533);
   U192 : INV_X1 port map( A => n13533, ZN => n3059);
   U193 : OAI22_X1 port map( A1 => n10072, A2 => n14490, B1 => n10415, B2 => 
                           n13916, ZN => n13534);
   U194 : INV_X1 port map( A => n13534, ZN => n3027);
   U195 : OAI22_X1 port map( A1 => n10071, A2 => n14285, B1 => n10495, B2 => 
                           n13921, ZN => n13535);
   U196 : INV_X1 port map( A => n13535, ZN => n3060);
   U197 : OAI22_X1 port map( A1 => n10072, A2 => n14276, B1 => n10525, B2 => 
                           n13916, ZN => n13536);
   U198 : INV_X1 port map( A => n13536, ZN => n2995);
   U199 : OAI22_X1 port map( A1 => n10073, A2 => n14220, B1 => n10995, B2 => 
                           n13918, ZN => n13537);
   U200 : INV_X1 port map( A => n13537, ZN => n3314);
   U201 : OAI22_X1 port map( A1 => n10072, A2 => n14274, B1 => n10617, B2 => 
                           n13916, ZN => n13538);
   U202 : INV_X1 port map( A => n13538, ZN => n2963);
   U203 : OAI22_X1 port map( A1 => n11196, A2 => n14210, B1 => n10904, B2 => 
                           n13912, ZN => n13539);
   U204 : INV_X1 port map( A => n13539, ZN => n3217);
   U205 : OAI22_X1 port map( A1 => n11196, A2 => n14218, B1 => n10964, B2 => 
                           n13912, ZN => n13540);
   U206 : INV_X1 port map( A => n13540, ZN => n3281);
   U207 : OAI22_X1 port map( A1 => n10074, A2 => n14490, B1 => n10433, B2 => 
                           n13912, ZN => n13541);
   U208 : INV_X1 port map( A => n13541, ZN => n3025);
   U209 : OAI22_X1 port map( A1 => n10074, A2 => n14220, B1 => n10994, B2 => 
                           n13912, ZN => n13542);
   U210 : INV_X1 port map( A => n13542, ZN => n3313);
   U211 : OAI22_X1 port map( A1 => n10074, A2 => n14285, B1 => n10492, B2 => 
                           n13912, ZN => n13543);
   U212 : INV_X1 port map( A => n13543, ZN => n3057);
   U213 : OAI22_X1 port map( A1 => n11194, A2 => n14271, B1 => n10402, B2 => 
                           n13916, ZN => n13544);
   U214 : INV_X1 port map( A => n13544, ZN => n2899);
   U215 : OAI22_X1 port map( A1 => n10074, A2 => n14484, B1 => n10795, B2 => 
                           n13912, ZN => n13545);
   U216 : INV_X1 port map( A => n13545, ZN => n3089);
   U217 : OAI22_X1 port map( A1 => n11195, A2 => n14241, B1 => n10289, B2 => 
                           n13918, ZN => n13546);
   U218 : INV_X1 port map( A => n13546, ZN => n2738);
   U219 : OAI22_X1 port map( A1 => n10074, A2 => n14282, B1 => n10764, B2 => 
                           n13912, ZN => n13547);
   U220 : INV_X1 port map( A => n13547, ZN => n3121);
   U221 : OAI22_X1 port map( A1 => n11195, A2 => n14218, B1 => n10965, B2 => 
                           n13918, ZN => n13548);
   U222 : INV_X1 port map( A => n13548, ZN => n3282);
   U223 : OAI22_X1 port map( A1 => n10074, A2 => n14280, B1 => n10824, B2 => 
                           n13912, ZN => n13549);
   U224 : INV_X1 port map( A => n13549, ZN => n3153);
   U225 : OAI22_X1 port map( A1 => n11194, A2 => n14267, B1 => n10445, B2 => 
                           n13916, ZN => n13550);
   U226 : INV_X1 port map( A => n13550, ZN => n2803);
   U227 : OAI22_X1 port map( A1 => n10073, A2 => n14287, B1 => n10855, B2 => 
                           n13918, ZN => n13551);
   U228 : INV_X1 port map( A => n13551, ZN => n3186);
   U229 : OAI22_X1 port map( A1 => n10071, A2 => n14280, B1 => n10827, B2 => 
                           n13921, ZN => n13552);
   U230 : INV_X1 port map( A => n13552, ZN => n3156);
   U231 : OAI22_X1 port map( A1 => n11194, A2 => n14261, B1 => n10169, B2 => 
                           n13916, ZN => n13553);
   U232 : INV_X1 port map( A => n13553, ZN => n2643);
   U233 : OAI22_X1 port map( A1 => n10073, A2 => n14276, B1 => n10524, B2 => 
                           n13918, ZN => n13554);
   U234 : INV_X1 port map( A => n13554, ZN => n2994);
   U235 : OAI22_X1 port map( A1 => n10071, A2 => n14287, B1 => n10857, B2 => 
                           n13921, ZN => n13555);
   U236 : INV_X1 port map( A => n13555, ZN => n3188);
   U237 : OAI22_X1 port map( A1 => n10073, A2 => n14484, B1 => n10796, B2 => 
                           n13918, ZN => n13556);
   U238 : INV_X1 port map( A => n13556, ZN => n3090);
   U239 : OAI22_X1 port map( A1 => n10073, A2 => n14274, B1 => n10616, B2 => 
                           n13918, ZN => n13557);
   U240 : INV_X1 port map( A => n13557, ZN => n2962);
   U241 : OAI22_X1 port map( A1 => n11195, A2 => n14267, B1 => n10463, B2 => 
                           n13918, ZN => n13558);
   U242 : INV_X1 port map( A => n13558, ZN => n2802);
   U243 : OAI22_X1 port map( A1 => n11193, A2 => n14210, B1 => n10887, B2 => 
                           n13921, ZN => n13559);
   U244 : INV_X1 port map( A => n13559, ZN => n3220);
   U245 : OAI22_X1 port map( A1 => n11193, A2 => n14218, B1 => n10947, B2 => 
                           n13921, ZN => n13560);
   U246 : INV_X1 port map( A => n13560, ZN => n3284);
   U247 : OAI22_X1 port map( A1 => n10073, A2 => n14285, B1 => n10493, B2 => 
                           n13918, ZN => n13561);
   U248 : INV_X1 port map( A => n13561, ZN => n3058);
   U249 : OAI22_X1 port map( A1 => n10071, A2 => n14220, B1 => n10997, B2 => 
                           n13921, ZN => n13562);
   U250 : INV_X1 port map( A => n13562, ZN => n3316);
   U251 : OAI22_X1 port map( A1 => n10074, A2 => n14287, B1 => n10854, B2 => 
                           n13912, ZN => n13563);
   U252 : INV_X1 port map( A => n13563, ZN => n3185);
   U253 : OAI22_X1 port map( A1 => n11195, A2 => n14271, B1 => n10401, B2 => 
                           n13918, ZN => n13564);
   U254 : INV_X1 port map( A => n13564, ZN => n2898);
   U255 : OAI22_X1 port map( A1 => n11194, A2 => n14241, B1 => n10290, B2 => 
                           n13916, ZN => n13565);
   U256 : INV_X1 port map( A => n13565, ZN => n2739);
   U257 : OAI22_X1 port map( A1 => n11195, A2 => n14261, B1 => n10168, B2 => 
                           n13918, ZN => n13566);
   U258 : INV_X1 port map( A => n13566, ZN => n2642);
   U259 : OAI22_X1 port map( A1 => n11195, A2 => n14210, B1 => n10885, B2 => 
                           n13918, ZN => n13567);
   U260 : INV_X1 port map( A => n13567, ZN => n3218);
   U261 : OAI22_X1 port map( A1 => n10073, A2 => n14282, B1 => n10765, B2 => 
                           n13918, ZN => n13568);
   U262 : INV_X1 port map( A => n13568, ZN => n3122);
   U263 : OAI22_X1 port map( A1 => n10073, A2 => n14280, B1 => n10825, B2 => 
                           n13918, ZN => n13569);
   U264 : INV_X1 port map( A => n13569, ZN => n3154);
   U265 : CLKBUF_X1 port map( A => n14218, Z => n14125);
   U266 : OAI22_X1 port map( A1 => n11221, A2 => n14125, B1 => n10978, B2 => 
                           n14358, ZN => n13570);
   U267 : INV_X1 port map( A => n13570, ZN => n3260);
   U268 : OAI22_X1 port map( A1 => n11218, A2 => n14125, B1 => n10981, B2 => 
                           n14422, ZN => n13571);
   U269 : INV_X1 port map( A => n13571, ZN => n3257);
   U270 : OAI22_X1 port map( A1 => n11219, A2 => n14125, B1 => n10980, B2 => 
                           n14406, ZN => n13572);
   U271 : INV_X1 port map( A => n13572, ZN => n3258);
   U272 : OAI22_X1 port map( A1 => n11217, A2 => n14125, B1 => n10982, B2 => 
                           n14404, ZN => n13573);
   U273 : INV_X1 port map( A => n13573, ZN => n3256);
   U274 : OAI22_X1 port map( A1 => n11220, A2 => n14125, B1 => n10979, B2 => 
                           n14365, ZN => n13574);
   U275 : INV_X1 port map( A => n13574, ZN => n3259);
   U276 : OAI22_X1 port map( A1 => n11222, A2 => n14125, B1 => n10983, B2 => 
                           n14408, ZN => n13575);
   U277 : INV_X1 port map( A => n13575, ZN => n3255);
   U278 : OAI22_X1 port map( A1 => n11215, A2 => n14125, B1 => n10985, B2 => 
                           n14410, ZN => n13576);
   U279 : INV_X1 port map( A => n13576, ZN => n3253);
   U280 : OAI22_X1 port map( A1 => n11216, A2 => n14125, B1 => n10984, B2 => 
                           n14419, ZN => n13577);
   U281 : INV_X1 port map( A => n13577, ZN => n3254);
   U282 : CLKBUF_X1 port map( A => n14267, Z => n14253);
   U283 : OAI22_X1 port map( A1 => n11216, A2 => n14253, B1 => n10358, B2 => 
                           n14419, ZN => n13578);
   U284 : INV_X1 port map( A => n13578, ZN => n2776);
   U285 : OAI22_X1 port map( A1 => n11222, A2 => n14253, B1 => n10357, B2 => 
                           n14408, ZN => n13579);
   U286 : INV_X1 port map( A => n13579, ZN => n2777);
   U287 : OAI22_X1 port map( A1 => n11198, A2 => n14253, B1 => n10460, B2 => 
                           n14414, ZN => n13580);
   U288 : INV_X1 port map( A => n13580, ZN => n2799);
   U289 : OAI22_X1 port map( A1 => n11218, A2 => n14253, B1 => n10355, B2 => 
                           n14422, ZN => n13581);
   U290 : INV_X1 port map( A => n13581, ZN => n2779);
   U291 : OAI22_X1 port map( A1 => n11219, A2 => n14253, B1 => n10354, B2 => 
                           n14406, ZN => n13582);
   U292 : INV_X1 port map( A => n13582, ZN => n2780);
   U293 : OAI22_X1 port map( A1 => n11215, A2 => n14253, B1 => n10359, B2 => 
                           n14410, ZN => n13583);
   U294 : INV_X1 port map( A => n13583, ZN => n2775);
   U295 : OAI22_X1 port map( A1 => n11217, A2 => n14253, B1 => n10356, B2 => 
                           n14404, ZN => n13584);
   U296 : INV_X1 port map( A => n13584, ZN => n2778);
   U297 : CLKBUF_X1 port map( A => n14220, Z => n14127);
   U298 : OAI22_X1 port map( A1 => n10095, A2 => n14127, B1 => n11016, B2 => 
                           n14410, ZN => n13585);
   U299 : INV_X1 port map( A => n13585, ZN => n3285);
   U300 : OAI22_X1 port map( A1 => n10098, A2 => n14127, B1 => n11013, B2 => 
                           n14404, ZN => n13586);
   U301 : INV_X1 port map( A => n13586, ZN => n3288);
   U302 : OAI22_X1 port map( A1 => n10100, A2 => n14127, B1 => n11011, B2 => 
                           n14406, ZN => n13587);
   U303 : INV_X1 port map( A => n13587, ZN => n3290);
   U304 : OAI22_X1 port map( A1 => n11221, A2 => n14127, B1 => n11009, B2 => 
                           n14358, ZN => n13588);
   U305 : INV_X1 port map( A => n13588, ZN => n3292);
   U306 : OAI22_X1 port map( A1 => n10101, A2 => n14127, B1 => n11010, B2 => 
                           n14365, ZN => n13589);
   U307 : INV_X1 port map( A => n13589, ZN => n3291);
   U308 : OAI22_X1 port map( A1 => n10099, A2 => n14127, B1 => n11012, B2 => 
                           n14422, ZN => n13590);
   U309 : INV_X1 port map( A => n13590, ZN => n3289);
   U310 : OAI22_X1 port map( A1 => n10097, A2 => n14127, B1 => n11014, B2 => 
                           n14408, ZN => n13591);
   U311 : INV_X1 port map( A => n13591, ZN => n3287);
   U312 : OAI22_X1 port map( A1 => n10096, A2 => n14127, B1 => n11015, B2 => 
                           n14419, ZN => n13592);
   U313 : INV_X1 port map( A => n13592, ZN => n3286);
   U314 : CLKBUF_X1 port map( A => n14261, Z => n14122);
   U315 : OAI22_X1 port map( A1 => n11215, A2 => n14122, B1 => n10188, B2 => 
                           n14410, ZN => n13593);
   U316 : INV_X1 port map( A => n13593, ZN => n2615);
   U317 : OAI22_X1 port map( A1 => n11216, A2 => n14122, B1 => n10187, B2 => 
                           n14419, ZN => n13594);
   U318 : INV_X1 port map( A => n13594, ZN => n2616);
   U319 : OAI22_X1 port map( A1 => n11222, A2 => n14122, B1 => n10186, B2 => 
                           n14408, ZN => n13595);
   U320 : INV_X1 port map( A => n13595, ZN => n2617);
   U321 : CLKBUF_X1 port map( A => n14163, Z => n14229);
   U322 : OAI22_X1 port map( A1 => n11194, A2 => n14229, B1 => n10106, B2 => 
                           n13916, ZN => n13596);
   U323 : INV_X1 port map( A => n13596, ZN => n2550);
   U324 : OAI22_X1 port map( A1 => n11217, A2 => n14122, B1 => n10185, B2 => 
                           n14404, ZN => n13597);
   U325 : INV_X1 port map( A => n13597, ZN => n2618);
   U326 : OAI22_X1 port map( A1 => n11218, A2 => n14122, B1 => n10184, B2 => 
                           n14422, ZN => n13598);
   U327 : INV_X1 port map( A => n13598, ZN => n2619);
   U328 : OAI22_X1 port map( A1 => n11219, A2 => n14122, B1 => n10183, B2 => 
                           n14406, ZN => n13599);
   U329 : INV_X1 port map( A => n13599, ZN => n2620);
   U330 : CLKBUF_X1 port map( A => n14241, Z => n14093);
   U331 : OAI22_X1 port map( A1 => n11216, A2 => n14093, B1 => n10308, B2 => 
                           n14419, ZN => n13600);
   U332 : INV_X1 port map( A => n13600, ZN => n2712);
   U333 : OAI22_X1 port map( A1 => n11215, A2 => n14093, B1 => n10309, B2 => 
                           n14410, ZN => n13601);
   U334 : INV_X1 port map( A => n13601, ZN => n2711);
   U335 : CLKBUF_X1 port map( A => n14282, Z => n14171);
   U336 : OAI22_X1 port map( A1 => n10100, A2 => n14171, B1 => n10800, B2 => 
                           n14406, ZN => n13602);
   U337 : INV_X1 port map( A => n13602, ZN => n3098);
   U338 : OAI22_X1 port map( A1 => n10101, A2 => n14171, B1 => n10799, B2 => 
                           n14365, ZN => n13603);
   U339 : INV_X1 port map( A => n13603, ZN => n3099);
   U340 : OAI22_X1 port map( A1 => n10095, A2 => n14171, B1 => n10786, B2 => 
                           n14410, ZN => n13604);
   U341 : INV_X1 port map( A => n13604, ZN => n3093);
   U342 : OAI22_X1 port map( A1 => n10096, A2 => n14171, B1 => n10785, B2 => 
                           n14419, ZN => n13605);
   U343 : INV_X1 port map( A => n13605, ZN => n3094);
   U344 : CLKBUF_X1 port map( A => n14484, Z => n14169);
   U345 : OAI22_X1 port map( A1 => n10102, A2 => n14169, B1 => n10828, B2 => 
                           n14358, ZN => n13606);
   U346 : INV_X1 port map( A => n13606, ZN => n3068);
   U347 : OAI22_X1 port map( A1 => n10097, A2 => n14171, B1 => n10784, B2 => 
                           n14408, ZN => n13607);
   U348 : INV_X1 port map( A => n13607, ZN => n3095);
   U349 : OAI22_X1 port map( A1 => n10098, A2 => n14171, B1 => n10783, B2 => 
                           n14404, ZN => n13608);
   U350 : INV_X1 port map( A => n13608, ZN => n3096);
   U351 : OAI22_X1 port map( A1 => n10099, A2 => n14171, B1 => n10782, B2 => 
                           n14422, ZN => n13609);
   U352 : INV_X1 port map( A => n13609, ZN => n3097);
   U353 : OAI22_X1 port map( A1 => n11196, A2 => n14229, B1 => n10104, B2 => 
                           n13912, ZN => n13610);
   U354 : INV_X1 port map( A => n13610, ZN => n2552);
   U355 : OAI22_X1 port map( A1 => n11219, A2 => n14093, B1 => n10325, B2 => 
                           n14406, ZN => n13611);
   U356 : INV_X1 port map( A => n13611, ZN => n2716);
   U357 : OAI22_X1 port map( A1 => n11218, A2 => n14093, B1 => n10326, B2 => 
                           n14422, ZN => n13612);
   U358 : INV_X1 port map( A => n13612, ZN => n2715);
   U359 : OAI22_X1 port map( A1 => n11217, A2 => n14093, B1 => n10327, B2 => 
                           n14404, ZN => n13613);
   U360 : INV_X1 port map( A => n13613, ZN => n2714);
   U361 : OAI22_X1 port map( A1 => n11222, A2 => n14093, B1 => n10328, B2 => 
                           n14408, ZN => n13614);
   U362 : INV_X1 port map( A => n13614, ZN => n2713);
   U363 : OAI22_X1 port map( A1 => n11197, A2 => n14229, B1 => n10103, B2 => 
                           n13900, ZN => n13615);
   U364 : INV_X1 port map( A => n13615, ZN => n2553);
   U365 : CLKBUF_X1 port map( A => n14280, Z => n14173);
   U366 : OAI22_X1 port map( A1 => n10097, A2 => n14173, B1 => n10843, B2 => 
                           n14408, ZN => n13616);
   U367 : INV_X1 port map( A => n13616, ZN => n3127);
   U368 : OAI22_X1 port map( A1 => n10096, A2 => n14173, B1 => n10844, B2 => 
                           n14419, ZN => n13617);
   U369 : INV_X1 port map( A => n13617, ZN => n3126);
   U370 : OAI22_X1 port map( A1 => n10095, A2 => n14173, B1 => n10845, B2 => 
                           n14410, ZN => n13618);
   U371 : INV_X1 port map( A => n13618, ZN => n3125);
   U372 : OAI22_X1 port map( A1 => n11195, A2 => n14229, B1 => n10105, B2 => 
                           n13918, ZN => n13619);
   U373 : INV_X1 port map( A => n13619, ZN => n2551);
   U374 : OAI22_X1 port map( A1 => n11198, A2 => n14093, B1 => n10306, B2 => 
                           n14414, ZN => n13620);
   U375 : INV_X1 port map( A => n13620, ZN => n2735);
   U376 : OAI22_X1 port map( A1 => n11198, A2 => n14122, B1 => n10165, B2 => 
                           n14414, ZN => n13621);
   U377 : INV_X1 port map( A => n13621, ZN => n2639);
   U378 : OAI22_X1 port map( A1 => n10102, A2 => n14173, B1 => n10858, B2 => 
                           n14358, ZN => n13622);
   U379 : INV_X1 port map( A => n13622, ZN => n3132);
   U380 : OAI22_X1 port map( A1 => n10101, A2 => n14173, B1 => n10859, B2 => 
                           n14365, ZN => n13623);
   U381 : INV_X1 port map( A => n13623, ZN => n3131);
   U382 : OAI22_X1 port map( A1 => n10100, A2 => n14173, B1 => n10860, B2 => 
                           n14406, ZN => n13624);
   U383 : INV_X1 port map( A => n13624, ZN => n3130);
   U384 : OAI22_X1 port map( A1 => n10099, A2 => n14173, B1 => n10861, B2 => 
                           n14422, ZN => n13625);
   U385 : INV_X1 port map( A => n13625, ZN => n3129);
   U386 : OAI22_X1 port map( A1 => n10098, A2 => n14173, B1 => n10862, B2 => 
                           n14404, ZN => n13626);
   U387 : INV_X1 port map( A => n13626, ZN => n3128);
   U388 : CLKBUF_X1 port map( A => n14287, Z => n14131);
   U389 : OAI22_X1 port map( A1 => n10096, A2 => n14131, B1 => n10874, B2 => 
                           n14419, ZN => n13627);
   U390 : INV_X1 port map( A => n13627, ZN => n3158);
   U391 : OAI22_X1 port map( A1 => n10095, A2 => n14131, B1 => n10875, B2 => 
                           n14410, ZN => n13628);
   U392 : INV_X1 port map( A => n13628, ZN => n3157);
   U393 : CLKBUF_X1 port map( A => n14276, Z => n14167);
   U394 : OAI22_X1 port map( A1 => n10102, A2 => n14167, B1 => n11125, B2 => 
                           n14358, ZN => n13629);
   U395 : INV_X1 port map( A => n13629, ZN => n2972);
   U396 : OAI22_X1 port map( A1 => n11193, A2 => n14229, B1 => n11124, B2 => 
                           n13921, ZN => n13630);
   U397 : INV_X1 port map( A => n13630, ZN => n2549);
   U398 : OAI22_X1 port map( A1 => n11221, A2 => n14131, B1 => n10888, B2 => 
                           n14358, ZN => n13631);
   U399 : INV_X1 port map( A => n13631, ZN => n3164);
   U400 : OAI22_X1 port map( A1 => n10101, A2 => n14131, B1 => n10889, B2 => 
                           n14365, ZN => n13632);
   U401 : INV_X1 port map( A => n13632, ZN => n3163);
   U402 : OAI22_X1 port map( A1 => n10100, A2 => n14131, B1 => n10890, B2 => 
                           n14406, ZN => n13633);
   U403 : INV_X1 port map( A => n13633, ZN => n3162);
   U404 : OAI22_X1 port map( A1 => n10099, A2 => n14131, B1 => n10891, B2 => 
                           n14422, ZN => n13634);
   U405 : INV_X1 port map( A => n13634, ZN => n3161);
   U406 : OAI22_X1 port map( A1 => n10098, A2 => n14131, B1 => n10892, B2 => 
                           n14404, ZN => n13635);
   U407 : INV_X1 port map( A => n13635, ZN => n3160);
   U408 : OAI22_X1 port map( A1 => n10097, A2 => n14131, B1 => n10893, B2 => 
                           n14408, ZN => n13636);
   U409 : INV_X1 port map( A => n13636, ZN => n3159);
   U410 : CLKBUF_X1 port map( A => n14490, Z => n14224);
   U411 : OAI22_X1 port map( A1 => n10102, A2 => n14224, B1 => n10447, B2 => 
                           n14358, ZN => n13637);
   U412 : INV_X1 port map( A => n13637, ZN => n3004);
   U413 : OAI22_X1 port map( A1 => n11198, A2 => n14229, B1 => n11122, B2 => 
                           n14414, ZN => n13638);
   U414 : INV_X1 port map( A => n13638, ZN => n2554);
   U415 : CLKBUF_X1 port map( A => n14210, Z => n14129);
   U416 : OAI22_X1 port map( A1 => n11215, A2 => n14129, B1 => n10905, B2 => 
                           n14410, ZN => n13639);
   U417 : INV_X1 port map( A => n13639, ZN => n3189);
   U418 : OAI22_X1 port map( A1 => n11221, A2 => n14129, B1 => n10918, B2 => 
                           n14358, ZN => n13640);
   U419 : INV_X1 port map( A => n13640, ZN => n3196);
   U420 : OAI22_X1 port map( A1 => n11220, A2 => n14129, B1 => n10919, B2 => 
                           n14365, ZN => n13641);
   U421 : INV_X1 port map( A => n13641, ZN => n3195);
   U422 : OAI22_X1 port map( A1 => n11219, A2 => n14129, B1 => n10920, B2 => 
                           n14406, ZN => n13642);
   U423 : INV_X1 port map( A => n13642, ZN => n3194);
   U424 : OAI22_X1 port map( A1 => n11218, A2 => n14129, B1 => n10921, B2 => 
                           n14422, ZN => n13643);
   U425 : INV_X1 port map( A => n13643, ZN => n3193);
   U426 : CLKBUF_X1 port map( A => n14274, Z => n14165);
   U427 : OAI22_X1 port map( A1 => n10102, A2 => n14165, B1 => n10648, B2 => 
                           n14358, ZN => n13644);
   U428 : INV_X1 port map( A => n13644, ZN => n2940);
   U429 : OAI22_X1 port map( A1 => n11217, A2 => n14129, B1 => n10922, B2 => 
                           n14404, ZN => n13645);
   U430 : INV_X1 port map( A => n13645, ZN => n3192);
   U431 : OAI22_X1 port map( A1 => n11222, A2 => n14129, B1 => n10923, B2 => 
                           n14408, ZN => n13646);
   U432 : INV_X1 port map( A => n13646, ZN => n3191);
   U433 : CLKBUF_X1 port map( A => n14285, Z => n14247);
   U434 : OAI22_X1 port map( A1 => n10101, A2 => n14247, B1 => n10508, B2 => 
                           n14365, ZN => n13647);
   U435 : INV_X1 port map( A => n13647, ZN => n3035);
   U436 : OAI22_X1 port map( A1 => n10100, A2 => n14247, B1 => n10509, B2 => 
                           n14406, ZN => n13648);
   U437 : INV_X1 port map( A => n13648, ZN => n3034);
   U438 : OAI22_X1 port map( A1 => n10099, A2 => n14247, B1 => n10510, B2 => 
                           n14422, ZN => n13649);
   U439 : INV_X1 port map( A => n13649, ZN => n3033);
   U440 : OAI22_X1 port map( A1 => n10098, A2 => n14247, B1 => n10511, B2 => 
                           n14404, ZN => n13650);
   U441 : INV_X1 port map( A => n13650, ZN => n3032);
   U442 : OAI22_X1 port map( A1 => n10097, A2 => n14247, B1 => n10512, B2 => 
                           n14408, ZN => n13651);
   U443 : INV_X1 port map( A => n13651, ZN => n3031);
   U444 : OAI22_X1 port map( A1 => n10096, A2 => n14247, B1 => n10513, B2 => 
                           n14419, ZN => n13652);
   U445 : INV_X1 port map( A => n13652, ZN => n3030);
   U446 : OAI22_X1 port map( A1 => n11216, A2 => n14129, B1 => n10924, B2 => 
                           n14419, ZN => n13653);
   U447 : INV_X1 port map( A => n13653, ZN => n3190);
   U448 : OAI22_X1 port map( A1 => n10095, A2 => n14247, B1 => n10514, B2 => 
                           n14410, ZN => n13654);
   U449 : INV_X1 port map( A => n13654, ZN => n3029);
   U450 : CLKBUF_X1 port map( A => n14271, Z => n14195);
   U451 : OAI22_X1 port map( A1 => n10102, A2 => n14195, B1 => n10538, B2 => 
                           n14358, ZN => n13655);
   U452 : INV_X1 port map( A => n13655, ZN => n2876);
   U453 : OAI22_X1 port map( A1 => n10101, A2 => n14165, B1 => n10649, B2 => 
                           n14365, ZN => n13656);
   U454 : INV_X1 port map( A => n13656, ZN => n2939);
   U455 : OAI22_X1 port map( A1 => n11220, A2 => n14195, B1 => n10539, B2 => 
                           n14365, ZN => n13657);
   U456 : INV_X1 port map( A => n13657, ZN => n2875);
   U457 : OAI22_X1 port map( A1 => n11219, A2 => n14195, B1 => n10540, B2 => 
                           n14406, ZN => n13658);
   U458 : INV_X1 port map( A => n13658, ZN => n2874);
   U459 : OAI22_X1 port map( A1 => n10098, A2 => n14165, B1 => n10632, B2 => 
                           n14404, ZN => n13659);
   U460 : INV_X1 port map( A => n13659, ZN => n2936);
   U461 : OAI22_X1 port map( A1 => n11218, A2 => n14195, B1 => n10541, B2 => 
                           n14422, ZN => n13660);
   U462 : INV_X1 port map( A => n13660, ZN => n2873);
   U463 : OAI22_X1 port map( A1 => n11217, A2 => n14195, B1 => n10542, B2 => 
                           n14404, ZN => n13661);
   U464 : INV_X1 port map( A => n13661, ZN => n2872);
   U465 : OAI22_X1 port map( A1 => n11222, A2 => n14195, B1 => n10543, B2 => 
                           n14408, ZN => n13662);
   U466 : INV_X1 port map( A => n13662, ZN => n2871);
   U467 : OAI22_X1 port map( A1 => n11216, A2 => n14195, B1 => n10544, B2 => 
                           n14419, ZN => n13663);
   U468 : INV_X1 port map( A => n13663, ZN => n2870);
   U469 : OAI22_X1 port map( A1 => n11215, A2 => n14195, B1 => n10545, B2 => 
                           n14410, ZN => n13664);
   U470 : INV_X1 port map( A => n13664, ZN => n2869);
   U471 : OAI22_X1 port map( A1 => n10101, A2 => n14167, B1 => n10600, B2 => 
                           n14365, ZN => n13665);
   U472 : INV_X1 port map( A => n13665, ZN => n2971);
   U473 : OAI22_X1 port map( A1 => n10100, A2 => n14167, B1 => n10601, B2 => 
                           n14406, ZN => n13666);
   U474 : INV_X1 port map( A => n13666, ZN => n2970);
   U475 : OAI22_X1 port map( A1 => n10099, A2 => n14167, B1 => n10602, B2 => 
                           n14422, ZN => n13667);
   U476 : INV_X1 port map( A => n13667, ZN => n2969);
   U477 : OAI22_X1 port map( A1 => n10098, A2 => n14167, B1 => n10603, B2 => 
                           n14404, ZN => n13668);
   U478 : INV_X1 port map( A => n13668, ZN => n2968);
   U479 : OAI22_X1 port map( A1 => n10097, A2 => n14167, B1 => n10604, B2 => 
                           n14408, ZN => n13669);
   U480 : INV_X1 port map( A => n13669, ZN => n2967);
   U481 : OAI22_X1 port map( A1 => n10096, A2 => n14167, B1 => n10605, B2 => 
                           n14419, ZN => n13670);
   U482 : INV_X1 port map( A => n13670, ZN => n2966);
   U483 : OAI22_X1 port map( A1 => n10095, A2 => n14167, B1 => n10606, B2 => 
                           n14410, ZN => n13671);
   U484 : INV_X1 port map( A => n13671, ZN => n2965);
   U485 : OAI22_X1 port map( A1 => n10100, A2 => n14165, B1 => n10630, B2 => 
                           n14406, ZN => n13672);
   U486 : INV_X1 port map( A => n13672, ZN => n2938);
   U487 : OAI22_X1 port map( A1 => n10099, A2 => n14165, B1 => n10631, B2 => 
                           n14422, ZN => n13673);
   U488 : INV_X1 port map( A => n13673, ZN => n2937);
   U489 : OAI22_X1 port map( A1 => n10095, A2 => n14165, B1 => n10635, B2 => 
                           n14410, ZN => n13674);
   U490 : INV_X1 port map( A => n13674, ZN => n2933);
   U491 : OAI22_X1 port map( A1 => n10097, A2 => n14165, B1 => n10633, B2 => 
                           n14408, ZN => n13675);
   U492 : INV_X1 port map( A => n13675, ZN => n2935);
   U493 : OAI22_X1 port map( A1 => n10096, A2 => n14165, B1 => n10634, B2 => 
                           n14419, ZN => n13676);
   U494 : INV_X1 port map( A => n13676, ZN => n2934);
   U495 : CLKBUF_X1 port map( A => n14414, Z => n13844);
   U496 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11233, ZN => n14479);
   U497 : OAI22_X1 port map( A1 => n10151, A2 => n13844, B1 => n10076, B2 => 
                           n14479, ZN => n13677);
   U498 : INV_X1 port map( A => n13677, ZN => n3567);
   U499 : CLKBUF_X1 port map( A => n13916, Z => n13846);
   U500 : OAI22_X1 port map( A1 => n10135, A2 => n13846, B1 => n10072, B2 => 
                           n14479, ZN => n13678);
   U501 : INV_X1 port map( A => n13678, ZN => n3571);
   U502 : CLKBUF_X1 port map( A => n13918, Z => n13850);
   U503 : OAI22_X1 port map( A1 => n10134, A2 => n13850, B1 => n10073, B2 => 
                           n14479, ZN => n13679);
   U504 : INV_X1 port map( A => n13679, ZN => n3570);
   U505 : CLKBUF_X1 port map( A => n13900, Z => n13852);
   U506 : OAI22_X1 port map( A1 => n10132, A2 => n13852, B1 => n10075, B2 => 
                           n14479, ZN => n13680);
   U507 : INV_X1 port map( A => n13680, ZN => n3568);
   U508 : CLKBUF_X1 port map( A => n13921, Z => n13848);
   U509 : OAI22_X1 port map( A1 => n10136, A2 => n13848, B1 => n10071, B2 => 
                           n14479, ZN => n13681);
   U510 : INV_X1 port map( A => n13681, ZN => n3572);
   U511 : CLKBUF_X1 port map( A => n13912, Z => n13842);
   U512 : OAI22_X1 port map( A1 => n10133, A2 => n13842, B1 => n10074, B2 => 
                           n14479, ZN => n13682);
   U513 : INV_X1 port map( A => n13682, ZN => n3569);
   U514 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11238, ZN => n14573);
   U515 : CLKBUF_X1 port map( A => n14573, Z => n14502);
   U516 : CLKBUF_X1 port map( A => n14408, Z => n14323);
   U517 : OAI22_X1 port map( A1 => n10097, A2 => n14502, B1 => n11105, B2 => 
                           n14323, ZN => n13683);
   U518 : INV_X1 port map( A => n13683, ZN => n3383);
   U519 : CLKBUF_X1 port map( A => n14404, Z => n14314);
   U520 : OAI22_X1 port map( A1 => n10098, A2 => n14502, B1 => n11104, B2 => 
                           n14314, ZN => n13684);
   U521 : INV_X1 port map( A => n13684, ZN => n3384);
   U522 : CLKBUF_X1 port map( A => n14419, Z => n14316);
   U523 : OAI22_X1 port map( A1 => n10096, A2 => n14502, B1 => n11106, B2 => 
                           n14316, ZN => n13685);
   U524 : INV_X1 port map( A => n13685, ZN => n3382);
   U525 : CLKBUF_X1 port map( A => n14422, Z => n14327);
   U526 : OAI22_X1 port map( A1 => n10099, A2 => n14502, B1 => n11103, B2 => 
                           n14327, ZN => n13686);
   U527 : INV_X1 port map( A => n13686, ZN => n3385);
   U528 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11239, ZN => n14610);
   U529 : CLKBUF_X1 port map( A => n14610, Z => n14508);
   U530 : OAI22_X1 port map( A1 => n10099, A2 => n14508, B1 => n11073, B2 => 
                           n14327, ZN => n13687);
   U531 : INV_X1 port map( A => n13687, ZN => n3353);
   U532 : OAI22_X1 port map( A1 => n10098, A2 => n14508, B1 => n11074, B2 => 
                           n14314, ZN => n13688);
   U533 : INV_X1 port map( A => n13688, ZN => n3352);
   U534 : OAI22_X1 port map( A1 => n10099, A2 => n14169, B1 => n10831, B2 => 
                           n14327, ZN => n13689);
   U535 : INV_X1 port map( A => n13689, ZN => n3065);
   U536 : OAI22_X1 port map( A1 => n10097, A2 => n14508, B1 => n11075, B2 => 
                           n14323, ZN => n13690);
   U537 : INV_X1 port map( A => n13690, ZN => n3351);
   U538 : OAI22_X1 port map( A1 => n10096, A2 => n14508, B1 => n11076, B2 => 
                           n14316, ZN => n13691);
   U539 : INV_X1 port map( A => n13691, ZN => n3350);
   U540 : CLKBUF_X1 port map( A => n14410, Z => n14318);
   U541 : OAI22_X1 port map( A1 => n10095, A2 => n14508, B1 => n11077, B2 => 
                           n14318, ZN => n13692);
   U542 : INV_X1 port map( A => n13692, ZN => n3349);
   U543 : OAI22_X1 port map( A1 => n10095, A2 => n14502, B1 => n11107, B2 => 
                           n14318, ZN => n13693);
   U544 : INV_X1 port map( A => n13693, ZN => n3381);
   U545 : OAI22_X1 port map( A1 => n10095, A2 => n14169, B1 => n10815, B2 => 
                           n14318, ZN => n13694);
   U546 : INV_X1 port map( A => n13694, ZN => n3061);
   U547 : OAI22_X1 port map( A1 => n10096, A2 => n14169, B1 => n10814, B2 => 
                           n14316, ZN => n13695);
   U548 : INV_X1 port map( A => n13695, ZN => n3062);
   U549 : CLKBUF_X1 port map( A => n14406, Z => n14332);
   U550 : OAI22_X1 port map( A1 => n10100, A2 => n14502, B1 => n11102, B2 => 
                           n14332, ZN => n13696);
   U551 : INV_X1 port map( A => n13696, ZN => n3386);
   U552 : OAI22_X1 port map( A1 => n10100, A2 => n14508, B1 => n11072, B2 => 
                           n14332, ZN => n13697);
   U553 : INV_X1 port map( A => n13697, ZN => n3354);
   U554 : OAI22_X1 port map( A1 => n10097, A2 => n14169, B1 => n10813, B2 => 
                           n14323, ZN => n13698);
   U555 : INV_X1 port map( A => n13698, ZN => n3063);
   U556 : OAI22_X1 port map( A1 => n10098, A2 => n14169, B1 => n10812, B2 => 
                           n14314, ZN => n13699);
   U557 : INV_X1 port map( A => n13699, ZN => n3064);
   U558 : OAI22_X1 port map( A1 => n10100, A2 => n14169, B1 => n10830, B2 => 
                           n14332, ZN => n13700);
   U559 : INV_X1 port map( A => n13700, ZN => n3066);
   U560 : CLKBUF_X1 port map( A => n14358, Z => n14330);
   U561 : OAI22_X1 port map( A1 => n10102, A2 => n14502, B1 => n11120, B2 => 
                           n14330, ZN => n13701);
   U562 : INV_X1 port map( A => n13701, ZN => n3388);
   U563 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11236, ZN => n14599);
   U564 : CLKBUF_X1 port map( A => n14599, Z => n14511);
   U565 : OAI22_X1 port map( A1 => n10099, A2 => n14511, B1 => n10749, B2 => 
                           n14327, ZN => n13702);
   U566 : INV_X1 port map( A => n13702, ZN => n3449);
   U567 : OAI22_X1 port map( A1 => n10100, A2 => n14511, B1 => n10748, B2 => 
                           n14332, ZN => n13703);
   U568 : INV_X1 port map( A => n13703, ZN => n3450);
   U569 : CLKBUF_X1 port map( A => n14365, Z => n14320);
   U570 : OAI22_X1 port map( A1 => n10101, A2 => n14502, B1 => n11121, B2 => 
                           n14320, ZN => n13704);
   U571 : INV_X1 port map( A => n13704, ZN => n3387);
   U572 : OAI22_X1 port map( A1 => n10101, A2 => n14508, B1 => n11071, B2 => 
                           n14320, ZN => n13705);
   U573 : INV_X1 port map( A => n13705, ZN => n3355);
   U574 : OAI22_X1 port map( A1 => n10101, A2 => n14511, B1 => n10747, B2 => 
                           n14320, ZN => n13706);
   U575 : INV_X1 port map( A => n13706, ZN => n3451);
   U576 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11237, ZN => n14604);
   U577 : CLKBUF_X1 port map( A => n14604, Z => n14516);
   U578 : OAI22_X1 port map( A1 => n10096, A2 => n14516, B1 => n10702, B2 => 
                           n14316, ZN => n13707);
   U579 : INV_X1 port map( A => n13707, ZN => n3414);
   U580 : OAI22_X1 port map( A1 => n10097, A2 => n14516, B1 => n10701, B2 => 
                           n14323, ZN => n13708);
   U581 : INV_X1 port map( A => n13708, ZN => n3415);
   U582 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11235, ZN => n14594);
   U583 : CLKBUF_X1 port map( A => n14594, Z => n14505);
   U584 : OAI22_X1 port map( A1 => n10096, A2 => n14505, B1 => n10340, B2 => 
                           n14316, ZN => n13709);
   U585 : INV_X1 port map( A => n13709, ZN => n3478);
   U586 : OAI22_X1 port map( A1 => n10095, A2 => n14505, B1 => n10341, B2 => 
                           n14318, ZN => n13710);
   U587 : INV_X1 port map( A => n13710, ZN => n3477);
   U588 : OAI22_X1 port map( A1 => n10101, A2 => n14169, B1 => n10829, B2 => 
                           n14320, ZN => n13711);
   U589 : INV_X1 port map( A => n13711, ZN => n3067);
   U590 : OAI22_X1 port map( A1 => n10102, A2 => n14516, B1 => n10716, B2 => 
                           n14330, ZN => n13712);
   U591 : INV_X1 port map( A => n13712, ZN => n3420);
   U592 : OAI22_X1 port map( A1 => n10101, A2 => n14505, B1 => n10418, B2 => 
                           n14320, ZN => n13713);
   U593 : INV_X1 port map( A => n13713, ZN => n3483);
   U594 : OAI22_X1 port map( A1 => n10095, A2 => n14511, B1 => n10733, B2 => 
                           n14318, ZN => n13714);
   U595 : INV_X1 port map( A => n13714, ZN => n3445);
   U596 : OAI22_X1 port map( A1 => n10096, A2 => n14511, B1 => n10732, B2 => 
                           n14316, ZN => n13715);
   U597 : INV_X1 port map( A => n13715, ZN => n3446);
   U598 : OAI22_X1 port map( A1 => n10097, A2 => n14511, B1 => n10731, B2 => 
                           n14323, ZN => n13716);
   U599 : INV_X1 port map( A => n13716, ZN => n3447);
   U600 : OAI22_X1 port map( A1 => n10098, A2 => n14511, B1 => n10730, B2 => 
                           n14314, ZN => n13717);
   U601 : INV_X1 port map( A => n13717, ZN => n3448);
   U602 : OAI22_X1 port map( A1 => n10100, A2 => n14516, B1 => n10718, B2 => 
                           n14332, ZN => n13718);
   U603 : INV_X1 port map( A => n13718, ZN => n3418);
   U604 : OAI22_X1 port map( A1 => n10101, A2 => n14516, B1 => n10717, B2 => 
                           n14320, ZN => n13719);
   U605 : INV_X1 port map( A => n13719, ZN => n3419);
   U606 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11234, ZN => n14591);
   U607 : CLKBUF_X1 port map( A => n14591, Z => n14513);
   U608 : OAI22_X1 port map( A1 => n10096, A2 => n14513, B1 => n10673, B2 => 
                           n14316, ZN => n13720);
   U609 : INV_X1 port map( A => n13720, ZN => n3510);
   U610 : OAI22_X1 port map( A1 => n10100, A2 => n14505, B1 => n10419, B2 => 
                           n14332, ZN => n13721);
   U611 : INV_X1 port map( A => n13721, ZN => n3482);
   U612 : OAI22_X1 port map( A1 => n10102, A2 => n14505, B1 => n10417, B2 => 
                           n14330, ZN => n13722);
   U613 : INV_X1 port map( A => n13722, ZN => n3484);
   U614 : OAI22_X1 port map( A1 => n10102, A2 => n14511, B1 => n10746, B2 => 
                           n14330, ZN => n13723);
   U615 : INV_X1 port map( A => n13723, ZN => n3452);
   U616 : OAI22_X1 port map( A1 => n10097, A2 => n14513, B1 => n10672, B2 => 
                           n14323, ZN => n13724);
   U617 : INV_X1 port map( A => n13724, ZN => n3511);
   U618 : OAI22_X1 port map( A1 => n10098, A2 => n14516, B1 => n10700, B2 => 
                           n14314, ZN => n13725);
   U619 : INV_X1 port map( A => n13725, ZN => n3416);
   U620 : OAI22_X1 port map( A1 => n10102, A2 => n14508, B1 => n11090, B2 => 
                           n14330, ZN => n13726);
   U621 : INV_X1 port map( A => n13726, ZN => n3356);
   U622 : OAI22_X1 port map( A1 => n10098, A2 => n14513, B1 => n10687, B2 => 
                           n14314, ZN => n13727);
   U623 : INV_X1 port map( A => n13727, ZN => n3512);
   U624 : OAI22_X1 port map( A1 => n10099, A2 => n14513, B1 => n10686, B2 => 
                           n14327, ZN => n13728);
   U625 : INV_X1 port map( A => n13728, ZN => n3513);
   U626 : OAI22_X1 port map( A1 => n10100, A2 => n14513, B1 => n10685, B2 => 
                           n14332, ZN => n13729);
   U627 : INV_X1 port map( A => n13729, ZN => n3514);
   U628 : OAI22_X1 port map( A1 => n10101, A2 => n14513, B1 => n10684, B2 => 
                           n14320, ZN => n13730);
   U629 : INV_X1 port map( A => n13730, ZN => n3515);
   U630 : OAI22_X1 port map( A1 => n10099, A2 => n14505, B1 => n10420, B2 => 
                           n14327, ZN => n13731);
   U631 : INV_X1 port map( A => n13731, ZN => n3481);
   U632 : OAI22_X1 port map( A1 => n10102, A2 => n14171, B1 => n11126, B2 => 
                           n14330, ZN => n13732);
   U633 : INV_X1 port map( A => n13732, ZN => n3100);
   U634 : OAI22_X1 port map( A1 => n10098, A2 => n14505, B1 => n10421, B2 => 
                           n14314, ZN => n13733);
   U635 : INV_X1 port map( A => n13733, ZN => n3480);
   U636 : OAI22_X1 port map( A1 => n10097, A2 => n14505, B1 => n10422, B2 => 
                           n14323, ZN => n13734);
   U637 : INV_X1 port map( A => n13734, ZN => n3479);
   U638 : OAI22_X1 port map( A1 => n10095, A2 => n14516, B1 => n10703, B2 => 
                           n14318, ZN => n13735);
   U639 : INV_X1 port map( A => n13735, ZN => n3413);
   U640 : OAI22_X1 port map( A1 => n10099, A2 => n14224, B1 => n10450, B2 => 
                           n14327, ZN => n13736);
   U641 : INV_X1 port map( A => n13736, ZN => n3001);
   U642 : OAI22_X1 port map( A1 => n10095, A2 => n14513, B1 => n10674, B2 => 
                           n14318, ZN => n13737);
   U643 : INV_X1 port map( A => n13737, ZN => n3509);
   U644 : OAI22_X1 port map( A1 => n10098, A2 => n14224, B1 => n10451, B2 => 
                           n14314, ZN => n13738);
   U645 : INV_X1 port map( A => n13738, ZN => n3000);
   U646 : OAI22_X1 port map( A1 => n10099, A2 => n14516, B1 => n10699, B2 => 
                           n14327, ZN => n13739);
   U647 : INV_X1 port map( A => n13739, ZN => n3417);
   U648 : OAI22_X1 port map( A1 => n10096, A2 => n14224, B1 => n10453, B2 => 
                           n14316, ZN => n13740);
   U649 : INV_X1 port map( A => n13740, ZN => n2998);
   U650 : OAI22_X1 port map( A1 => n10102, A2 => n14247, B1 => n10507, B2 => 
                           n14330, ZN => n13741);
   U651 : INV_X1 port map( A => n13741, ZN => n3036);
   U652 : OAI22_X1 port map( A1 => n10095, A2 => n14224, B1 => n10434, B2 => 
                           n14318, ZN => n13742);
   U653 : INV_X1 port map( A => n13742, ZN => n2997);
   U654 : OAI22_X1 port map( A1 => n10102, A2 => n14513, B1 => n10683, B2 => 
                           n14330, ZN => n13743);
   U655 : INV_X1 port map( A => n13743, ZN => n3516);
   U656 : OAI22_X1 port map( A1 => n10101, A2 => n14224, B1 => n10448, B2 => 
                           n14320, ZN => n13744);
   U657 : INV_X1 port map( A => n13744, ZN => n3003);
   U658 : OAI22_X1 port map( A1 => n10100, A2 => n14224, B1 => n10449, B2 => 
                           n14332, ZN => n13745);
   U659 : INV_X1 port map( A => n13745, ZN => n3002);
   U660 : OAI22_X1 port map( A1 => n10097, A2 => n14224, B1 => n10452, B2 => 
                           n14323, ZN => n13746);
   U661 : INV_X1 port map( A => n13746, ZN => n2999);
   U662 : CLKBUF_X1 port map( A => n14479, Z => n14373);
   U663 : OAI22_X1 port map( A1 => n10294, A2 => n14332, B1 => n10100, B2 => 
                           n14373, ZN => n13747);
   U664 : INV_X1 port map( A => n13747, ZN => n3546);
   U665 : OAI22_X1 port map( A1 => n10153, A2 => n14316, B1 => n10096, B2 => 
                           n14373, ZN => n13748);
   U666 : INV_X1 port map( A => n13748, ZN => n3542);
   U667 : OAI22_X1 port map( A1 => n10292, A2 => n14330, B1 => n10102, B2 => 
                           n14373, ZN => n13749);
   U668 : INV_X1 port map( A => n13749, ZN => n3548);
   U669 : OAI22_X1 port map( A1 => n10293, A2 => n14320, B1 => n10101, B2 => 
                           n14373, ZN => n13750);
   U670 : INV_X1 port map( A => n13750, ZN => n3547);
   U671 : OAI22_X1 port map( A1 => n10295, A2 => n14327, B1 => n10099, B2 => 
                           n14373, ZN => n13751);
   U672 : INV_X1 port map( A => n13751, ZN => n3545);
   U673 : OAI22_X1 port map( A1 => n10152, A2 => n14323, B1 => n10097, B2 => 
                           n14373, ZN => n13752);
   U674 : INV_X1 port map( A => n13752, ZN => n3543);
   U675 : OAI22_X1 port map( A1 => n10296, A2 => n14314, B1 => n10098, B2 => 
                           n14373, ZN => n13753);
   U676 : INV_X1 port map( A => n13753, ZN => n3544);
   U677 : OAI22_X1 port map( A1 => n10154, A2 => n14318, B1 => n10095, B2 => 
                           n14373, ZN => n13754);
   U678 : INV_X1 port map( A => n13754, ZN => n3541);
   U679 : OAI22_X1 port map( A1 => n10073, A2 => n14599, B1 => n10713, B2 => 
                           n13850, ZN => n13755);
   U680 : INV_X1 port map( A => n13755, ZN => n3474);
   U681 : OAI22_X1 port map( A1 => n10071, A2 => n14610, B1 => n11059, B2 => 
                           n13848, ZN => n13756);
   U682 : INV_X1 port map( A => n13756, ZN => n3380);
   U683 : OAI22_X1 port map( A1 => n10072, A2 => n14591, B1 => n10744, B2 => 
                           n13846, ZN => n13757);
   U684 : INV_X1 port map( A => n13757, ZN => n3539);
   U685 : OAI22_X1 port map( A1 => n10076, A2 => n14573, B1 => n11084, B2 => 
                           n13844, ZN => n13758);
   U686 : INV_X1 port map( A => n13758, ZN => n3407);
   U687 : OAI22_X1 port map( A1 => n10071, A2 => n14573, B1 => n11089, B2 => 
                           n13848, ZN => n13759);
   U688 : INV_X1 port map( A => n13759, ZN => n3412);
   U689 : OAI22_X1 port map( A1 => n10071, A2 => n14604, B1 => n11119, B2 => 
                           n13848, ZN => n13760);
   U690 : INV_X1 port map( A => n13760, ZN => n3444);
   U691 : OAI22_X1 port map( A1 => n10071, A2 => n14599, B1 => n10715, B2 => 
                           n13848, ZN => n13761);
   U692 : INV_X1 port map( A => n13761, ZN => n3476);
   U693 : OAI22_X1 port map( A1 => n10071, A2 => n14594, B1 => n10322, B2 => 
                           n13848, ZN => n13762);
   U694 : INV_X1 port map( A => n13762, ZN => n3508);
   U695 : OAI22_X1 port map( A1 => n10076, A2 => n14591, B1 => n10671, B2 => 
                           n13844, ZN => n13763);
   U696 : INV_X1 port map( A => n13763, ZN => n3535);
   U697 : OAI22_X1 port map( A1 => n10071, A2 => n14591, B1 => n10745, B2 => 
                           n13848, ZN => n13764);
   U698 : INV_X1 port map( A => n13764, ZN => n3540);
   U699 : OAI22_X1 port map( A1 => n10073, A2 => n14610, B1 => n11057, B2 => 
                           n13850, ZN => n13765);
   U700 : INV_X1 port map( A => n13765, ZN => n3378);
   U701 : OAI22_X1 port map( A1 => n10074, A2 => n14610, B1 => n11056, B2 => 
                           n13842, ZN => n13766);
   U702 : INV_X1 port map( A => n13766, ZN => n3377);
   U703 : OAI22_X1 port map( A1 => n10072, A2 => n14594, B1 => n10321, B2 => 
                           n13846, ZN => n13767);
   U704 : INV_X1 port map( A => n13767, ZN => n3507);
   U705 : OAI22_X1 port map( A1 => n10073, A2 => n14591, B1 => n10743, B2 => 
                           n13850, ZN => n13768);
   U706 : INV_X1 port map( A => n13768, ZN => n3538);
   U707 : OAI22_X1 port map( A1 => n10073, A2 => n14594, B1 => n10320, B2 => 
                           n13850, ZN => n13769);
   U708 : INV_X1 port map( A => n13769, ZN => n3506);
   U709 : OAI22_X1 port map( A1 => n10072, A2 => n14599, B1 => n10714, B2 => 
                           n13846, ZN => n13770);
   U710 : INV_X1 port map( A => n13770, ZN => n3475);
   U711 : OAI22_X1 port map( A1 => n10074, A2 => n14591, B1 => n10742, B2 => 
                           n13842, ZN => n13771);
   U712 : INV_X1 port map( A => n13771, ZN => n3537);
   U713 : OAI22_X1 port map( A1 => n10072, A2 => n14604, B1 => n11118, B2 => 
                           n13846, ZN => n13772);
   U714 : INV_X1 port map( A => n13772, ZN => n3443);
   U715 : OAI22_X1 port map( A1 => n10072, A2 => n14573, B1 => n11088, B2 => 
                           n13846, ZN => n13773);
   U716 : INV_X1 port map( A => n13773, ZN => n3411);
   U717 : OAI22_X1 port map( A1 => n10072, A2 => n14610, B1 => n11058, B2 => 
                           n13846, ZN => n13774);
   U718 : INV_X1 port map( A => n13774, ZN => n3379);
   U719 : OAI22_X1 port map( A1 => n10074, A2 => n14604, B1 => n11116, B2 => 
                           n13842, ZN => n13775);
   U720 : INV_X1 port map( A => n13775, ZN => n3441);
   U721 : OAI22_X1 port map( A1 => n10074, A2 => n14573, B1 => n11086, B2 => 
                           n13842, ZN => n13776);
   U722 : INV_X1 port map( A => n13776, ZN => n3409);
   U723 : OAI22_X1 port map( A1 => n10075, A2 => n14604, B1 => n11115, B2 => 
                           n13852, ZN => n13777);
   U724 : INV_X1 port map( A => n13777, ZN => n3440);
   U725 : OAI22_X1 port map( A1 => n10073, A2 => n14573, B1 => n11087, B2 => 
                           n13850, ZN => n13778);
   U726 : INV_X1 port map( A => n13778, ZN => n3410);
   U727 : OAI22_X1 port map( A1 => n10075, A2 => n14594, B1 => n10339, B2 => 
                           n13852, ZN => n13779);
   U728 : INV_X1 port map( A => n13779, ZN => n3504);
   U729 : OAI22_X1 port map( A1 => n10076, A2 => n14604, B1 => n11114, B2 => 
                           n13844, ZN => n13780);
   U730 : INV_X1 port map( A => n13780, ZN => n3439);
   U731 : OAI22_X1 port map( A1 => n10073, A2 => n14604, B1 => n11117, B2 => 
                           n13850, ZN => n13781);
   U732 : INV_X1 port map( A => n13781, ZN => n3442);
   U733 : OAI22_X1 port map( A1 => n10076, A2 => n14610, B1 => n11054, B2 => 
                           n13844, ZN => n13782);
   U734 : INV_X1 port map( A => n13782, ZN => n3375);
   U735 : OAI22_X1 port map( A1 => n10075, A2 => n14599, B1 => n10711, B2 => 
                           n13852, ZN => n13783);
   U736 : INV_X1 port map( A => n13783, ZN => n3472);
   U737 : OAI22_X1 port map( A1 => n10075, A2 => n14610, B1 => n11055, B2 => 
                           n13852, ZN => n13784);
   U738 : INV_X1 port map( A => n13784, ZN => n3376);
   U739 : OAI22_X1 port map( A1 => n10076, A2 => n14594, B1 => n10338, B2 => 
                           n13844, ZN => n13785);
   U740 : INV_X1 port map( A => n13785, ZN => n3503);
   U741 : OAI22_X1 port map( A1 => n10076, A2 => n14599, B1 => n10710, B2 => 
                           n13844, ZN => n13786);
   U742 : INV_X1 port map( A => n13786, ZN => n3471);
   U743 : OAI22_X1 port map( A1 => n10075, A2 => n14573, B1 => n11085, B2 => 
                           n13852, ZN => n13787);
   U744 : INV_X1 port map( A => n13787, ZN => n3408);
   U745 : OAI22_X1 port map( A1 => n10075, A2 => n14591, B1 => n10741, B2 => 
                           n13852, ZN => n13788);
   U746 : INV_X1 port map( A => n13788, ZN => n3536);
   U747 : OAI22_X1 port map( A1 => n10074, A2 => n14599, B1 => n10712, B2 => 
                           n13842, ZN => n13789);
   U748 : INV_X1 port map( A => n13789, ZN => n3473);
   U749 : OAI22_X1 port map( A1 => n10074, A2 => n14594, B1 => n10319, B2 => 
                           n13842, ZN => n13790);
   U750 : INV_X1 port map( A => n13790, ZN => n3505);
   U751 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11243, ZN => n14295);
   U752 : OAI22_X1 port map( A1 => n11198, A2 => n14295, B1 => n10932, B2 => 
                           n14414, ZN => n13791);
   U753 : INV_X1 port map( A => n13791, ZN => n3247);
   U754 : OAI22_X1 port map( A1 => n11194, A2 => n14295, B1 => n10916, B2 => 
                           n13916, ZN => n13792);
   U755 : INV_X1 port map( A => n13792, ZN => n3251);
   U756 : OAI22_X1 port map( A1 => n11193, A2 => n14295, B1 => n10917, B2 => 
                           n13921, ZN => n13793);
   U757 : INV_X1 port map( A => n13793, ZN => n3252);
   U758 : OAI22_X1 port map( A1 => n11197, A2 => n14295, B1 => n10933, B2 => 
                           n13900, ZN => n13794);
   U759 : INV_X1 port map( A => n13794, ZN => n3248);
   U760 : OAI22_X1 port map( A1 => n11195, A2 => n14295, B1 => n10935, B2 => 
                           n13918, ZN => n13795);
   U761 : INV_X1 port map( A => n13795, ZN => n3250);
   U762 : OAI22_X1 port map( A1 => n11196, A2 => n14295, B1 => n10934, B2 => 
                           n13912, ZN => n13796);
   U763 : INV_X1 port map( A => n13796, ZN => n3249);
   U764 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11214, ZN => n14293);
   U765 : OAI22_X1 port map( A1 => n11214, A2 => n14163, B1 => n10125, B2 => 
                           n14293, ZN => n13797);
   U766 : INV_X1 port map( A => n13797, ZN => n2565);
   U767 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11213, ZN => n14289);
   U768 : OAI22_X1 port map( A1 => n11213, A2 => n14267, B1 => n10465, B2 => 
                           n14289, ZN => n13798);
   U769 : INV_X1 port map( A => n13798, ZN => n2784);
   U770 : OAI22_X1 port map( A1 => n11214, A2 => n14218, B1 => n10986, B2 => 
                           n14293, ZN => n13799);
   U771 : INV_X1 port map( A => n13799, ZN => n3261);
   U772 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11212, ZN => n14291);
   U773 : OAI22_X1 port map( A1 => n11212, A2 => n14295, B1 => n10938, B2 => 
                           n14291, ZN => n13800);
   U774 : INV_X1 port map( A => n13800, ZN => n3231);
   U775 : OAI22_X1 port map( A1 => n10094, A2 => n14276, B1 => n10607, B2 => 
                           n14293, ZN => n13801);
   U776 : INV_X1 port map( A => n13801, ZN => n2973);
   U777 : OAI22_X1 port map( A1 => n10092, A2 => n14280, B1 => n10848, B2 => 
                           n14291, ZN => n13802);
   U778 : INV_X1 port map( A => n13802, ZN => n3135);
   U779 : OAI22_X1 port map( A1 => n11214, A2 => n14261, B1 => n10189, B2 => 
                           n14293, ZN => n13803);
   U780 : INV_X1 port map( A => n13803, ZN => n2623);
   U781 : OAI22_X1 port map( A1 => n11212, A2 => n14261, B1 => n10191, B2 => 
                           n14291, ZN => n13804);
   U782 : INV_X1 port map( A => n13804, ZN => n2625);
   U783 : OAI22_X1 port map( A1 => n10092, A2 => n14220, B1 => n10998, B2 => 
                           n14291, ZN => n13805);
   U784 : INV_X1 port map( A => n13805, ZN => n3295);
   U785 : OAI22_X1 port map( A1 => n11214, A2 => n14241, B1 => n10310, B2 => 
                           n14293, ZN => n13806);
   U786 : INV_X1 port map( A => n13806, ZN => n2719);
   U787 : OAI22_X1 port map( A1 => n11213, A2 => n14210, B1 => n10907, B2 => 
                           n14289, ZN => n13807);
   U788 : INV_X1 port map( A => n13807, ZN => n3198);
   U789 : OAI22_X1 port map( A1 => n11212, A2 => n14218, B1 => n10968, B2 => 
                           n14291, ZN => n13808);
   U790 : INV_X1 port map( A => n13808, ZN => n3263);
   U791 : OAI22_X1 port map( A1 => n10093, A2 => n14280, B1 => n10847, B2 => 
                           n14289, ZN => n13809);
   U792 : INV_X1 port map( A => n13809, ZN => n3134);
   U793 : OAI22_X1 port map( A1 => n11212, A2 => n14210, B1 => n10908, B2 => 
                           n14291, ZN => n13810);
   U794 : INV_X1 port map( A => n13810, ZN => n3199);
   U795 : OAI22_X1 port map( A1 => n10092, A2 => n14287, B1 => n10878, B2 => 
                           n14291, ZN => n13811);
   U796 : INV_X1 port map( A => n13811, ZN => n3167);
   U797 : OAI22_X1 port map( A1 => n11214, A2 => n14271, B1 => n10546, B2 => 
                           n14293, ZN => n13812);
   U798 : INV_X1 port map( A => n13812, ZN => n2877);
   U799 : OAI22_X1 port map( A1 => n10094, A2 => n14285, B1 => n10515, B2 => 
                           n14293, ZN => n13813);
   U800 : INV_X1 port map( A => n13813, ZN => n3037);
   U801 : OAI22_X1 port map( A1 => n11213, A2 => n14261, B1 => n10190, B2 => 
                           n14289, ZN => n13814);
   U802 : INV_X1 port map( A => n13814, ZN => n2624);
   U803 : OAI22_X1 port map( A1 => n10092, A2 => n14282, B1 => n10789, B2 => 
                           n14291, ZN => n13815);
   U804 : INV_X1 port map( A => n13815, ZN => n3103);
   U805 : OAI22_X1 port map( A1 => n11213, A2 => n14163, B1 => n10126, B2 => 
                           n14289, ZN => n13816);
   U806 : INV_X1 port map( A => n13816, ZN => n2566);
   U807 : OAI22_X1 port map( A1 => n10092, A2 => n14285, B1 => n10517, B2 => 
                           n14291, ZN => n13817);
   U808 : INV_X1 port map( A => n13817, ZN => n3039);
   U809 : OAI22_X1 port map( A1 => n11214, A2 => n14267, B1 => n10464, B2 => 
                           n14293, ZN => n13818);
   U810 : INV_X1 port map( A => n13818, ZN => n2783);
   U811 : OAI22_X1 port map( A1 => n10094, A2 => n14280, B1 => n10846, B2 => 
                           n14293, ZN => n13819);
   U812 : INV_X1 port map( A => n13819, ZN => n3133);
   U813 : OAI22_X1 port map( A1 => n10094, A2 => n14274, B1 => n10636, B2 => 
                           n14293, ZN => n13820);
   U814 : INV_X1 port map( A => n13820, ZN => n2941);
   U815 : OAI22_X1 port map( A1 => n10092, A2 => n14276, B1 => n10609, B2 => 
                           n14291, ZN => n13821);
   U816 : INV_X1 port map( A => n13821, ZN => n2975);
   U817 : OAI22_X1 port map( A1 => n10092, A2 => n14274, B1 => n10638, B2 => 
                           n14291, ZN => n13822);
   U818 : INV_X1 port map( A => n13822, ZN => n2943);
   U819 : OAI22_X1 port map( A1 => n11212, A2 => n14271, B1 => n10404, B2 => 
                           n14291, ZN => n13823);
   U820 : INV_X1 port map( A => n13823, ZN => n2879);
   U821 : OAI22_X1 port map( A1 => n11214, A2 => n14295, B1 => n10936, B2 => 
                           n14293, ZN => n13824);
   U822 : INV_X1 port map( A => n13824, ZN => n3229);
   U823 : OAI22_X1 port map( A1 => n10093, A2 => n14274, B1 => n10637, B2 => 
                           n14289, ZN => n13825);
   U824 : INV_X1 port map( A => n13825, ZN => n2942);
   U825 : OAI22_X1 port map( A1 => n11212, A2 => n14267, B1 => n10466, B2 => 
                           n14291, ZN => n13826);
   U826 : INV_X1 port map( A => n13826, ZN => n2785);
   U827 : OAI22_X1 port map( A1 => n11214, A2 => n14210, B1 => n10906, B2 => 
                           n14293, ZN => n13827);
   U828 : INV_X1 port map( A => n13827, ZN => n3197);
   U829 : OAI22_X1 port map( A1 => n11212, A2 => n14241, B1 => n10312, B2 => 
                           n14291, ZN => n13828);
   U830 : INV_X1 port map( A => n13828, ZN => n2721);
   U831 : OAI22_X1 port map( A1 => n11213, A2 => n14241, B1 => n10311, B2 => 
                           n14289, ZN => n13829);
   U832 : INV_X1 port map( A => n13829, ZN => n2720);
   U833 : OAI22_X1 port map( A1 => n10093, A2 => n14285, B1 => n10516, B2 => 
                           n14289, ZN => n13830);
   U834 : INV_X1 port map( A => n13830, ZN => n3038);
   U835 : OAI22_X1 port map( A1 => n10093, A2 => n14276, B1 => n10608, B2 => 
                           n14289, ZN => n13831);
   U836 : INV_X1 port map( A => n13831, ZN => n2974);
   U837 : OAI22_X1 port map( A1 => n10094, A2 => n14220, B1 => n11017, B2 => 
                           n14293, ZN => n13832);
   U838 : INV_X1 port map( A => n13832, ZN => n3293);
   U839 : OAI22_X1 port map( A1 => n11213, A2 => n14218, B1 => n10967, B2 => 
                           n14289, ZN => n13833);
   U840 : INV_X1 port map( A => n13833, ZN => n3262);
   U841 : OAI22_X1 port map( A1 => n11213, A2 => n14295, B1 => n10937, B2 => 
                           n14289, ZN => n13834);
   U842 : INV_X1 port map( A => n13834, ZN => n3230);
   U843 : OAI22_X1 port map( A1 => n11212, A2 => n14163, B1 => n10127, B2 => 
                           n14291, ZN => n13835);
   U844 : INV_X1 port map( A => n13835, ZN => n2567);
   U845 : OAI22_X1 port map( A1 => n10094, A2 => n14282, B1 => n10787, B2 => 
                           n14293, ZN => n13836);
   U846 : INV_X1 port map( A => n13836, ZN => n3101);
   U847 : OAI22_X1 port map( A1 => n10093, A2 => n14220, B1 => n11018, B2 => 
                           n14289, ZN => n13837);
   U848 : INV_X1 port map( A => n13837, ZN => n3294);
   U849 : OAI22_X1 port map( A1 => n10093, A2 => n14282, B1 => n10788, B2 => 
                           n14289, ZN => n13838);
   U850 : INV_X1 port map( A => n13838, ZN => n3102);
   U851 : OAI22_X1 port map( A1 => n11213, A2 => n14271, B1 => n10403, B2 => 
                           n14289, ZN => n13839);
   U852 : INV_X1 port map( A => n13839, ZN => n2878);
   U853 : OAI22_X1 port map( A1 => n10094, A2 => n14287, B1 => n10876, B2 => 
                           n14293, ZN => n13840);
   U854 : INV_X1 port map( A => n13840, ZN => n3165);
   U855 : OAI22_X1 port map( A1 => n10093, A2 => n14287, B1 => n10877, B2 => 
                           n14289, ZN => n13841);
   U856 : INV_X1 port map( A => n13841, ZN => n3166);
   U857 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11240, ZN => n14619);
   U858 : OAI22_X1 port map( A1 => n10074, A2 => n14619, B1 => n11025, B2 => 
                           n13842, ZN => n13843);
   U859 : INV_X1 port map( A => n13843, ZN => n3345);
   U860 : OAI22_X1 port map( A1 => n10076, A2 => n14619, B1 => n11023, B2 => 
                           n13844, ZN => n13845);
   U861 : INV_X1 port map( A => n13845, ZN => n3343);
   U862 : OAI22_X1 port map( A1 => n10072, A2 => n14619, B1 => n11027, B2 => 
                           n13846, ZN => n13847);
   U863 : INV_X1 port map( A => n13847, ZN => n3347);
   U864 : OAI22_X1 port map( A1 => n10071, A2 => n14619, B1 => n11028, B2 => 
                           n13848, ZN => n13849);
   U865 : INV_X1 port map( A => n13849, ZN => n3348);
   U866 : OAI22_X1 port map( A1 => n10073, A2 => n14619, B1 => n11026, B2 => 
                           n13850, ZN => n13851);
   U867 : INV_X1 port map( A => n13851, ZN => n3346);
   U868 : OAI22_X1 port map( A1 => n10075, A2 => n14619, B1 => n11024, B2 => 
                           n13852, ZN => n13853);
   U869 : INV_X1 port map( A => n13853, ZN => n3344);
   U870 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11263, ZN => n14363);
   U871 : OAI22_X1 port map( A1 => n11214, A2 => n14363, B1 => n10219, B2 => 
                           n14293, ZN => n13854);
   U872 : INV_X1 port map( A => n13854, ZN => n2591);
   U873 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11260, ZN => n14384);
   U874 : OAI22_X1 port map( A1 => n11214, A2 => n14384, B1 => n10254, B2 => 
                           n14293, ZN => n13855);
   U875 : INV_X1 port map( A => n13855, ZN => n2687);
   U876 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11256, ZN => n14334);
   U877 : OAI22_X1 port map( A1 => n11197, A2 => n14334, B1 => n10584, B2 => 
                           n13900, ZN => n13856);
   U878 : INV_X1 port map( A => n13856, ZN => n2832);
   U879 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11258, ZN => n14344);
   U880 : OAI22_X1 port map( A1 => n11214, A2 => n14344, B1 => n10391, B2 => 
                           n14293, ZN => n13857);
   U881 : INV_X1 port map( A => n13857, ZN => n2751);
   U882 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11255, ZN => n14337);
   U883 : OAI22_X1 port map( A1 => n11197, A2 => n14337, B1 => n10553, B2 => 
                           n13900, ZN => n13858);
   U884 : INV_X1 port map( A => n13858, ZN => n2864);
   U885 : OAI22_X1 port map( A1 => n11214, A2 => n14334, B1 => n10483, B2 => 
                           n14293, ZN => n13859);
   U886 : INV_X1 port map( A => n13859, ZN => n2813);
   U887 : OAI22_X1 port map( A1 => n11214, A2 => n14337, B1 => n10577, B2 => 
                           n14293, ZN => n13860);
   U888 : INV_X1 port map( A => n13860, ZN => n2845);
   U889 : OAI22_X1 port map( A1 => n11213, A2 => n14363, B1 => n10220, B2 => 
                           n14289, ZN => n13861);
   U890 : INV_X1 port map( A => n13861, ZN => n2592);
   U891 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11261, ZN => n14375);
   U892 : OAI22_X1 port map( A1 => n11213, A2 => n14375, B1 => n10285, B2 => 
                           n14289, ZN => n13862);
   U893 : INV_X1 port map( A => n13862, ZN => n2656);
   U894 : OAI22_X1 port map( A1 => n11213, A2 => n14384, B1 => n10255, B2 => 
                           n14289, ZN => n13863);
   U895 : INV_X1 port map( A => n13863, ZN => n2688);
   U896 : OAI22_X1 port map( A1 => n11213, A2 => n14344, B1 => n10371, B2 => 
                           n14289, ZN => n13864);
   U897 : INV_X1 port map( A => n13864, ZN => n2752);
   U898 : OAI22_X1 port map( A1 => n11213, A2 => n14334, B1 => n10484, B2 => 
                           n14289, ZN => n13865);
   U899 : INV_X1 port map( A => n13865, ZN => n2814);
   U900 : OAI22_X1 port map( A1 => n11213, A2 => n14337, B1 => n10578, B2 => 
                           n14289, ZN => n13866);
   U901 : INV_X1 port map( A => n13866, ZN => n2846);
   U902 : OAI22_X1 port map( A1 => n11198, A2 => n14334, B1 => n10583, B2 => 
                           n14414, ZN => n13867);
   U903 : INV_X1 port map( A => n13867, ZN => n2831);
   U904 : OAI22_X1 port map( A1 => n11212, A2 => n14363, B1 => n10221, B2 => 
                           n14291, ZN => n13868);
   U905 : INV_X1 port map( A => n13868, ZN => n2593);
   U906 : OAI22_X1 port map( A1 => n11212, A2 => n14375, B1 => n10286, B2 => 
                           n14291, ZN => n13869);
   U907 : INV_X1 port map( A => n13869, ZN => n2657);
   U908 : OAI22_X1 port map( A1 => n11212, A2 => n14384, B1 => n10256, B2 => 
                           n14291, ZN => n13870);
   U909 : INV_X1 port map( A => n13870, ZN => n2689);
   U910 : OAI22_X1 port map( A1 => n11212, A2 => n14344, B1 => n10372, B2 => 
                           n14291, ZN => n13871);
   U911 : INV_X1 port map( A => n13871, ZN => n2753);
   U912 : OAI22_X1 port map( A1 => n11212, A2 => n14334, B1 => n10485, B2 => 
                           n14291, ZN => n13872);
   U913 : INV_X1 port map( A => n13872, ZN => n2815);
   U914 : OAI22_X1 port map( A1 => n11212, A2 => n14337, B1 => n10558, B2 => 
                           n14291, ZN => n13873);
   U915 : INV_X1 port map( A => n13873, ZN => n2847);
   U916 : OAI22_X1 port map( A1 => n11196, A2 => n14337, B1 => n10554, B2 => 
                           n13912, ZN => n13874);
   U917 : INV_X1 port map( A => n13874, ZN => n2865);
   U918 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11253, ZN => n14488);
   U919 : OAI22_X1 port map( A1 => n10074, A2 => n14488, B1 => n10644, B2 => 
                           n13912, ZN => n13875);
   U920 : INV_X1 port map( A => n13875, ZN => n2929);
   U921 : OAI22_X1 port map( A1 => n11195, A2 => n14363, B1 => n10198, B2 => 
                           n13918, ZN => n13876);
   U922 : INV_X1 port map( A => n13876, ZN => n2610);
   U923 : OAI22_X1 port map( A1 => n11195, A2 => n14375, B1 => n10263, B2 => 
                           n13918, ZN => n13877);
   U924 : INV_X1 port map( A => n13877, ZN => n2674);
   U925 : OAI22_X1 port map( A1 => n11195, A2 => n14384, B1 => n10232, B2 => 
                           n13918, ZN => n13878);
   U926 : INV_X1 port map( A => n13878, ZN => n2706);
   U927 : OAI22_X1 port map( A1 => n11195, A2 => n14344, B1 => n10369, B2 => 
                           n13918, ZN => n13879);
   U928 : INV_X1 port map( A => n13879, ZN => n2770);
   U929 : OAI22_X1 port map( A1 => n11221, A2 => n14363, B1 => n10107, B2 => 
                           n14358, ZN => n13880);
   U930 : INV_X1 port map( A => n13880, ZN => n2590);
   U931 : OAI22_X1 port map( A1 => n11221, A2 => n14375, B1 => n10171, B2 => 
                           n14358, ZN => n13881);
   U932 : INV_X1 port map( A => n13881, ZN => n2654);
   U933 : OAI22_X1 port map( A1 => n11221, A2 => n14384, B1 => n10246, B2 => 
                           n14358, ZN => n13882);
   U934 : INV_X1 port map( A => n13882, ZN => n2686);
   U935 : OAI22_X1 port map( A1 => n11221, A2 => n14344, B1 => n10383, B2 => 
                           n14358, ZN => n13883);
   U936 : INV_X1 port map( A => n13883, ZN => n2750);
   U937 : OAI22_X1 port map( A1 => n11214, A2 => n14375, B1 => n10284, B2 => 
                           n14293, ZN => n13884);
   U938 : INV_X1 port map( A => n13884, ZN => n2655);
   U939 : OAI22_X1 port map( A1 => n11220, A2 => n14384, B1 => n10247, B2 => 
                           n14365, ZN => n13885);
   U940 : INV_X1 port map( A => n13885, ZN => n2685);
   U941 : OAI22_X1 port map( A1 => n11198, A2 => n14337, B1 => n10552, B2 => 
                           n14414, ZN => n13886);
   U942 : INV_X1 port map( A => n13886, ZN => n2863);
   U943 : OAI22_X1 port map( A1 => n11195, A2 => n14337, B1 => n10555, B2 => 
                           n13918, ZN => n13887);
   U944 : INV_X1 port map( A => n13887, ZN => n2866);
   U945 : OAI22_X1 port map( A1 => n10076, A2 => n14488, B1 => n10642, B2 => 
                           n14414, ZN => n13888);
   U946 : INV_X1 port map( A => n13888, ZN => n2927);
   U947 : OAI22_X1 port map( A1 => n11197, A2 => n14363, B1 => n10196, B2 => 
                           n13900, ZN => n13889);
   U948 : INV_X1 port map( A => n13889, ZN => n2608);
   U949 : OAI22_X1 port map( A1 => n11197, A2 => n14375, B1 => n10261, B2 => 
                           n13900, ZN => n13890);
   U950 : INV_X1 port map( A => n13890, ZN => n2672);
   U951 : OAI22_X1 port map( A1 => n11197, A2 => n14384, B1 => n10230, B2 => 
                           n13900, ZN => n13891);
   U952 : INV_X1 port map( A => n13891, ZN => n2704);
   U953 : OAI22_X1 port map( A1 => n11197, A2 => n14344, B1 => n10367, B2 => 
                           n13900, ZN => n13892);
   U954 : INV_X1 port map( A => n13892, ZN => n2768);
   U955 : OAI22_X1 port map( A1 => n11194, A2 => n14384, B1 => n10233, B2 => 
                           n13916, ZN => n13893);
   U956 : INV_X1 port map( A => n13893, ZN => n2707);
   U957 : OAI22_X1 port map( A1 => n11194, A2 => n14344, B1 => n10370, B2 => 
                           n13916, ZN => n13894);
   U958 : INV_X1 port map( A => n13894, ZN => n2771);
   U959 : OAI22_X1 port map( A1 => n11194, A2 => n14334, B1 => n10587, B2 => 
                           n13916, ZN => n13895);
   U960 : INV_X1 port map( A => n13895, ZN => n2835);
   U961 : OAI22_X1 port map( A1 => n11194, A2 => n14337, B1 => n10556, B2 => 
                           n13916, ZN => n13896);
   U962 : INV_X1 port map( A => n13896, ZN => n2867);
   U963 : OAI22_X1 port map( A1 => n11194, A2 => n14375, B1 => n10264, B2 => 
                           n13916, ZN => n13897);
   U964 : INV_X1 port map( A => n13897, ZN => n2675);
   U965 : OAI22_X1 port map( A1 => n11196, A2 => n14375, B1 => n10262, B2 => 
                           n13912, ZN => n13898);
   U966 : INV_X1 port map( A => n13898, ZN => n2673);
   U967 : OAI22_X1 port map( A1 => n11193, A2 => n14384, B1 => n10234, B2 => 
                           n13921, ZN => n13899);
   U968 : INV_X1 port map( A => n13899, ZN => n2708);
   U969 : OAI22_X1 port map( A1 => n10075, A2 => n14488, B1 => n10643, B2 => 
                           n13900, ZN => n13901);
   U970 : INV_X1 port map( A => n13901, ZN => n2928);
   U971 : OAI22_X1 port map( A1 => n11220, A2 => n14363, B1 => n10108, B2 => 
                           n14365, ZN => n13902);
   U972 : INV_X1 port map( A => n13902, ZN => n2589);
   U973 : OAI22_X1 port map( A1 => n11220, A2 => n14375, B1 => n10277, B2 => 
                           n14365, ZN => n13903);
   U974 : INV_X1 port map( A => n13903, ZN => n2653);
   U975 : OAI22_X1 port map( A1 => n11193, A2 => n14337, B1 => n10557, B2 => 
                           n13921, ZN => n13904);
   U976 : INV_X1 port map( A => n13904, ZN => n2868);
   U977 : OAI22_X1 port map( A1 => n11220, A2 => n14344, B1 => n10384, B2 => 
                           n14365, ZN => n13905);
   U978 : INV_X1 port map( A => n13905, ZN => n2749);
   U979 : OAI22_X1 port map( A1 => n11196, A2 => n14363, B1 => n10197, B2 => 
                           n13912, ZN => n13906);
   U980 : INV_X1 port map( A => n13906, ZN => n2609);
   U981 : OAI22_X1 port map( A1 => n11196, A2 => n14334, B1 => n10585, B2 => 
                           n13912, ZN => n13907);
   U982 : INV_X1 port map( A => n13907, ZN => n2833);
   U983 : OAI22_X1 port map( A1 => n11193, A2 => n14334, B1 => n10588, B2 => 
                           n13921, ZN => n13908);
   U984 : INV_X1 port map( A => n13908, ZN => n2836);
   U985 : OAI22_X1 port map( A1 => n11193, A2 => n14375, B1 => n10265, B2 => 
                           n13921, ZN => n13909);
   U986 : INV_X1 port map( A => n13909, ZN => n2676);
   U987 : OAI22_X1 port map( A1 => n11195, A2 => n14334, B1 => n10586, B2 => 
                           n13918, ZN => n13910);
   U988 : INV_X1 port map( A => n13910, ZN => n2834);
   U989 : OAI22_X1 port map( A1 => n11196, A2 => n14384, B1 => n10231, B2 => 
                           n13912, ZN => n13911);
   U990 : INV_X1 port map( A => n13911, ZN => n2705);
   U991 : OAI22_X1 port map( A1 => n11196, A2 => n14344, B1 => n10368, B2 => 
                           n13912, ZN => n13913);
   U992 : INV_X1 port map( A => n13913, ZN => n2769);
   U993 : OAI22_X1 port map( A1 => n11194, A2 => n14363, B1 => n10199, B2 => 
                           n13916, ZN => n13914);
   U994 : INV_X1 port map( A => n13914, ZN => n2611);
   U995 : OAI22_X1 port map( A1 => n10071, A2 => n14488, B1 => n10647, B2 => 
                           n13921, ZN => n13915);
   U996 : INV_X1 port map( A => n13915, ZN => n2932);
   U997 : OAI22_X1 port map( A1 => n10072, A2 => n14488, B1 => n10646, B2 => 
                           n13916, ZN => n13917);
   U998 : INV_X1 port map( A => n13917, ZN => n2931);
   U999 : OAI22_X1 port map( A1 => n10073, A2 => n14488, B1 => n10645, B2 => 
                           n13918, ZN => n13919);
   U1000 : INV_X1 port map( A => n13919, ZN => n2930);
   U1001 : OAI22_X1 port map( A1 => n11193, A2 => n14344, B1 => n10351, B2 => 
                           n13921, ZN => n13920);
   U1002 : INV_X1 port map( A => n13920, ZN => n2772);
   U1003 : OAI22_X1 port map( A1 => n11193, A2 => n14363, B1 => n10200, B2 => 
                           n13921, ZN => n13922);
   U1004 : INV_X1 port map( A => n13922, ZN => n2612);
   U1005 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11211, ZN => n14308);
   U1006 : OAI22_X1 port map( A1 => n11211, A2 => n14363, B1 => n10222, B2 => 
                           n14308, ZN => n13923);
   U1007 : INV_X1 port map( A => n13923, ZN => n2594);
   U1008 : OAI22_X1 port map( A1 => n11211, A2 => n14384, B1 => n10235, B2 => 
                           n14308, ZN => n13924);
   U1009 : INV_X1 port map( A => n13924, ZN => n2690);
   U1010 : OAI22_X1 port map( A1 => n10091, A2 => n14274, B1 => n10639, B2 => 
                           n14308, ZN => n13925);
   U1011 : INV_X1 port map( A => n13925, ZN => n2944);
   U1012 : OAI22_X1 port map( A1 => n11211, A2 => n14261, B1 => n10192, B2 => 
                           n14308, ZN => n13926);
   U1013 : INV_X1 port map( A => n13926, ZN => n2626);
   U1014 : OAI22_X1 port map( A1 => n11211, A2 => n14344, B1 => n10373, B2 => 
                           n14308, ZN => n13927);
   U1015 : INV_X1 port map( A => n13927, ZN => n2754);
   U1016 : OAI22_X1 port map( A1 => n10091, A2 => n14287, B1 => n10879, B2 => 
                           n14308, ZN => n13928);
   U1017 : INV_X1 port map( A => n13928, ZN => n3168);
   U1018 : OAI22_X1 port map( A1 => n11211, A2 => n14210, B1 => n10909, B2 => 
                           n14308, ZN => n13929);
   U1019 : INV_X1 port map( A => n13929, ZN => n3200);
   U1020 : OAI22_X1 port map( A1 => n11211, A2 => n14271, B1 => n10405, B2 => 
                           n14308, ZN => n13930);
   U1021 : INV_X1 port map( A => n13930, ZN => n2880);
   U1022 : OAI22_X1 port map( A1 => n11211, A2 => n14295, B1 => n10939, B2 => 
                           n14308, ZN => n13931);
   U1023 : INV_X1 port map( A => n13931, ZN => n3232);
   U1024 : OAI22_X1 port map( A1 => n11211, A2 => n14337, B1 => n10559, B2 => 
                           n14308, ZN => n13932);
   U1025 : INV_X1 port map( A => n13932, ZN => n2848);
   U1026 : OAI22_X1 port map( A1 => n11211, A2 => n14267, B1 => n10467, B2 => 
                           n14308, ZN => n13933);
   U1027 : INV_X1 port map( A => n13933, ZN => n2786);
   U1028 : OAI22_X1 port map( A1 => n11211, A2 => n14241, B1 => n10313, B2 => 
                           n14308, ZN => n13934);
   U1029 : INV_X1 port map( A => n13934, ZN => n2722);
   U1030 : OAI22_X1 port map( A1 => n10091, A2 => n14285, B1 => n10496, B2 => 
                           n14308, ZN => n13935);
   U1031 : INV_X1 port map( A => n13935, ZN => n3040);
   U1032 : OAI22_X1 port map( A1 => n10091, A2 => n14280, B1 => n10849, B2 => 
                           n14308, ZN => n13936);
   U1033 : INV_X1 port map( A => n13936, ZN => n3136);
   U1034 : OAI22_X1 port map( A1 => n10091, A2 => n14276, B1 => n10610, B2 => 
                           n14308, ZN => n13937);
   U1035 : INV_X1 port map( A => n13937, ZN => n2976);
   U1036 : OAI22_X1 port map( A1 => n11211, A2 => n14375, B1 => n10287, B2 => 
                           n14308, ZN => n13938);
   U1037 : INV_X1 port map( A => n13938, ZN => n2658);
   U1038 : OAI22_X1 port map( A1 => n10091, A2 => n14220, B1 => n10999, B2 => 
                           n14308, ZN => n13939);
   U1039 : INV_X1 port map( A => n13939, ZN => n3296);
   U1040 : OAI22_X1 port map( A1 => n11211, A2 => n14334, B1 => n10589, B2 => 
                           n14308, ZN => n13940);
   U1041 : INV_X1 port map( A => n13940, ZN => n2816);
   U1042 : OAI22_X1 port map( A1 => n11211, A2 => n14218, B1 => n10969, B2 => 
                           n14308, ZN => n13941);
   U1043 : INV_X1 port map( A => n13941, ZN => n3264);
   U1044 : OAI22_X1 port map( A1 => n11211, A2 => n14163, B1 => n10128, B2 => 
                           n14308, ZN => n13942);
   U1045 : INV_X1 port map( A => n13942, ZN => n2568);
   U1046 : OAI22_X1 port map( A1 => n10091, A2 => n14282, B1 => n10790, B2 => 
                           n14308, ZN => n13943);
   U1047 : INV_X1 port map( A => n13943, ZN => n3104);
   U1048 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11203, ZN => n14417);
   U1049 : OAI22_X1 port map( A1 => n10082, A2 => n14282, B1 => n10777, B2 => 
                           n14417, ZN => n13944);
   U1050 : INV_X1 port map( A => n13944, ZN => n3113);
   U1051 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11202, ZN => n14466);
   U1052 : OAI22_X1 port map( A1 => n10081, A2 => n14488, B1 => n10657, B2 => 
                           n14466, ZN => n13945);
   U1053 : INV_X1 port map( A => n13945, ZN => n2922);
   U1054 : OAI22_X1 port map( A1 => n10082, A2 => n14488, B1 => n10656, B2 => 
                           n14417, ZN => n13946);
   U1055 : INV_X1 port map( A => n13946, ZN => n2921);
   U1056 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11204, ZN => n14458);
   U1057 : OAI22_X1 port map( A1 => n10083, A2 => n14282, B1 => n10776, B2 => 
                           n14458, ZN => n13947);
   U1058 : INV_X1 port map( A => n13947, ZN => n3112);
   U1059 : OAI22_X1 port map( A1 => n10081, A2 => n14274, B1 => n10627, B2 => 
                           n14466, ZN => n13948);
   U1060 : INV_X1 port map( A => n13948, ZN => n2954);
   U1061 : OAI22_X1 port map( A1 => n10082, A2 => n14274, B1 => n10626, B2 => 
                           n14417, ZN => n13949);
   U1062 : INV_X1 port map( A => n13949, ZN => n2953);
   U1063 : OAI22_X1 port map( A1 => n10083, A2 => n14274, B1 => n10625, B2 => 
                           n14458, ZN => n13950);
   U1064 : INV_X1 port map( A => n13950, ZN => n2952);
   U1065 : OAI22_X1 port map( A1 => n10083, A2 => n14488, B1 => n10655, B2 => 
                           n14458, ZN => n13951);
   U1066 : INV_X1 port map( A => n13951, ZN => n2920);
   U1067 : OAI22_X1 port map( A1 => n11202, A2 => n14334, B1 => n10599, B2 => 
                           n14466, ZN => n13952);
   U1068 : INV_X1 port map( A => n13952, ZN => n2826);
   U1069 : OAI22_X1 port map( A1 => n11203, A2 => n14334, B1 => n10598, B2 => 
                           n14417, ZN => n13953);
   U1070 : INV_X1 port map( A => n13953, ZN => n2825);
   U1071 : OAI22_X1 port map( A1 => n11204, A2 => n14334, B1 => n10597, B2 => 
                           n14458, ZN => n13954);
   U1072 : INV_X1 port map( A => n13954, ZN => n2824);
   U1073 : OAI22_X1 port map( A1 => n11203, A2 => n14337, B1 => n10568, B2 => 
                           n14417, ZN => n13955);
   U1074 : INV_X1 port map( A => n13955, ZN => n2857);
   U1075 : OAI22_X1 port map( A1 => n11204, A2 => n14337, B1 => n10567, B2 => 
                           n14458, ZN => n13956);
   U1076 : INV_X1 port map( A => n13956, ZN => n2856);
   U1077 : OAI22_X1 port map( A1 => n11202, A2 => n14337, B1 => n10547, B2 => 
                           n14466, ZN => n13957);
   U1078 : INV_X1 port map( A => n13957, ZN => n2858);
   U1079 : OAI22_X1 port map( A1 => n10082, A2 => n14276, B1 => n10535, B2 => 
                           n14417, ZN => n13958);
   U1080 : INV_X1 port map( A => n13958, ZN => n2985);
   U1081 : OAI22_X1 port map( A1 => n10083, A2 => n14276, B1 => n10534, B2 => 
                           n14458, ZN => n13959);
   U1082 : INV_X1 port map( A => n13959, ZN => n2984);
   U1083 : OAI22_X1 port map( A1 => n10081, A2 => n14276, B1 => n10536, B2 => 
                           n14466, ZN => n13960);
   U1084 : INV_X1 port map( A => n13960, ZN => n2986);
   U1085 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11199, ZN => n14474);
   U1086 : OAI22_X1 port map( A1 => n10077, A2 => n14282, B1 => n10761, B2 => 
                           n14474, ZN => n13961);
   U1087 : INV_X1 port map( A => n13961, ZN => n3118);
   U1088 : OAI22_X1 port map( A1 => n10077, A2 => n14276, B1 => n10520, B2 => 
                           n14474, ZN => n13962);
   U1089 : INV_X1 port map( A => n13962, ZN => n2990);
   U1090 : OAI22_X1 port map( A1 => n10077, A2 => n14274, B1 => n10612, B2 => 
                           n14474, ZN => n13963);
   U1091 : INV_X1 port map( A => n13963, ZN => n2958);
   U1092 : OAI22_X1 port map( A1 => n10077, A2 => n14488, B1 => n10641, B2 => 
                           n14474, ZN => n13964);
   U1093 : INV_X1 port map( A => n13964, ZN => n2926);
   U1094 : OAI22_X1 port map( A1 => n11199, A2 => n14337, B1 => n10551, B2 => 
                           n14474, ZN => n13965);
   U1095 : INV_X1 port map( A => n13965, ZN => n2862);
   U1096 : OAI22_X1 port map( A1 => n11199, A2 => n14334, B1 => n10582, B2 => 
                           n14474, ZN => n13966);
   U1097 : INV_X1 port map( A => n13966, ZN => n2830);
   U1098 : OAI22_X1 port map( A1 => n11203, A2 => n14253, B1 => n11123, B2 => 
                           n14417, ZN => n13967);
   U1099 : INV_X1 port map( A => n13967, ZN => n2773);
   U1100 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11200, ZN => n14476);
   U1101 : OAI22_X1 port map( A1 => n10078, A2 => n14282, B1 => n10781, B2 => 
                           n14476, ZN => n13968);
   U1102 : INV_X1 port map( A => n13968, ZN => n3117);
   U1103 : OAI22_X1 port map( A1 => n10078, A2 => n14276, B1 => n10519, B2 => 
                           n14476, ZN => n13969);
   U1104 : INV_X1 port map( A => n13969, ZN => n2989);
   U1105 : OAI22_X1 port map( A1 => n10078, A2 => n14274, B1 => n10611, B2 => 
                           n14476, ZN => n13970);
   U1106 : INV_X1 port map( A => n13970, ZN => n2957);
   U1107 : OAI22_X1 port map( A1 => n10078, A2 => n14488, B1 => n10660, B2 => 
                           n14476, ZN => n13971);
   U1108 : INV_X1 port map( A => n13971, ZN => n2925);
   U1109 : OAI22_X1 port map( A1 => n11200, A2 => n14337, B1 => n10550, B2 => 
                           n14476, ZN => n13972);
   U1110 : INV_X1 port map( A => n13972, ZN => n2861);
   U1111 : OAI22_X1 port map( A1 => n11200, A2 => n14334, B1 => n10581, B2 => 
                           n14476, ZN => n13973);
   U1112 : INV_X1 port map( A => n13973, ZN => n2829);
   U1113 : OAI22_X1 port map( A1 => n10082, A2 => n14220, B1 => n11008, B2 => 
                           n14417, ZN => n13974);
   U1114 : INV_X1 port map( A => n13974, ZN => n3305);
   U1115 : OAI22_X1 port map( A1 => n10083, A2 => n14220, B1 => n11007, B2 => 
                           n14458, ZN => n13975);
   U1116 : INV_X1 port map( A => n13975, ZN => n3304);
   U1117 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11205, ZN => n14470);
   U1118 : OAI22_X1 port map( A1 => n10084, A2 => n14220, B1 => n11006, B2 => 
                           n14470, ZN => n13976);
   U1119 : INV_X1 port map( A => n13976, ZN => n3303);
   U1120 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11201, ZN => n14460);
   U1121 : OAI22_X1 port map( A1 => n10079, A2 => n14282, B1 => n10780, B2 => 
                           n14460, ZN => n13977);
   U1122 : INV_X1 port map( A => n13977, ZN => n3116);
   U1123 : OAI22_X1 port map( A1 => n10077, A2 => n14220, B1 => n10991, B2 => 
                           n14474, ZN => n13978);
   U1124 : INV_X1 port map( A => n13978, ZN => n3310);
   U1125 : OAI22_X1 port map( A1 => n10078, A2 => n14220, B1 => n10990, B2 => 
                           n14476, ZN => n13979);
   U1126 : INV_X1 port map( A => n13979, ZN => n3309);
   U1127 : OAI22_X1 port map( A1 => n10079, A2 => n14220, B1 => n10989, B2 => 
                           n14460, ZN => n13980);
   U1128 : INV_X1 port map( A => n13980, ZN => n3308);
   U1129 : OAI22_X1 port map( A1 => n10079, A2 => n14276, B1 => n10518, B2 => 
                           n14460, ZN => n13981);
   U1130 : INV_X1 port map( A => n13981, ZN => n2988);
   U1131 : OAI22_X1 port map( A1 => n10079, A2 => n14274, B1 => n10629, B2 => 
                           n14460, ZN => n13982);
   U1132 : INV_X1 port map( A => n13982, ZN => n2956);
   U1133 : OAI22_X1 port map( A1 => n10079, A2 => n14488, B1 => n10659, B2 => 
                           n14460, ZN => n13983);
   U1134 : INV_X1 port map( A => n13983, ZN => n2924);
   U1135 : OAI22_X1 port map( A1 => n11201, A2 => n14337, B1 => n10549, B2 => 
                           n14460, ZN => n13984);
   U1136 : INV_X1 port map( A => n13984, ZN => n2860);
   U1137 : OAI22_X1 port map( A1 => n11201, A2 => n14334, B1 => n10580, B2 => 
                           n14460, ZN => n13985);
   U1138 : INV_X1 port map( A => n13985, ZN => n2828);
   U1139 : OAI22_X1 port map( A1 => n11204, A2 => n14218, B1 => n10977, B2 => 
                           n14458, ZN => n13986);
   U1140 : INV_X1 port map( A => n13986, ZN => n3272);
   U1141 : OAI22_X1 port map( A1 => n11205, A2 => n14218, B1 => n10976, B2 => 
                           n14470, ZN => n13987);
   U1142 : INV_X1 port map( A => n13987, ZN => n3271);
   U1143 : OAI22_X1 port map( A1 => n11200, A2 => n14218, B1 => n10960, B2 => 
                           n14476, ZN => n13988);
   U1144 : INV_X1 port map( A => n13988, ZN => n3277);
   U1145 : OAI22_X1 port map( A1 => n11201, A2 => n14218, B1 => n10959, B2 => 
                           n14460, ZN => n13989);
   U1146 : INV_X1 port map( A => n13989, ZN => n3276);
   U1147 : OAI22_X1 port map( A1 => n11203, A2 => n14125, B1 => n10956, B2 => 
                           n14417, ZN => n13990);
   U1148 : INV_X1 port map( A => n13990, ZN => n3273);
   U1149 : OAI22_X1 port map( A1 => n11205, A2 => n14295, B1 => n10946, B2 => 
                           n14470, ZN => n13991);
   U1150 : INV_X1 port map( A => n13991, ZN => n3239);
   U1151 : OAI22_X1 port map( A1 => n10083, A2 => n14484, B1 => n10805, B2 => 
                           n14458, ZN => n13992);
   U1152 : INV_X1 port map( A => n13992, ZN => n3080);
   U1153 : OAI22_X1 port map( A1 => n10082, A2 => n14484, B1 => n10806, B2 => 
                           n14417, ZN => n13993);
   U1154 : INV_X1 port map( A => n13993, ZN => n3081);
   U1155 : OAI22_X1 port map( A1 => n10079, A2 => n14484, B1 => n10809, B2 => 
                           n14460, ZN => n13994);
   U1156 : INV_X1 port map( A => n13994, ZN => n3084);
   U1157 : OAI22_X1 port map( A1 => n10078, A2 => n14484, B1 => n10810, B2 => 
                           n14476, ZN => n13995);
   U1158 : INV_X1 port map( A => n13995, ZN => n3085);
   U1159 : OAI22_X1 port map( A1 => n10077, A2 => n14484, B1 => n10811, B2 => 
                           n14474, ZN => n13996);
   U1160 : INV_X1 port map( A => n13996, ZN => n3086);
   U1161 : OAI22_X1 port map( A1 => n10081, A2 => n14484, B1 => n10807, B2 => 
                           n14466, ZN => n13997);
   U1162 : INV_X1 port map( A => n13997, ZN => n3082);
   U1163 : OAI22_X1 port map( A1 => n10081, A2 => n14282, B1 => n10778, B2 => 
                           n14466, ZN => n13998);
   U1164 : INV_X1 port map( A => n13998, ZN => n3114);
   U1165 : OAI22_X1 port map( A1 => n11202, A2 => n14218, B1 => n10957, B2 => 
                           n14466, ZN => n13999);
   U1166 : INV_X1 port map( A => n13999, ZN => n3274);
   U1167 : OAI22_X1 port map( A1 => n10081, A2 => n14220, B1 => n10987, B2 => 
                           n14466, ZN => n14000);
   U1168 : INV_X1 port map( A => n14000, ZN => n3306);
   U1169 : OAI22_X1 port map( A1 => n10083, A2 => n14280, B1 => n10835, B2 => 
                           n14458, ZN => n14001);
   U1170 : INV_X1 port map( A => n14001, ZN => n3144);
   U1171 : OAI22_X1 port map( A1 => n10082, A2 => n14280, B1 => n10836, B2 => 
                           n14417, ZN => n14002);
   U1172 : INV_X1 port map( A => n14002, ZN => n3145);
   U1173 : OAI22_X1 port map( A1 => n10081, A2 => n14280, B1 => n10837, B2 => 
                           n14466, ZN => n14003);
   U1174 : INV_X1 port map( A => n14003, ZN => n3146);
   U1175 : OAI22_X1 port map( A1 => n10079, A2 => n14280, B1 => n10839, B2 => 
                           n14460, ZN => n14004);
   U1176 : INV_X1 port map( A => n14004, ZN => n3148);
   U1177 : OAI22_X1 port map( A1 => n10078, A2 => n14280, B1 => n10840, B2 => 
                           n14476, ZN => n14005);
   U1178 : INV_X1 port map( A => n14005, ZN => n3149);
   U1179 : OAI22_X1 port map( A1 => n10077, A2 => n14280, B1 => n10841, B2 => 
                           n14474, ZN => n14006);
   U1180 : INV_X1 port map( A => n14006, ZN => n3150);
   U1181 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11224, ZN => n14478);
   U1182 : OAI22_X1 port map( A1 => n11224, A2 => n14334, B1 => n10579, B2 => 
                           n14478, ZN => n14007);
   U1183 : INV_X1 port map( A => n14007, ZN => n2827);
   U1184 : OAI22_X1 port map( A1 => n10083, A2 => n14287, B1 => n10865, B2 => 
                           n14458, ZN => n14008);
   U1185 : INV_X1 port map( A => n14008, ZN => n3176);
   U1186 : OAI22_X1 port map( A1 => n10082, A2 => n14287, B1 => n10866, B2 => 
                           n14417, ZN => n14009);
   U1187 : INV_X1 port map( A => n14009, ZN => n3177);
   U1188 : OAI22_X1 port map( A1 => n10081, A2 => n14287, B1 => n10867, B2 => 
                           n14466, ZN => n14010);
   U1189 : INV_X1 port map( A => n14010, ZN => n3178);
   U1190 : OAI22_X1 port map( A1 => n10079, A2 => n14287, B1 => n10869, B2 => 
                           n14460, ZN => n14011);
   U1191 : INV_X1 port map( A => n14011, ZN => n3180);
   U1192 : OAI22_X1 port map( A1 => n10078, A2 => n14287, B1 => n10870, B2 => 
                           n14476, ZN => n14012);
   U1193 : INV_X1 port map( A => n14012, ZN => n3181);
   U1194 : OAI22_X1 port map( A1 => n10077, A2 => n14287, B1 => n10871, B2 => 
                           n14474, ZN => n14013);
   U1195 : INV_X1 port map( A => n14013, ZN => n3182);
   U1196 : OAI22_X1 port map( A1 => n11224, A2 => n14337, B1 => n10548, B2 => 
                           n14478, ZN => n14014);
   U1197 : INV_X1 port map( A => n14014, ZN => n2859);
   U1198 : OAI22_X1 port map( A1 => n10080, A2 => n14488, B1 => n10658, B2 => 
                           n14478, ZN => n14015);
   U1199 : INV_X1 port map( A => n14015, ZN => n2923);
   U1200 : OAI22_X1 port map( A1 => n10080, A2 => n14274, B1 => n10628, B2 => 
                           n14478, ZN => n14016);
   U1201 : INV_X1 port map( A => n14016, ZN => n2955);
   U1202 : OAI22_X1 port map( A1 => n10080, A2 => n14276, B1 => n10537, B2 => 
                           n14478, ZN => n14017);
   U1203 : INV_X1 port map( A => n14017, ZN => n2987);
   U1204 : OAI22_X1 port map( A1 => n10080, A2 => n14484, B1 => n10808, B2 => 
                           n14478, ZN => n14018);
   U1205 : INV_X1 port map( A => n14018, ZN => n3083);
   U1206 : OAI22_X1 port map( A1 => n10080, A2 => n14282, B1 => n10779, B2 => 
                           n14478, ZN => n14019);
   U1207 : INV_X1 port map( A => n14019, ZN => n3115);
   U1208 : OAI22_X1 port map( A1 => n10080, A2 => n14280, B1 => n10838, B2 => 
                           n14478, ZN => n14020);
   U1209 : INV_X1 port map( A => n14020, ZN => n3147);
   U1210 : OAI22_X1 port map( A1 => n10080, A2 => n14287, B1 => n10868, B2 => 
                           n14478, ZN => n14021);
   U1211 : INV_X1 port map( A => n14021, ZN => n3179);
   U1212 : OAI22_X1 port map( A1 => n11204, A2 => n14210, B1 => n10895, B2 => 
                           n14458, ZN => n14022);
   U1213 : INV_X1 port map( A => n14022, ZN => n3208);
   U1214 : OAI22_X1 port map( A1 => n11203, A2 => n14210, B1 => n10896, B2 => 
                           n14417, ZN => n14023);
   U1215 : INV_X1 port map( A => n14023, ZN => n3209);
   U1216 : OAI22_X1 port map( A1 => n11202, A2 => n14210, B1 => n10897, B2 => 
                           n14466, ZN => n14024);
   U1217 : INV_X1 port map( A => n14024, ZN => n3210);
   U1218 : OAI22_X1 port map( A1 => n11224, A2 => n14210, B1 => n10898, B2 => 
                           n14478, ZN => n14025);
   U1219 : INV_X1 port map( A => n14025, ZN => n3211);
   U1220 : OAI22_X1 port map( A1 => n11201, A2 => n14210, B1 => n10899, B2 => 
                           n14460, ZN => n14026);
   U1221 : INV_X1 port map( A => n14026, ZN => n3212);
   U1222 : OAI22_X1 port map( A1 => n11200, A2 => n14210, B1 => n10900, B2 => 
                           n14476, ZN => n14027);
   U1223 : INV_X1 port map( A => n14027, ZN => n3213);
   U1224 : OAI22_X1 port map( A1 => n11199, A2 => n14210, B1 => n10901, B2 => 
                           n14474, ZN => n14028);
   U1225 : INV_X1 port map( A => n14028, ZN => n3214);
   U1226 : OAI22_X1 port map( A1 => n11224, A2 => n14218, B1 => n10958, B2 => 
                           n14478, ZN => n14029);
   U1227 : INV_X1 port map( A => n14029, ZN => n3275);
   U1228 : OAI22_X1 port map( A1 => n10080, A2 => n14220, B1 => n10988, B2 => 
                           n14478, ZN => n14030);
   U1229 : INV_X1 port map( A => n14030, ZN => n3307);
   U1230 : OAI22_X1 port map( A1 => n11204, A2 => n14295, B1 => n10925, B2 => 
                           n14458, ZN => n14031);
   U1231 : INV_X1 port map( A => n14031, ZN => n3240);
   U1232 : OAI22_X1 port map( A1 => n11202, A2 => n14295, B1 => n10927, B2 => 
                           n14466, ZN => n14032);
   U1233 : INV_X1 port map( A => n14032, ZN => n3242);
   U1234 : OAI22_X1 port map( A1 => n11224, A2 => n14295, B1 => n10928, B2 => 
                           n14478, ZN => n14033);
   U1235 : INV_X1 port map( A => n14033, ZN => n3243);
   U1236 : OAI22_X1 port map( A1 => n11201, A2 => n14295, B1 => n10929, B2 => 
                           n14460, ZN => n14034);
   U1237 : INV_X1 port map( A => n14034, ZN => n3244);
   U1238 : OAI22_X1 port map( A1 => n11200, A2 => n14295, B1 => n10930, B2 => 
                           n14476, ZN => n14035);
   U1239 : INV_X1 port map( A => n14035, ZN => n3245);
   U1240 : OAI22_X1 port map( A1 => n11199, A2 => n14295, B1 => n10931, B2 => 
                           n14474, ZN => n14036);
   U1241 : INV_X1 port map( A => n14036, ZN => n3246);
   U1242 : OAI22_X1 port map( A1 => n11199, A2 => n14218, B1 => n10961, B2 => 
                           n14474, ZN => n14037);
   U1243 : INV_X1 port map( A => n14037, ZN => n3278);
   U1244 : OAI22_X1 port map( A1 => n11199, A2 => n14344, B1 => n10365, B2 => 
                           n14474, ZN => n14038);
   U1245 : INV_X1 port map( A => n14038, ZN => n2766);
   U1246 : OAI22_X1 port map( A1 => n11201, A2 => n14344, B1 => n10363, B2 => 
                           n14460, ZN => n14039);
   U1247 : INV_X1 port map( A => n14039, ZN => n2764);
   U1248 : OAI22_X1 port map( A1 => n11224, A2 => n14344, B1 => n10362, B2 => 
                           n14478, ZN => n14040);
   U1249 : INV_X1 port map( A => n14040, ZN => n2763);
   U1250 : OAI22_X1 port map( A1 => n11202, A2 => n14344, B1 => n10361, B2 => 
                           n14466, ZN => n14041);
   U1251 : INV_X1 port map( A => n14041, ZN => n2762);
   U1252 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11207, ZN => n14468);
   U1253 : OAI22_X1 port map( A1 => n10086, A2 => n14220, B1 => n11004, B2 => 
                           n14468, ZN => n14042);
   U1254 : INV_X1 port map( A => n14042, ZN => n3301);
   U1255 : OAI22_X1 port map( A1 => n11207, A2 => n14218, B1 => n10974, B2 => 
                           n14468, ZN => n14043);
   U1256 : INV_X1 port map( A => n14043, ZN => n3269);
   U1257 : OAI22_X1 port map( A1 => n11207, A2 => n14295, B1 => n10944, B2 => 
                           n14468, ZN => n14044);
   U1258 : INV_X1 port map( A => n14044, ZN => n3237);
   U1259 : OAI22_X1 port map( A1 => n11207, A2 => n14210, B1 => n10914, B2 => 
                           n14468, ZN => n14045);
   U1260 : INV_X1 port map( A => n14045, ZN => n3205);
   U1261 : OAI22_X1 port map( A1 => n10086, A2 => n14287, B1 => n10884, B2 => 
                           n14468, ZN => n14046);
   U1262 : INV_X1 port map( A => n14046, ZN => n3173);
   U1263 : OAI22_X1 port map( A1 => n10086, A2 => n14280, B1 => n10832, B2 => 
                           n14468, ZN => n14047);
   U1264 : INV_X1 port map( A => n14047, ZN => n3141);
   U1265 : OAI22_X1 port map( A1 => n10086, A2 => n14282, B1 => n10773, B2 => 
                           n14468, ZN => n14048);
   U1266 : INV_X1 port map( A => n14048, ZN => n3109);
   U1267 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11210, ZN => n14464);
   U1268 : OAI22_X1 port map( A1 => n11210, A2 => n14241, B1 => n10314, B2 => 
                           n14464, ZN => n14049);
   U1269 : INV_X1 port map( A => n14049, ZN => n2723);
   U1270 : OAI22_X1 port map( A1 => n10086, A2 => n14484, B1 => n10802, B2 => 
                           n14468, ZN => n14050);
   U1271 : INV_X1 port map( A => n14050, ZN => n3077);
   U1272 : OAI22_X1 port map( A1 => n10086, A2 => n14276, B1 => n10531, B2 => 
                           n14468, ZN => n14051);
   U1273 : INV_X1 port map( A => n14051, ZN => n2981);
   U1274 : OAI22_X1 port map( A1 => n11199, A2 => n14241, B1 => n10305, B2 => 
                           n14474, ZN => n14052);
   U1275 : INV_X1 port map( A => n14052, ZN => n2734);
   U1276 : OAI22_X1 port map( A1 => n11200, A2 => n14093, B1 => n10304, B2 => 
                           n14476, ZN => n14053);
   U1277 : INV_X1 port map( A => n14053, ZN => n2733);
   U1278 : OAI22_X1 port map( A1 => n11201, A2 => n14241, B1 => n10303, B2 => 
                           n14460, ZN => n14054);
   U1279 : INV_X1 port map( A => n14054, ZN => n2732);
   U1280 : OAI22_X1 port map( A1 => n11224, A2 => n14241, B1 => n10302, B2 => 
                           n14478, ZN => n14055);
   U1281 : INV_X1 port map( A => n14055, ZN => n2731);
   U1282 : OAI22_X1 port map( A1 => n11202, A2 => n14241, B1 => n10301, B2 => 
                           n14466, ZN => n14056);
   U1283 : INV_X1 port map( A => n14056, ZN => n2730);
   U1284 : OAI22_X1 port map( A1 => n11203, A2 => n14093, B1 => n10300, B2 => 
                           n14417, ZN => n14057);
   U1285 : INV_X1 port map( A => n14057, ZN => n2709);
   U1286 : OAI22_X1 port map( A1 => n11204, A2 => n14241, B1 => n10299, B2 => 
                           n14458, ZN => n14058);
   U1287 : INV_X1 port map( A => n14058, ZN => n2729);
   U1288 : OAI22_X1 port map( A1 => n11210, A2 => n14334, B1 => n10590, B2 => 
                           n14464, ZN => n14059);
   U1289 : INV_X1 port map( A => n14059, ZN => n2817);
   U1290 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11206, ZN => n14353);
   U1291 : OAI22_X1 port map( A1 => n11206, A2 => n14241, B1 => n10297, B2 => 
                           n14353, ZN => n14060);
   U1292 : INV_X1 port map( A => n14060, ZN => n2727);
   U1293 : OAI22_X1 port map( A1 => n10086, A2 => n14274, B1 => n10622, B2 => 
                           n14468, ZN => n14061);
   U1294 : INV_X1 port map( A => n14061, ZN => n2949);
   U1295 : OAI22_X1 port map( A1 => n10086, A2 => n14488, B1 => n10652, B2 => 
                           n14468, ZN => n14062);
   U1296 : INV_X1 port map( A => n14062, ZN => n2917);
   U1297 : OAI22_X1 port map( A1 => n11207, A2 => n14337, B1 => n10564, B2 => 
                           n14468, ZN => n14063);
   U1298 : INV_X1 port map( A => n14063, ZN => n2853);
   U1299 : OAI22_X1 port map( A1 => n11207, A2 => n14334, B1 => n10594, B2 => 
                           n14468, ZN => n14064);
   U1300 : INV_X1 port map( A => n14064, ZN => n2821);
   U1301 : OAI22_X1 port map( A1 => n11210, A2 => n14337, B1 => n10560, B2 => 
                           n14464, ZN => n14065);
   U1302 : INV_X1 port map( A => n14065, ZN => n2849);
   U1303 : OAI22_X1 port map( A1 => n10090, A2 => n14488, B1 => n10759, B2 => 
                           n14464, ZN => n14066);
   U1304 : INV_X1 port map( A => n14066, ZN => n2913);
   U1305 : OAI22_X1 port map( A1 => n10090, A2 => n14274, B1 => n10640, B2 => 
                           n14464, ZN => n14067);
   U1306 : INV_X1 port map( A => n14067, ZN => n2945);
   U1307 : OAI22_X1 port map( A1 => n11207, A2 => n14241, B1 => n10318, B2 => 
                           n14468, ZN => n14068);
   U1308 : INV_X1 port map( A => n14068, ZN => n2726);
   U1309 : OAI22_X1 port map( A1 => n10090, A2 => n14276, B1 => n10527, B2 => 
                           n14464, ZN => n14069);
   U1310 : INV_X1 port map( A => n14069, ZN => n2977);
   U1311 : OAI22_X1 port map( A1 => n10090, A2 => n14484, B1 => n10820, B2 => 
                           n14464, ZN => n14070);
   U1312 : INV_X1 port map( A => n14070, ZN => n3073);
   U1313 : OAI22_X1 port map( A1 => n11224, A2 => n14375, B1 => n10276, B2 => 
                           n14478, ZN => n14071);
   U1314 : INV_X1 port map( A => n14071, ZN => n2667);
   U1315 : OAI22_X1 port map( A1 => n11202, A2 => n14375, B1 => n10275, B2 => 
                           n14466, ZN => n14072);
   U1316 : INV_X1 port map( A => n14072, ZN => n2666);
   U1317 : OAI22_X1 port map( A1 => n10090, A2 => n14282, B1 => n10791, B2 => 
                           n14464, ZN => n14073);
   U1318 : INV_X1 port map( A => n14073, ZN => n3105);
   U1319 : OAI22_X1 port map( A1 => n10090, A2 => n14280, B1 => n10850, B2 => 
                           n14464, ZN => n14074);
   U1320 : INV_X1 port map( A => n14074, ZN => n3137);
   U1321 : OAI22_X1 port map( A1 => n10090, A2 => n14287, B1 => n10880, B2 => 
                           n14464, ZN => n14075);
   U1322 : INV_X1 port map( A => n14075, ZN => n3169);
   U1323 : OAI22_X1 port map( A1 => n11210, A2 => n14210, B1 => n10910, B2 => 
                           n14464, ZN => n14076);
   U1324 : INV_X1 port map( A => n14076, ZN => n3201);
   U1325 : OAI22_X1 port map( A1 => n11204, A2 => n14375, B1 => n10273, B2 => 
                           n14458, ZN => n14077);
   U1326 : INV_X1 port map( A => n14077, ZN => n2665);
   U1327 : OAI22_X1 port map( A1 => n11206, A2 => n14375, B1 => n10271, B2 => 
                           n14353, ZN => n14078);
   U1328 : INV_X1 port map( A => n14078, ZN => n2663);
   U1329 : OAI22_X1 port map( A1 => n11210, A2 => n14295, B1 => n10940, B2 => 
                           n14464, ZN => n14079);
   U1330 : INV_X1 port map( A => n14079, ZN => n3233);
   U1331 : OAI22_X1 port map( A1 => n11210, A2 => n14375, B1 => n10266, B2 => 
                           n14464, ZN => n14080);
   U1332 : INV_X1 port map( A => n14080, ZN => n2659);
   U1333 : OAI22_X1 port map( A1 => n11210, A2 => n14218, B1 => n10970, B2 => 
                           n14464, ZN => n14081);
   U1334 : INV_X1 port map( A => n14081, ZN => n3265);
   U1335 : OAI22_X1 port map( A1 => n11199, A2 => n14375, B1 => n10259, B2 => 
                           n14474, ZN => n14082);
   U1336 : INV_X1 port map( A => n14082, ZN => n2670);
   U1337 : OAI22_X1 port map( A1 => n10090, A2 => n14220, B1 => n11000, B2 => 
                           n14464, ZN => n14083);
   U1338 : INV_X1 port map( A => n14083, ZN => n3297);
   U1339 : OAI22_X1 port map( A1 => n11201, A2 => n14375, B1 => n10257, B2 => 
                           n14460, ZN => n14084);
   U1340 : INV_X1 port map( A => n14084, ZN => n2668);
   U1341 : OAI22_X1 port map( A1 => n11202, A2 => n14384, B1 => n10245, B2 => 
                           n14466, ZN => n14085);
   U1342 : INV_X1 port map( A => n14085, ZN => n2698);
   U1343 : OAI22_X1 port map( A1 => n11204, A2 => n14384, B1 => n10243, B2 => 
                           n14458, ZN => n14086);
   U1344 : INV_X1 port map( A => n14086, ZN => n2697);
   U1345 : OAI22_X1 port map( A1 => n11206, A2 => n14384, B1 => n10241, B2 => 
                           n14353, ZN => n14087);
   U1346 : INV_X1 port map( A => n14087, ZN => n2695);
   U1347 : OAI22_X1 port map( A1 => n11207, A2 => n14384, B1 => n10240, B2 => 
                           n14468, ZN => n14088);
   U1348 : INV_X1 port map( A => n14088, ZN => n2694);
   U1349 : OAI22_X1 port map( A1 => n11210, A2 => n14384, B1 => n10236, B2 => 
                           n14464, ZN => n14089);
   U1350 : INV_X1 port map( A => n14089, ZN => n2691);
   U1351 : OAI22_X1 port map( A1 => n11199, A2 => n14384, B1 => n10228, B2 => 
                           n14474, ZN => n14090);
   U1352 : INV_X1 port map( A => n14090, ZN => n2702);
   U1353 : OAI22_X1 port map( A1 => n11201, A2 => n14384, B1 => n10226, B2 => 
                           n14460, ZN => n14091);
   U1354 : INV_X1 port map( A => n14091, ZN => n2700);
   U1355 : OAI22_X1 port map( A1 => n11224, A2 => n14384, B1 => n10225, B2 => 
                           n14478, ZN => n14092);
   U1356 : INV_X1 port map( A => n14092, ZN => n2699);
   U1357 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11209, ZN => n14462);
   U1358 : OAI22_X1 port map( A1 => n11209, A2 => n14093, B1 => n10315, B2 => 
                           n14462, ZN => n14094);
   U1359 : INV_X1 port map( A => n14094, ZN => n2710);
   U1360 : OAI22_X1 port map( A1 => n11210, A2 => n14363, B1 => n10223, B2 => 
                           n14464, ZN => n14095);
   U1361 : INV_X1 port map( A => n14095, ZN => n2595);
   U1362 : OAI22_X1 port map( A1 => n11201, A2 => n14363, B1 => n10212, B2 => 
                           n14460, ZN => n14096);
   U1363 : INV_X1 port map( A => n14096, ZN => n2604);
   U1364 : OAI22_X1 port map( A1 => n11210, A2 => n14344, B1 => n10374, B2 => 
                           n14464, ZN => n14097);
   U1365 : INV_X1 port map( A => n14097, ZN => n2755);
   U1366 : OAI22_X1 port map( A1 => n11224, A2 => n14363, B1 => n10211, B2 => 
                           n14478, ZN => n14098);
   U1367 : INV_X1 port map( A => n14098, ZN => n2603);
   U1368 : OAI22_X1 port map( A1 => n11202, A2 => n14363, B1 => n10210, B2 => 
                           n14466, ZN => n14099);
   U1369 : INV_X1 port map( A => n14099, ZN => n2602);
   U1370 : OAI22_X1 port map( A1 => n11204, A2 => n14363, B1 => n10208, B2 => 
                           n14458, ZN => n14100);
   U1371 : INV_X1 port map( A => n14100, ZN => n2601);
   U1372 : OAI22_X1 port map( A1 => n11206, A2 => n14363, B1 => n10206, B2 => 
                           n14353, ZN => n14101);
   U1373 : INV_X1 port map( A => n14101, ZN => n2599);
   U1374 : OAI22_X1 port map( A1 => n11207, A2 => n14375, B1 => n10270, B2 => 
                           n14468, ZN => n14102);
   U1375 : INV_X1 port map( A => n14102, ZN => n2662);
   U1376 : OAI22_X1 port map( A1 => n11199, A2 => n14363, B1 => n10194, B2 => 
                           n14474, ZN => n14103);
   U1377 : INV_X1 port map( A => n14103, ZN => n2606);
   U1378 : OAI22_X1 port map( A1 => n11207, A2 => n14363, B1 => n10205, B2 => 
                           n14468, ZN => n14104);
   U1379 : INV_X1 port map( A => n14104, ZN => n2598);
   U1380 : OAI22_X1 port map( A1 => n10089, A2 => n14165, B1 => n10619, B2 => 
                           n14462, ZN => n14105);
   U1381 : INV_X1 port map( A => n14105, ZN => n2946);
   U1382 : OAI22_X1 port map( A1 => n10089, A2 => n14167, B1 => n10528, B2 => 
                           n14462, ZN => n14106);
   U1383 : INV_X1 port map( A => n14106, ZN => n2978);
   U1384 : OAI22_X1 port map( A1 => n10089, A2 => n14169, B1 => n10821, B2 => 
                           n14462, ZN => n14107);
   U1385 : INV_X1 port map( A => n14107, ZN => n3074);
   U1386 : OAI22_X1 port map( A1 => n11201, A2 => n14261, B1 => n10182, B2 => 
                           n14460, ZN => n14108);
   U1387 : INV_X1 port map( A => n14108, ZN => n2636);
   U1388 : OAI22_X1 port map( A1 => n11224, A2 => n14261, B1 => n10181, B2 => 
                           n14478, ZN => n14109);
   U1389 : INV_X1 port map( A => n14109, ZN => n2635);
   U1390 : OAI22_X1 port map( A1 => n11202, A2 => n14261, B1 => n10180, B2 => 
                           n14466, ZN => n14110);
   U1391 : INV_X1 port map( A => n14110, ZN => n2634);
   U1392 : OAI22_X1 port map( A1 => n11203, A2 => n14122, B1 => n10179, B2 => 
                           n14417, ZN => n14111);
   U1393 : INV_X1 port map( A => n14111, ZN => n2613);
   U1394 : OAI22_X1 port map( A1 => n11204, A2 => n14261, B1 => n10178, B2 => 
                           n14458, ZN => n14112);
   U1395 : INV_X1 port map( A => n14112, ZN => n2633);
   U1396 : OAI22_X1 port map( A1 => n11206, A2 => n14261, B1 => n10176, B2 => 
                           n14353, ZN => n14113);
   U1397 : INV_X1 port map( A => n14113, ZN => n2631);
   U1398 : OAI22_X1 port map( A1 => n10089, A2 => n14171, B1 => n10792, B2 => 
                           n14462, ZN => n14114);
   U1399 : INV_X1 port map( A => n14114, ZN => n3106);
   U1400 : OAI22_X1 port map( A1 => n11207, A2 => n14261, B1 => n10175, B2 => 
                           n14468, ZN => n14115);
   U1401 : INV_X1 port map( A => n14115, ZN => n2630);
   U1402 : OAI22_X1 port map( A1 => n11209, A2 => n14122, B1 => n10172, B2 => 
                           n14462, ZN => n14116);
   U1403 : INV_X1 port map( A => n14116, ZN => n2614);
   U1404 : OAI22_X1 port map( A1 => n10089, A2 => n14173, B1 => n10851, B2 => 
                           n14462, ZN => n14117);
   U1405 : INV_X1 port map( A => n14117, ZN => n3138);
   U1406 : OAI22_X1 port map( A1 => n10089, A2 => n14131, B1 => n10881, B2 => 
                           n14462, ZN => n14118);
   U1407 : INV_X1 port map( A => n14118, ZN => n3170);
   U1408 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11223, ZN => n14361);
   U1409 : OAI22_X1 port map( A1 => n10087, A2 => n14127, B1 => n11003, B2 => 
                           n14361, ZN => n14119);
   U1410 : INV_X1 port map( A => n14119, ZN => n3300);
   U1411 : OAI22_X1 port map( A1 => n11223, A2 => n14125, B1 => n10973, B2 => 
                           n14361, ZN => n14120);
   U1412 : INV_X1 port map( A => n14120, ZN => n3268);
   U1413 : OAI22_X1 port map( A1 => n11199, A2 => n14261, B1 => n10164, B2 => 
                           n14474, ZN => n14121);
   U1414 : INV_X1 port map( A => n14121, ZN => n2638);
   U1415 : OAI22_X1 port map( A1 => n11200, A2 => n14122, B1 => n10163, B2 => 
                           n14476, ZN => n14123);
   U1416 : INV_X1 port map( A => n14123, ZN => n2637);
   U1417 : OAI22_X1 port map( A1 => n11209, A2 => n14129, B1 => n10911, B2 => 
                           n14462, ZN => n14124);
   U1418 : INV_X1 port map( A => n14124, ZN => n3202);
   U1419 : OAI22_X1 port map( A1 => n11209, A2 => n14125, B1 => n10971, B2 => 
                           n14462, ZN => n14126);
   U1420 : INV_X1 port map( A => n14126, ZN => n3266);
   U1421 : OAI22_X1 port map( A1 => n10089, A2 => n14127, B1 => n11001, B2 => 
                           n14462, ZN => n14128);
   U1422 : INV_X1 port map( A => n14128, ZN => n3298);
   U1423 : OAI22_X1 port map( A1 => n11223, A2 => n14129, B1 => n10913, B2 => 
                           n14361, ZN => n14130);
   U1424 : INV_X1 port map( A => n14130, ZN => n3204);
   U1425 : OAI22_X1 port map( A1 => n10087, A2 => n14131, B1 => n10883, B2 => 
                           n14361, ZN => n14132);
   U1426 : INV_X1 port map( A => n14132, ZN => n3172);
   U1427 : OAI22_X1 port map( A1 => n10087, A2 => n14280, B1 => n10853, B2 => 
                           n14361, ZN => n14133);
   U1428 : INV_X1 port map( A => n14133, ZN => n3140);
   U1429 : NAND2_X1 port map( A1 => RESET_BAR, A2 => n11208, ZN => n14472);
   U1430 : OAI22_X1 port map( A1 => n11208, A2 => n14363, B1 => n10203, B2 => 
                           n14472, ZN => n14134);
   U1431 : INV_X1 port map( A => n14134, ZN => n2596);
   U1432 : OAI22_X1 port map( A1 => n11208, A2 => n14261, B1 => n10173, B2 => 
                           n14472, ZN => n14135);
   U1433 : INV_X1 port map( A => n14135, ZN => n2628);
   U1434 : OAI22_X1 port map( A1 => n11208, A2 => n14375, B1 => n10268, B2 => 
                           n14472, ZN => n14136);
   U1435 : INV_X1 port map( A => n14136, ZN => n2660);
   U1436 : OAI22_X1 port map( A1 => n11208, A2 => n14384, B1 => n10238, B2 => 
                           n14472, ZN => n14137);
   U1437 : INV_X1 port map( A => n14137, ZN => n2692);
   U1438 : OAI22_X1 port map( A1 => n11208, A2 => n14241, B1 => n10316, B2 => 
                           n14472, ZN => n14138);
   U1439 : INV_X1 port map( A => n14138, ZN => n2724);
   U1440 : OAI22_X1 port map( A1 => n10087, A2 => n14282, B1 => n10772, B2 => 
                           n14361, ZN => n14139);
   U1441 : INV_X1 port map( A => n14139, ZN => n3108);
   U1442 : OAI22_X1 port map( A1 => n10087, A2 => n14484, B1 => n10801, B2 => 
                           n14361, ZN => n14140);
   U1443 : INV_X1 port map( A => n14140, ZN => n3076);
   U1444 : OAI22_X1 port map( A1 => n10087, A2 => n14276, B1 => n10530, B2 => 
                           n14361, ZN => n14141);
   U1445 : INV_X1 port map( A => n14141, ZN => n2980);
   U1446 : OAI22_X1 port map( A1 => n10087, A2 => n14274, B1 => n10621, B2 => 
                           n14361, ZN => n14142);
   U1447 : INV_X1 port map( A => n14142, ZN => n2948);
   U1448 : OAI22_X1 port map( A1 => n10087, A2 => n14488, B1 => n10651, B2 => 
                           n14361, ZN => n14143);
   U1449 : INV_X1 port map( A => n14143, ZN => n2916);
   U1450 : OAI22_X1 port map( A1 => n11223, A2 => n14337, B1 => n10563, B2 => 
                           n14361, ZN => n14144);
   U1451 : INV_X1 port map( A => n14144, ZN => n2852);
   U1452 : OAI22_X1 port map( A1 => n11208, A2 => n14163, B1 => n10131, B2 => 
                           n14472, ZN => n14145);
   U1453 : INV_X1 port map( A => n14145, ZN => n2571);
   U1454 : OAI22_X1 port map( A1 => n11209, A2 => n14163, B1 => n10130, B2 => 
                           n14462, ZN => n14146);
   U1455 : INV_X1 port map( A => n14146, ZN => n2570);
   U1456 : OAI22_X1 port map( A1 => n11210, A2 => n14163, B1 => n10129, B2 => 
                           n14464, ZN => n14147);
   U1457 : INV_X1 port map( A => n14147, ZN => n2569);
   U1458 : OAI22_X1 port map( A1 => n11223, A2 => n14334, B1 => n10593, B2 => 
                           n14361, ZN => n14148);
   U1459 : INV_X1 port map( A => n14148, ZN => n2820);
   U1460 : OAI22_X1 port map( A1 => n11223, A2 => n14241, B1 => n10317, B2 => 
                           n14361, ZN => n14149);
   U1461 : INV_X1 port map( A => n14149, ZN => n2725);
   U1462 : OAI22_X1 port map( A1 => n11199, A2 => n14229, B1 => n10120, B2 => 
                           n14474, ZN => n14150);
   U1463 : INV_X1 port map( A => n14150, ZN => n2555);
   U1464 : OAI22_X1 port map( A1 => n11200, A2 => n14229, B1 => n10119, B2 => 
                           n14476, ZN => n14151);
   U1465 : INV_X1 port map( A => n14151, ZN => n2556);
   U1466 : OAI22_X1 port map( A1 => n11201, A2 => n14163, B1 => n10118, B2 => 
                           n14460, ZN => n14152);
   U1467 : INV_X1 port map( A => n14152, ZN => n2580);
   U1468 : OAI22_X1 port map( A1 => n11224, A2 => n14163, B1 => n10117, B2 => 
                           n14478, ZN => n14153);
   U1469 : INV_X1 port map( A => n14153, ZN => n2579);
   U1470 : OAI22_X1 port map( A1 => n11202, A2 => n14163, B1 => n10116, B2 => 
                           n14466, ZN => n14154);
   U1471 : INV_X1 port map( A => n14154, ZN => n2578);
   U1472 : OAI22_X1 port map( A1 => n11203, A2 => n14163, B1 => n10115, B2 => 
                           n14417, ZN => n14155);
   U1473 : INV_X1 port map( A => n14155, ZN => n2577);
   U1474 : OAI22_X1 port map( A1 => n11204, A2 => n14163, B1 => n10114, B2 => 
                           n14458, ZN => n14156);
   U1475 : INV_X1 port map( A => n14156, ZN => n2576);
   U1476 : OAI22_X1 port map( A1 => n11206, A2 => n14163, B1 => n10112, B2 => 
                           n14353, ZN => n14157);
   U1477 : INV_X1 port map( A => n14157, ZN => n2574);
   U1478 : OAI22_X1 port map( A1 => n11207, A2 => n14229, B1 => n10111, B2 => 
                           n14468, ZN => n14158);
   U1479 : INV_X1 port map( A => n14158, ZN => n2573);
   U1480 : OAI22_X1 port map( A1 => n11223, A2 => n14384, B1 => n10239, B2 => 
                           n14361, ZN => n14159);
   U1481 : INV_X1 port map( A => n14159, ZN => n2693);
   U1482 : OAI22_X1 port map( A1 => n11223, A2 => n14375, B1 => n10269, B2 => 
                           n14361, ZN => n14160);
   U1483 : INV_X1 port map( A => n14160, ZN => n2661);
   U1484 : OAI22_X1 port map( A1 => n11223, A2 => n14261, B1 => n10174, B2 => 
                           n14361, ZN => n14161);
   U1485 : INV_X1 port map( A => n14161, ZN => n2629);
   U1486 : OAI22_X1 port map( A1 => n11223, A2 => n14363, B1 => n10204, B2 => 
                           n14361, ZN => n14162);
   U1487 : INV_X1 port map( A => n14162, ZN => n2597);
   U1488 : OAI22_X1 port map( A1 => n11223, A2 => n14163, B1 => n10110, B2 => 
                           n14361, ZN => n14164);
   U1489 : INV_X1 port map( A => n14164, ZN => n2572);
   U1490 : OAI22_X1 port map( A1 => n10088, A2 => n14165, B1 => n10620, B2 => 
                           n14472, ZN => n14166);
   U1491 : INV_X1 port map( A => n14166, ZN => n2947);
   U1492 : OAI22_X1 port map( A1 => n10088, A2 => n14167, B1 => n10529, B2 => 
                           n14472, ZN => n14168);
   U1493 : INV_X1 port map( A => n14168, ZN => n2979);
   U1494 : OAI22_X1 port map( A1 => n10088, A2 => n14169, B1 => n10822, B2 => 
                           n14472, ZN => n14170);
   U1495 : INV_X1 port map( A => n14170, ZN => n3075);
   U1496 : OAI22_X1 port map( A1 => n10088, A2 => n14171, B1 => n10771, B2 => 
                           n14472, ZN => n14172);
   U1497 : INV_X1 port map( A => n14172, ZN => n3107);
   U1498 : OAI22_X1 port map( A1 => n10088, A2 => n14173, B1 => n10852, B2 => 
                           n14472, ZN => n14174);
   U1499 : INV_X1 port map( A => n14174, ZN => n3139);
   U1500 : OAI22_X1 port map( A1 => n10088, A2 => n14287, B1 => n10882, B2 => 
                           n14472, ZN => n14175);
   U1501 : INV_X1 port map( A => n14175, ZN => n3171);
   U1502 : OAI22_X1 port map( A1 => n11208, A2 => n14210, B1 => n10912, B2 => 
                           n14472, ZN => n14176);
   U1503 : INV_X1 port map( A => n14176, ZN => n3203);
   U1504 : OAI22_X1 port map( A1 => n10088, A2 => n14220, B1 => n11002, B2 => 
                           n14472, ZN => n14177);
   U1505 : INV_X1 port map( A => n14177, ZN => n3299);
   U1506 : OAI22_X1 port map( A1 => n11208, A2 => n14218, B1 => n10972, B2 => 
                           n14472, ZN => n14178);
   U1507 : INV_X1 port map( A => n14178, ZN => n3267);
   U1508 : OAI22_X1 port map( A1 => n11208, A2 => n14295, B1 => n10942, B2 => 
                           n14472, ZN => n14179);
   U1509 : INV_X1 port map( A => n14179, ZN => n3235);
   U1510 : OAI22_X1 port map( A1 => n11206, A2 => n14344, B1 => n10379, B2 => 
                           n14353, ZN => n14180);
   U1511 : INV_X1 port map( A => n14180, ZN => n2759);
   U1512 : OAI22_X1 port map( A1 => n11207, A2 => n14344, B1 => n10378, B2 => 
                           n14468, ZN => n14181);
   U1513 : INV_X1 port map( A => n14181, ZN => n2758);
   U1514 : OAI22_X1 port map( A1 => n11204, A2 => n14344, B1 => n10381, B2 => 
                           n14458, ZN => n14182);
   U1515 : INV_X1 port map( A => n14182, ZN => n2761);
   U1516 : OAI22_X1 port map( A1 => n11203, A2 => n14271, B1 => n10392, B2 => 
                           n14417, ZN => n14183);
   U1517 : INV_X1 port map( A => n14183, ZN => n2889);
   U1518 : OAI22_X1 port map( A1 => n11202, A2 => n14271, B1 => n10393, B2 => 
                           n14466, ZN => n14184);
   U1519 : INV_X1 port map( A => n14184, ZN => n2890);
   U1520 : OAI22_X1 port map( A1 => n11224, A2 => n14271, B1 => n10394, B2 => 
                           n14478, ZN => n14185);
   U1521 : INV_X1 port map( A => n14185, ZN => n2891);
   U1522 : OAI22_X1 port map( A1 => n11201, A2 => n14271, B1 => n10395, B2 => 
                           n14460, ZN => n14186);
   U1523 : INV_X1 port map( A => n14186, ZN => n2892);
   U1524 : OAI22_X1 port map( A1 => n11200, A2 => n14271, B1 => n10396, B2 => 
                           n14476, ZN => n14187);
   U1525 : INV_X1 port map( A => n14187, ZN => n2893);
   U1526 : OAI22_X1 port map( A1 => n11199, A2 => n14271, B1 => n10397, B2 => 
                           n14474, ZN => n14188);
   U1527 : INV_X1 port map( A => n14188, ZN => n2894);
   U1528 : OAI22_X1 port map( A1 => n11206, A2 => n14334, B1 => n10595, B2 => 
                           n14353, ZN => n14189);
   U1529 : INV_X1 port map( A => n14189, ZN => n2822);
   U1530 : OAI22_X1 port map( A1 => n11206, A2 => n14337, B1 => n10565, B2 => 
                           n14353, ZN => n14190);
   U1531 : INV_X1 port map( A => n14190, ZN => n2854);
   U1532 : OAI22_X1 port map( A1 => n10085, A2 => n14488, B1 => n10653, B2 => 
                           n14353, ZN => n14191);
   U1533 : INV_X1 port map( A => n14191, ZN => n2918);
   U1534 : OAI22_X1 port map( A1 => n10085, A2 => n14274, B1 => n10623, B2 => 
                           n14353, ZN => n14192);
   U1535 : INV_X1 port map( A => n14192, ZN => n2950);
   U1536 : OAI22_X1 port map( A1 => n11210, A2 => n14271, B1 => n10406, B2 => 
                           n14464, ZN => n14193);
   U1537 : INV_X1 port map( A => n14193, ZN => n2881);
   U1538 : OAI22_X1 port map( A1 => n11209, A2 => n14195, B1 => n10407, B2 => 
                           n14462, ZN => n14194);
   U1539 : INV_X1 port map( A => n14194, ZN => n2882);
   U1540 : OAI22_X1 port map( A1 => n11208, A2 => n14195, B1 => n10408, B2 => 
                           n14472, ZN => n14196);
   U1541 : INV_X1 port map( A => n14196, ZN => n2883);
   U1542 : OAI22_X1 port map( A1 => n11223, A2 => n14271, B1 => n10409, B2 => 
                           n14361, ZN => n14197);
   U1543 : INV_X1 port map( A => n14197, ZN => n2884);
   U1544 : OAI22_X1 port map( A1 => n11207, A2 => n14271, B1 => n10410, B2 => 
                           n14468, ZN => n14198);
   U1545 : INV_X1 port map( A => n14198, ZN => n2885);
   U1546 : OAI22_X1 port map( A1 => n11206, A2 => n14271, B1 => n10411, B2 => 
                           n14353, ZN => n14199);
   U1547 : INV_X1 port map( A => n14199, ZN => n2886);
   U1548 : OAI22_X1 port map( A1 => n11204, A2 => n14271, B1 => n10413, B2 => 
                           n14458, ZN => n14200);
   U1549 : INV_X1 port map( A => n14200, ZN => n2888);
   U1550 : OAI22_X1 port map( A1 => n10085, A2 => n14276, B1 => n10532, B2 => 
                           n14353, ZN => n14201);
   U1551 : INV_X1 port map( A => n14201, ZN => n2982);
   U1552 : OAI22_X1 port map( A1 => n10085, A2 => n14484, B1 => n10803, B2 => 
                           n14353, ZN => n14202);
   U1553 : INV_X1 port map( A => n14202, ZN => n3078);
   U1554 : OAI22_X1 port map( A1 => n10085, A2 => n14282, B1 => n10774, B2 => 
                           n14353, ZN => n14203);
   U1555 : INV_X1 port map( A => n14203, ZN => n3110);
   U1556 : OAI22_X1 port map( A1 => n11223, A2 => n14344, B1 => n10377, B2 => 
                           n14361, ZN => n14204);
   U1557 : INV_X1 port map( A => n14204, ZN => n2757);
   U1558 : OAI22_X1 port map( A1 => n10085, A2 => n14280, B1 => n10833, B2 => 
                           n14353, ZN => n14205);
   U1559 : INV_X1 port map( A => n14205, ZN => n3142);
   U1560 : OAI22_X1 port map( A1 => n10085, A2 => n14287, B1 => n10863, B2 => 
                           n14353, ZN => n14206);
   U1561 : INV_X1 port map( A => n14206, ZN => n3174);
   U1562 : OAI22_X1 port map( A1 => n11206, A2 => n14210, B1 => n10915, B2 => 
                           n14353, ZN => n14207);
   U1563 : INV_X1 port map( A => n14207, ZN => n3206);
   U1564 : OAI22_X1 port map( A1 => n11206, A2 => n14295, B1 => n10945, B2 => 
                           n14353, ZN => n14208);
   U1565 : INV_X1 port map( A => n14208, ZN => n3238);
   U1566 : OAI22_X1 port map( A1 => n10083, A2 => n14490, B1 => n10424, B2 => 
                           n14458, ZN => n14209);
   U1567 : INV_X1 port map( A => n14209, ZN => n3016);
   U1568 : OAI22_X1 port map( A1 => n11205, A2 => n14210, B1 => n10894, B2 => 
                           n14470, ZN => n14211);
   U1569 : INV_X1 port map( A => n14211, ZN => n3207);
   U1570 : OAI22_X1 port map( A1 => n10082, A2 => n14490, B1 => n10425, B2 => 
                           n14417, ZN => n14212);
   U1571 : INV_X1 port map( A => n14212, ZN => n3017);
   U1572 : OAI22_X1 port map( A1 => n10081, A2 => n14490, B1 => n10426, B2 => 
                           n14466, ZN => n14213);
   U1573 : INV_X1 port map( A => n14213, ZN => n3018);
   U1574 : OAI22_X1 port map( A1 => n10080, A2 => n14490, B1 => n10427, B2 => 
                           n14478, ZN => n14214);
   U1575 : INV_X1 port map( A => n14214, ZN => n3019);
   U1576 : OAI22_X1 port map( A1 => n10079, A2 => n14490, B1 => n10428, B2 => 
                           n14460, ZN => n14215);
   U1577 : INV_X1 port map( A => n14215, ZN => n3020);
   U1578 : OAI22_X1 port map( A1 => n10078, A2 => n14490, B1 => n10429, B2 => 
                           n14476, ZN => n14216);
   U1579 : INV_X1 port map( A => n14216, ZN => n3021);
   U1580 : OAI22_X1 port map( A1 => n10077, A2 => n14490, B1 => n10430, B2 => 
                           n14474, ZN => n14217);
   U1581 : INV_X1 port map( A => n14217, ZN => n3022);
   U1582 : OAI22_X1 port map( A1 => n11206, A2 => n14218, B1 => n10975, B2 => 
                           n14353, ZN => n14219);
   U1583 : INV_X1 port map( A => n14219, ZN => n3270);
   U1584 : OAI22_X1 port map( A1 => n10085, A2 => n14220, B1 => n11005, B2 => 
                           n14353, ZN => n14221);
   U1585 : INV_X1 port map( A => n14221, ZN => n3302);
   U1586 : OAI22_X1 port map( A1 => n10090, A2 => n14490, B1 => n10439, B2 => 
                           n14464, ZN => n14222);
   U1587 : INV_X1 port map( A => n14222, ZN => n3009);
   U1588 : OAI22_X1 port map( A1 => n10089, A2 => n14224, B1 => n10440, B2 => 
                           n14462, ZN => n14223);
   U1589 : INV_X1 port map( A => n14223, ZN => n3010);
   U1590 : OAI22_X1 port map( A1 => n10088, A2 => n14224, B1 => n10441, B2 => 
                           n14472, ZN => n14225);
   U1591 : INV_X1 port map( A => n14225, ZN => n3011);
   U1592 : OAI22_X1 port map( A1 => n10087, A2 => n14490, B1 => n10442, B2 => 
                           n14361, ZN => n14226);
   U1593 : INV_X1 port map( A => n14226, ZN => n3012);
   U1594 : OAI22_X1 port map( A1 => n10086, A2 => n14490, B1 => n10443, B2 => 
                           n14468, ZN => n14227);
   U1595 : INV_X1 port map( A => n14227, ZN => n3013);
   U1596 : OAI22_X1 port map( A1 => n10085, A2 => n14490, B1 => n10444, B2 => 
                           n14353, ZN => n14228);
   U1597 : INV_X1 port map( A => n14228, ZN => n3014);
   U1598 : OAI22_X1 port map( A1 => n11205, A2 => n14229, B1 => n10113, B2 => 
                           n14470, ZN => n14230);
   U1599 : INV_X1 port map( A => n14230, ZN => n2575);
   U1600 : OAI22_X1 port map( A1 => n11205, A2 => n14363, B1 => n10207, B2 => 
                           n14470, ZN => n14231);
   U1601 : INV_X1 port map( A => n14231, ZN => n2600);
   U1602 : OAI22_X1 port map( A1 => n11205, A2 => n14261, B1 => n10177, B2 => 
                           n14470, ZN => n14232);
   U1603 : INV_X1 port map( A => n14232, ZN => n2632);
   U1604 : OAI22_X1 port map( A1 => n11204, A2 => n14253, B1 => n10454, B2 => 
                           n14458, ZN => n14233);
   U1605 : INV_X1 port map( A => n14233, ZN => n2793);
   U1606 : OAI22_X1 port map( A1 => n11202, A2 => n14267, B1 => n10455, B2 => 
                           n14466, ZN => n14234);
   U1607 : INV_X1 port map( A => n14234, ZN => n2794);
   U1608 : OAI22_X1 port map( A1 => n11224, A2 => n14267, B1 => n10456, B2 => 
                           n14478, ZN => n14235);
   U1609 : INV_X1 port map( A => n14235, ZN => n2795);
   U1610 : OAI22_X1 port map( A1 => n11201, A2 => n14267, B1 => n10457, B2 => 
                           n14460, ZN => n14236);
   U1611 : INV_X1 port map( A => n14236, ZN => n2796);
   U1612 : OAI22_X1 port map( A1 => n11200, A2 => n14253, B1 => n10458, B2 => 
                           n14476, ZN => n14237);
   U1613 : INV_X1 port map( A => n14237, ZN => n2797);
   U1614 : OAI22_X1 port map( A1 => n11199, A2 => n14267, B1 => n10459, B2 => 
                           n14474, ZN => n14238);
   U1615 : INV_X1 port map( A => n14238, ZN => n2798);
   U1616 : OAI22_X1 port map( A1 => n11205, A2 => n14375, B1 => n10272, B2 => 
                           n14470, ZN => n14239);
   U1617 : INV_X1 port map( A => n14239, ZN => n2664);
   U1618 : OAI22_X1 port map( A1 => n11205, A2 => n14384, B1 => n10242, B2 => 
                           n14470, ZN => n14240);
   U1619 : INV_X1 port map( A => n14240, ZN => n2696);
   U1620 : OAI22_X1 port map( A1 => n11205, A2 => n14241, B1 => n10298, B2 => 
                           n14470, ZN => n14242);
   U1621 : INV_X1 port map( A => n14242, ZN => n2728);
   U1622 : OAI22_X1 port map( A1 => n11205, A2 => n14344, B1 => n10380, B2 => 
                           n14470, ZN => n14243);
   U1623 : INV_X1 port map( A => n14243, ZN => n2760);
   U1624 : OAI22_X1 port map( A1 => n11210, A2 => n14267, B1 => n10468, B2 => 
                           n14464, ZN => n14244);
   U1625 : INV_X1 port map( A => n14244, ZN => n2787);
   U1626 : OAI22_X1 port map( A1 => n10090, A2 => n14285, B1 => n10497, B2 => 
                           n14464, ZN => n14245);
   U1627 : INV_X1 port map( A => n14245, ZN => n3041);
   U1628 : OAI22_X1 port map( A1 => n10089, A2 => n14247, B1 => n10498, B2 => 
                           n14462, ZN => n14246);
   U1629 : INV_X1 port map( A => n14246, ZN => n3042);
   U1630 : OAI22_X1 port map( A1 => n10088, A2 => n14247, B1 => n10499, B2 => 
                           n14472, ZN => n14248);
   U1631 : INV_X1 port map( A => n14248, ZN => n3043);
   U1632 : OAI22_X1 port map( A1 => n10087, A2 => n14285, B1 => n10500, B2 => 
                           n14361, ZN => n14249);
   U1633 : INV_X1 port map( A => n14249, ZN => n3044);
   U1634 : OAI22_X1 port map( A1 => n10080, A2 => n14285, B1 => n10486, B2 => 
                           n14478, ZN => n14250);
   U1635 : INV_X1 port map( A => n14250, ZN => n3051);
   U1636 : OAI22_X1 port map( A1 => n10086, A2 => n14285, B1 => n10501, B2 => 
                           n14468, ZN => n14251);
   U1637 : INV_X1 port map( A => n14251, ZN => n3045);
   U1638 : OAI22_X1 port map( A1 => n10085, A2 => n14285, B1 => n10502, B2 => 
                           n14353, ZN => n14252);
   U1639 : INV_X1 port map( A => n14252, ZN => n3046);
   U1640 : OAI22_X1 port map( A1 => n11209, A2 => n14253, B1 => n10469, B2 => 
                           n14462, ZN => n14254);
   U1641 : INV_X1 port map( A => n14254, ZN => n2774);
   U1642 : OAI22_X1 port map( A1 => n11208, A2 => n14267, B1 => n10470, B2 => 
                           n14472, ZN => n14255);
   U1643 : INV_X1 port map( A => n14255, ZN => n2788);
   U1644 : OAI22_X1 port map( A1 => n11223, A2 => n14267, B1 => n10471, B2 => 
                           n14361, ZN => n14256);
   U1645 : INV_X1 port map( A => n14256, ZN => n2789);
   U1646 : OAI22_X1 port map( A1 => n10081, A2 => n14285, B1 => n10506, B2 => 
                           n14466, ZN => n14257);
   U1647 : INV_X1 port map( A => n14257, ZN => n3050);
   U1648 : OAI22_X1 port map( A1 => n11207, A2 => n14267, B1 => n10472, B2 => 
                           n14468, ZN => n14258);
   U1649 : INV_X1 port map( A => n14258, ZN => n2790);
   U1650 : OAI22_X1 port map( A1 => n11206, A2 => n14267, B1 => n10473, B2 => 
                           n14353, ZN => n14259);
   U1651 : INV_X1 port map( A => n14259, ZN => n2791);
   U1652 : OAI22_X1 port map( A1 => n10084, A2 => n14490, B1 => n10423, B2 => 
                           n14470, ZN => n14260);
   U1653 : INV_X1 port map( A => n14260, ZN => n3015);
   U1654 : OAI22_X1 port map( A1 => n11210, A2 => n14261, B1 => n10193, B2 => 
                           n14464, ZN => n14262);
   U1655 : INV_X1 port map( A => n14262, ZN => n2627);
   U1656 : OAI22_X1 port map( A1 => n10079, A2 => n14285, B1 => n10487, B2 => 
                           n14460, ZN => n14263);
   U1657 : INV_X1 port map( A => n14263, ZN => n3052);
   U1658 : OAI22_X1 port map( A1 => n10078, A2 => n14285, B1 => n10488, B2 => 
                           n14476, ZN => n14264);
   U1659 : INV_X1 port map( A => n14264, ZN => n3053);
   U1660 : OAI22_X1 port map( A1 => n11208, A2 => n14344, B1 => n10376, B2 => 
                           n14472, ZN => n14265);
   U1661 : INV_X1 port map( A => n14265, ZN => n2756);
   U1662 : OAI22_X1 port map( A1 => n10077, A2 => n14285, B1 => n10489, B2 => 
                           n14474, ZN => n14266);
   U1663 : INV_X1 port map( A => n14266, ZN => n3054);
   U1664 : OAI22_X1 port map( A1 => n11205, A2 => n14267, B1 => n10474, B2 => 
                           n14470, ZN => n14268);
   U1665 : INV_X1 port map( A => n14268, ZN => n2792);
   U1666 : OAI22_X1 port map( A1 => n11205, A2 => n14334, B1 => n10596, B2 => 
                           n14470, ZN => n14269);
   U1667 : INV_X1 port map( A => n14269, ZN => n2823);
   U1668 : OAI22_X1 port map( A1 => n11205, A2 => n14337, B1 => n10566, B2 => 
                           n14470, ZN => n14270);
   U1669 : INV_X1 port map( A => n14270, ZN => n2855);
   U1670 : OAI22_X1 port map( A1 => n11205, A2 => n14271, B1 => n10412, B2 => 
                           n14470, ZN => n14272);
   U1671 : INV_X1 port map( A => n14272, ZN => n2887);
   U1672 : OAI22_X1 port map( A1 => n10084, A2 => n14488, B1 => n10654, B2 => 
                           n14470, ZN => n14273);
   U1673 : INV_X1 port map( A => n14273, ZN => n2919);
   U1674 : OAI22_X1 port map( A1 => n10084, A2 => n14274, B1 => n10624, B2 => 
                           n14470, ZN => n14275);
   U1675 : INV_X1 port map( A => n14275, ZN => n2951);
   U1676 : OAI22_X1 port map( A1 => n10084, A2 => n14276, B1 => n10533, B2 => 
                           n14470, ZN => n14277);
   U1677 : INV_X1 port map( A => n14277, ZN => n2983);
   U1678 : OAI22_X1 port map( A1 => n10084, A2 => n14484, B1 => n10804, B2 => 
                           n14470, ZN => n14278);
   U1679 : INV_X1 port map( A => n14278, ZN => n3079);
   U1680 : OAI22_X1 port map( A1 => n10084, A2 => n14285, B1 => n10503, B2 => 
                           n14470, ZN => n14279);
   U1681 : INV_X1 port map( A => n14279, ZN => n3047);
   U1682 : OAI22_X1 port map( A1 => n10084, A2 => n14280, B1 => n10834, B2 => 
                           n14470, ZN => n14281);
   U1683 : INV_X1 port map( A => n14281, ZN => n3143);
   U1684 : OAI22_X1 port map( A1 => n10084, A2 => n14282, B1 => n10775, B2 => 
                           n14470, ZN => n14283);
   U1685 : INV_X1 port map( A => n14283, ZN => n3111);
   U1686 : OAI22_X1 port map( A1 => n10082, A2 => n14285, B1 => n10505, B2 => 
                           n14417, ZN => n14284);
   U1687 : INV_X1 port map( A => n14284, ZN => n3049);
   U1688 : OAI22_X1 port map( A1 => n10083, A2 => n14285, B1 => n10504, B2 => 
                           n14458, ZN => n14286);
   U1689 : INV_X1 port map( A => n14286, ZN => n3048);
   U1690 : OAI22_X1 port map( A1 => n10084, A2 => n14287, B1 => n10864, B2 => 
                           n14470, ZN => n14288);
   U1691 : INV_X1 port map( A => n14288, ZN => n3175);
   U1692 : CLKBUF_X1 port map( A => n14289, Z => n14450);
   U1693 : OAI22_X1 port map( A1 => n10156, A2 => n14450, B1 => n10093, B2 => 
                           n14479, ZN => n14290);
   U1694 : INV_X1 port map( A => n14290, ZN => n3550);
   U1695 : CLKBUF_X1 port map( A => n14291, Z => n14456);
   U1696 : OAI22_X1 port map( A1 => n10157, A2 => n14456, B1 => n10092, B2 => 
                           n14479, ZN => n14292);
   U1697 : INV_X1 port map( A => n14292, ZN => n3551);
   U1698 : CLKBUF_X1 port map( A => n14293, Z => n14454);
   U1699 : OAI22_X1 port map( A1 => n10155, A2 => n14454, B1 => n10094, B2 => 
                           n14479, ZN => n14294);
   U1700 : INV_X1 port map( A => n14294, ZN => n3549);
   U1701 : CLKBUF_X1 port map( A => n14295, Z => n14306);
   U1702 : OAI22_X1 port map( A1 => n11222, A2 => n14306, B1 => n10953, B2 => 
                           n14408, ZN => n14296);
   U1703 : INV_X1 port map( A => n14296, ZN => n3223);
   U1704 : OAI22_X1 port map( A1 => n11209, A2 => n14306, B1 => n10941, B2 => 
                           n14462, ZN => n14297);
   U1705 : INV_X1 port map( A => n14297, ZN => n3234);
   U1706 : OAI22_X1 port map( A1 => n11215, A2 => n14306, B1 => n10955, B2 => 
                           n14410, ZN => n14298);
   U1707 : INV_X1 port map( A => n14298, ZN => n3221);
   U1708 : OAI22_X1 port map( A1 => n11218, A2 => n14306, B1 => n10951, B2 => 
                           n14422, ZN => n14299);
   U1709 : INV_X1 port map( A => n14299, ZN => n3225);
   U1710 : OAI22_X1 port map( A1 => n11223, A2 => n14306, B1 => n10943, B2 => 
                           n14361, ZN => n14300);
   U1711 : INV_X1 port map( A => n14300, ZN => n3236);
   U1712 : OAI22_X1 port map( A1 => n11216, A2 => n14306, B1 => n10954, B2 => 
                           n14419, ZN => n14301);
   U1713 : INV_X1 port map( A => n14301, ZN => n3222);
   U1714 : OAI22_X1 port map( A1 => n11217, A2 => n14306, B1 => n10952, B2 => 
                           n14404, ZN => n14302);
   U1715 : INV_X1 port map( A => n14302, ZN => n3224);
   U1716 : OAI22_X1 port map( A1 => n11219, A2 => n14306, B1 => n10950, B2 => 
                           n14406, ZN => n14303);
   U1717 : INV_X1 port map( A => n14303, ZN => n3226);
   U1718 : OAI22_X1 port map( A1 => n11203, A2 => n14306, B1 => n10926, B2 => 
                           n14417, ZN => n14304);
   U1719 : INV_X1 port map( A => n14304, ZN => n3241);
   U1720 : OAI22_X1 port map( A1 => n11221, A2 => n14306, B1 => n10948, B2 => 
                           n14358, ZN => n14305);
   U1721 : INV_X1 port map( A => n14305, ZN => n3228);
   U1722 : OAI22_X1 port map( A1 => n11220, A2 => n14306, B1 => n10949, B2 => 
                           n14365, ZN => n14307);
   U1723 : INV_X1 port map( A => n14307, ZN => n3227);
   U1724 : CLKBUF_X1 port map( A => n14308, Z => n14493);
   U1725 : OAI22_X1 port map( A1 => n10158, A2 => n14493, B1 => n10091, B2 => 
                           n14479, ZN => n14309);
   U1726 : INV_X1 port map( A => n14309, ZN => n3552);
   U1727 : CLKBUF_X1 port map( A => n14619, Z => n14499);
   U1728 : OAI22_X1 port map( A1 => n10098, A2 => n14499, B1 => n11044, B2 => 
                           n14314, ZN => n14310);
   U1729 : INV_X1 port map( A => n14310, ZN => n3320);
   U1730 : OAI22_X1 port map( A1 => n10096, A2 => n14499, B1 => n11046, B2 => 
                           n14316, ZN => n14311);
   U1731 : INV_X1 port map( A => n14311, ZN => n3318);
   U1732 : OAI22_X1 port map( A1 => n10095, A2 => n14499, B1 => n11047, B2 => 
                           n14318, ZN => n14312);
   U1733 : INV_X1 port map( A => n14312, ZN => n3317);
   U1734 : OAI22_X1 port map( A1 => n10101, A2 => n14499, B1 => n11041, B2 => 
                           n14320, ZN => n14313);
   U1735 : INV_X1 port map( A => n14313, ZN => n3323);
   U1736 : CLKBUF_X1 port map( A => n14488, Z => n14412);
   U1737 : OAI22_X1 port map( A1 => n10098, A2 => n14412, B1 => n10751, B2 => 
                           n14314, ZN => n14315);
   U1738 : INV_X1 port map( A => n14315, ZN => n2904);
   U1739 : OAI22_X1 port map( A1 => n10096, A2 => n14412, B1 => n10753, B2 => 
                           n14316, ZN => n14317);
   U1740 : INV_X1 port map( A => n14317, ZN => n2902);
   U1741 : OAI22_X1 port map( A1 => n10095, A2 => n14412, B1 => n10754, B2 => 
                           n14318, ZN => n14319);
   U1742 : INV_X1 port map( A => n14319, ZN => n2901);
   U1743 : OAI22_X1 port map( A1 => n10101, A2 => n14412, B1 => n10769, B2 => 
                           n14320, ZN => n14321);
   U1744 : INV_X1 port map( A => n14321, ZN => n2907);
   U1745 : OAI22_X1 port map( A1 => n10097, A2 => n14499, B1 => n11045, B2 => 
                           n14323, ZN => n14322);
   U1746 : INV_X1 port map( A => n14322, ZN => n3319);
   U1747 : OAI22_X1 port map( A1 => n10097, A2 => n14412, B1 => n10752, B2 => 
                           n14323, ZN => n14324);
   U1748 : INV_X1 port map( A => n14324, ZN => n2903);
   U1749 : OAI22_X1 port map( A1 => n10100, A2 => n14499, B1 => n11042, B2 => 
                           n14332, ZN => n14325);
   U1750 : INV_X1 port map( A => n14325, ZN => n3322);
   U1751 : OAI22_X1 port map( A1 => n10099, A2 => n14499, B1 => n11043, B2 => 
                           n14327, ZN => n14326);
   U1752 : INV_X1 port map( A => n14326, ZN => n3321);
   U1753 : OAI22_X1 port map( A1 => n10099, A2 => n14412, B1 => n10750, B2 => 
                           n14327, ZN => n14328);
   U1754 : INV_X1 port map( A => n14328, ZN => n2905);
   U1755 : OAI22_X1 port map( A1 => n10102, A2 => n14412, B1 => n10768, B2 => 
                           n14330, ZN => n14329);
   U1756 : INV_X1 port map( A => n14329, ZN => n2908);
   U1757 : OAI22_X1 port map( A1 => n10102, A2 => n14499, B1 => n11040, B2 => 
                           n14330, ZN => n14331);
   U1758 : INV_X1 port map( A => n14331, ZN => n3324);
   U1759 : OAI22_X1 port map( A1 => n10100, A2 => n14412, B1 => n10770, B2 => 
                           n14332, ZN => n14333);
   U1760 : INV_X1 port map( A => n14333, ZN => n2906);
   U1761 : CLKBUF_X1 port map( A => n14334, Z => n14381);
   U1762 : OAI22_X1 port map( A1 => n11215, A2 => n14381, B1 => n10482, B2 => 
                           n14410, ZN => n14335);
   U1763 : INV_X1 port map( A => n14335, ZN => n2805);
   U1764 : OAI22_X1 port map( A1 => n11209, A2 => n14381, B1 => n10591, B2 => 
                           n14462, ZN => n14336);
   U1765 : INV_X1 port map( A => n14336, ZN => n2818);
   U1766 : CLKBUF_X1 port map( A => n14337, Z => n14355);
   U1767 : OAI22_X1 port map( A1 => n11215, A2 => n14355, B1 => n10576, B2 => 
                           n14410, ZN => n14338);
   U1768 : INV_X1 port map( A => n14338, ZN => n2837);
   U1769 : OAI22_X1 port map( A1 => n11216, A2 => n14381, B1 => n10481, B2 => 
                           n14419, ZN => n14339);
   U1770 : INV_X1 port map( A => n14339, ZN => n2806);
   U1771 : OAI22_X1 port map( A1 => n11216, A2 => n14355, B1 => n10575, B2 => 
                           n14419, ZN => n14340);
   U1772 : INV_X1 port map( A => n14340, ZN => n2838);
   U1773 : OAI22_X1 port map( A1 => n11222, A2 => n14381, B1 => n10480, B2 => 
                           n14408, ZN => n14341);
   U1774 : INV_X1 port map( A => n14341, ZN => n2807);
   U1775 : OAI22_X1 port map( A1 => n11217, A2 => n14381, B1 => n10479, B2 => 
                           n14404, ZN => n14342);
   U1776 : INV_X1 port map( A => n14342, ZN => n2808);
   U1777 : OAI22_X1 port map( A1 => n11222, A2 => n14355, B1 => n10574, B2 => 
                           n14408, ZN => n14343);
   U1778 : INV_X1 port map( A => n14343, ZN => n2839);
   U1779 : CLKBUF_X1 port map( A => n14344, Z => n14420);
   U1780 : OAI22_X1 port map( A1 => n11219, A2 => n14420, B1 => n10385, B2 => 
                           n14406, ZN => n14345);
   U1781 : INV_X1 port map( A => n14345, ZN => n2748);
   U1782 : OAI22_X1 port map( A1 => n11217, A2 => n14355, B1 => n10573, B2 => 
                           n14404, ZN => n14346);
   U1783 : INV_X1 port map( A => n14346, ZN => n2840);
   U1784 : OAI22_X1 port map( A1 => n11208, A2 => n14381, B1 => n10592, B2 => 
                           n14472, ZN => n14347);
   U1785 : INV_X1 port map( A => n14347, ZN => n2819);
   U1786 : OAI22_X1 port map( A1 => n11218, A2 => n14355, B1 => n10572, B2 => 
                           n14422, ZN => n14348);
   U1787 : INV_X1 port map( A => n14348, ZN => n2841);
   U1788 : OAI22_X1 port map( A1 => n11219, A2 => n14355, B1 => n10571, B2 => 
                           n14406, ZN => n14349);
   U1789 : INV_X1 port map( A => n14349, ZN => n2842);
   U1790 : OAI22_X1 port map( A1 => n11220, A2 => n14355, B1 => n10570, B2 => 
                           n14365, ZN => n14350);
   U1791 : INV_X1 port map( A => n14350, ZN => n2843);
   U1792 : OAI22_X1 port map( A1 => n10102, A2 => n14355, B1 => n10569, B2 => 
                           n14358, ZN => n14351);
   U1793 : INV_X1 port map( A => n14351, ZN => n2844);
   U1794 : OAI22_X1 port map( A1 => n11208, A2 => n14355, B1 => n10562, B2 => 
                           n14472, ZN => n14352);
   U1795 : INV_X1 port map( A => n14352, ZN => n2851);
   U1796 : CLKBUF_X1 port map( A => n14353, Z => n14583);
   U1797 : OAI22_X1 port map( A1 => n10142, A2 => n14583, B1 => n10085, B2 => 
                           n14373, ZN => n14354);
   U1798 : INV_X1 port map( A => n14354, ZN => n3558);
   U1799 : OAI22_X1 port map( A1 => n11209, A2 => n14355, B1 => n10561, B2 => 
                           n14462, ZN => n14356);
   U1800 : INV_X1 port map( A => n14356, ZN => n2850);
   U1801 : OAI22_X1 port map( A1 => n11218, A2 => n14420, B1 => n10386, B2 => 
                           n14422, ZN => n14357);
   U1802 : INV_X1 port map( A => n14357, ZN => n2747);
   U1803 : OAI22_X1 port map( A1 => n10102, A2 => n14381, B1 => n10475, B2 => 
                           n14358, ZN => n14359);
   U1804 : INV_X1 port map( A => n14359, ZN => n2812);
   U1805 : OAI22_X1 port map( A1 => n10089, A2 => n14412, B1 => n10760, B2 => 
                           n14462, ZN => n14360);
   U1806 : INV_X1 port map( A => n14360, ZN => n2914);
   U1807 : CLKBUF_X1 port map( A => n14361, Z => n14580);
   U1808 : OAI22_X1 port map( A1 => n10162, A2 => n14580, B1 => n10087, B2 => 
                           n14373, ZN => n14362);
   U1809 : INV_X1 port map( A => n14362, ZN => n3556);
   U1810 : CLKBUF_X1 port map( A => n14363, Z => n14400);
   U1811 : OAI22_X1 port map( A1 => n11198, A2 => n14400, B1 => n10195, B2 => 
                           n14414, ZN => n14364);
   U1812 : INV_X1 port map( A => n14364, ZN => n2607);
   U1813 : OAI22_X1 port map( A1 => n11220, A2 => n14381, B1 => n10476, B2 => 
                           n14365, ZN => n14366);
   U1814 : INV_X1 port map( A => n14366, ZN => n2811);
   U1815 : OAI22_X1 port map( A1 => n11219, A2 => n14381, B1 => n10477, B2 => 
                           n14406, ZN => n14367);
   U1816 : INV_X1 port map( A => n14367, ZN => n2810);
   U1817 : OAI22_X1 port map( A1 => n11200, A2 => n14400, B1 => n10213, B2 => 
                           n14476, ZN => n14368);
   U1818 : INV_X1 port map( A => n14368, ZN => n2605);
   U1819 : OAI22_X1 port map( A1 => n11218, A2 => n14400, B1 => n10214, B2 => 
                           n14422, ZN => n14369);
   U1820 : INV_X1 port map( A => n14369, ZN => n2587);
   U1821 : OAI22_X1 port map( A1 => n11217, A2 => n14400, B1 => n10215, B2 => 
                           n14404, ZN => n14370);
   U1822 : INV_X1 port map( A => n14370, ZN => n2586);
   U1823 : OAI22_X1 port map( A1 => n11222, A2 => n14400, B1 => n10216, B2 => 
                           n14408, ZN => n14371);
   U1824 : INV_X1 port map( A => n14371, ZN => n2585);
   U1825 : OAI22_X1 port map( A1 => n11216, A2 => n14400, B1 => n10217, B2 => 
                           n14419, ZN => n14372);
   U1826 : INV_X1 port map( A => n14372, ZN => n2584);
   U1827 : CLKBUF_X1 port map( A => n14417, Z => n14618);
   U1828 : OAI22_X1 port map( A1 => n10145, A2 => n14618, B1 => n10082, B2 => 
                           n14373, ZN => n14374);
   U1829 : INV_X1 port map( A => n14374, ZN => n3561);
   U1830 : CLKBUF_X1 port map( A => n14375, Z => n14395);
   U1831 : OAI22_X1 port map( A1 => n11215, A2 => n14395, B1 => n10283, B2 => 
                           n14410, ZN => n14376);
   U1832 : INV_X1 port map( A => n14376, ZN => n2647);
   U1833 : OAI22_X1 port map( A1 => n11215, A2 => n14400, B1 => n10218, B2 => 
                           n14410, ZN => n14377);
   U1834 : INV_X1 port map( A => n14377, ZN => n2583);
   U1835 : OAI22_X1 port map( A1 => n11216, A2 => n14395, B1 => n10282, B2 => 
                           n14419, ZN => n14378);
   U1836 : INV_X1 port map( A => n14378, ZN => n2648);
   U1837 : OAI22_X1 port map( A1 => n11222, A2 => n14395, B1 => n10281, B2 => 
                           n14408, ZN => n14379);
   U1838 : INV_X1 port map( A => n14379, ZN => n2649);
   U1839 : OAI22_X1 port map( A1 => n11217, A2 => n14395, B1 => n10280, B2 => 
                           n14404, ZN => n14380);
   U1840 : INV_X1 port map( A => n14380, ZN => n2650);
   U1841 : OAI22_X1 port map( A1 => n11218, A2 => n14381, B1 => n10478, B2 => 
                           n14422, ZN => n14382);
   U1842 : INV_X1 port map( A => n14382, ZN => n2809);
   U1843 : OAI22_X1 port map( A1 => n11203, A2 => n14400, B1 => n10209, B2 => 
                           n14417, ZN => n14383);
   U1844 : INV_X1 port map( A => n14383, ZN => n2581);
   U1845 : CLKBUF_X1 port map( A => n14384, Z => n14423);
   U1846 : OAI22_X1 port map( A1 => n11203, A2 => n14423, B1 => n10244, B2 => 
                           n14417, ZN => n14385);
   U1847 : INV_X1 port map( A => n14385, ZN => n2677);
   U1848 : OAI22_X1 port map( A1 => n11209, A2 => n14420, B1 => n10375, B2 => 
                           n14462, ZN => n14386);
   U1849 : INV_X1 port map( A => n14386, ZN => n2742);
   U1850 : OAI22_X1 port map( A1 => n11218, A2 => n14395, B1 => n10279, B2 => 
                           n14422, ZN => n14387);
   U1851 : INV_X1 port map( A => n14387, ZN => n2651);
   U1852 : OAI22_X1 port map( A1 => n11219, A2 => n14395, B1 => n10278, B2 => 
                           n14406, ZN => n14388);
   U1853 : INV_X1 port map( A => n14388, ZN => n2652);
   U1854 : OAI22_X1 port map( A1 => n11209, A2 => n14400, B1 => n10224, B2 => 
                           n14462, ZN => n14389);
   U1855 : INV_X1 port map( A => n14389, ZN => n2582);
   U1856 : OAI22_X1 port map( A1 => n11200, A2 => n14423, B1 => n10227, B2 => 
                           n14476, ZN => n14390);
   U1857 : INV_X1 port map( A => n14390, ZN => n2701);
   U1858 : OAI22_X1 port map( A1 => n11198, A2 => n14423, B1 => n10229, B2 => 
                           n14414, ZN => n14391);
   U1859 : INV_X1 port map( A => n14391, ZN => n2703);
   U1860 : OAI22_X1 port map( A1 => n11203, A2 => n14395, B1 => n10274, B2 => 
                           n14417, ZN => n14392);
   U1861 : INV_X1 port map( A => n14392, ZN => n2645);
   U1862 : OAI22_X1 port map( A1 => n11209, A2 => n14395, B1 => n10267, B2 => 
                           n14462, ZN => n14393);
   U1863 : INV_X1 port map( A => n14393, ZN => n2646);
   U1864 : OAI22_X1 port map( A1 => n11198, A2 => n14395, B1 => n10260, B2 => 
                           n14414, ZN => n14394);
   U1865 : INV_X1 port map( A => n14394, ZN => n2671);
   U1866 : OAI22_X1 port map( A1 => n11200, A2 => n14395, B1 => n10258, B2 => 
                           n14476, ZN => n14396);
   U1867 : INV_X1 port map( A => n14396, ZN => n2669);
   U1868 : OAI22_X1 port map( A1 => n11215, A2 => n14423, B1 => n10253, B2 => 
                           n14410, ZN => n14397);
   U1869 : INV_X1 port map( A => n14397, ZN => n2679);
   U1870 : OAI22_X1 port map( A1 => n11209, A2 => n14423, B1 => n10237, B2 => 
                           n14462, ZN => n14398);
   U1871 : INV_X1 port map( A => n14398, ZN => n2678);
   U1872 : OAI22_X1 port map( A1 => n11216, A2 => n14423, B1 => n10252, B2 => 
                           n14419, ZN => n14399);
   U1873 : INV_X1 port map( A => n14399, ZN => n2680);
   U1874 : OAI22_X1 port map( A1 => n11219, A2 => n14400, B1 => n10109, B2 => 
                           n14406, ZN => n14401);
   U1875 : INV_X1 port map( A => n14401, ZN => n2588);
   U1876 : OAI22_X1 port map( A1 => n11222, A2 => n14423, B1 => n10251, B2 => 
                           n14408, ZN => n14402);
   U1877 : INV_X1 port map( A => n14402, ZN => n2681);
   U1878 : OAI22_X1 port map( A1 => n11217, A2 => n14423, B1 => n10250, B2 => 
                           n14404, ZN => n14403);
   U1879 : INV_X1 port map( A => n14403, ZN => n2682);
   U1880 : OAI22_X1 port map( A1 => n11217, A2 => n14420, B1 => n10387, B2 => 
                           n14404, ZN => n14405);
   U1881 : INV_X1 port map( A => n14405, ZN => n2746);
   U1882 : OAI22_X1 port map( A1 => n11219, A2 => n14423, B1 => n10248, B2 => 
                           n14406, ZN => n14407);
   U1883 : INV_X1 port map( A => n14407, ZN => n2684);
   U1884 : OAI22_X1 port map( A1 => n11222, A2 => n14420, B1 => n10388, B2 => 
                           n14408, ZN => n14409);
   U1885 : INV_X1 port map( A => n14409, ZN => n2745);
   U1886 : OAI22_X1 port map( A1 => n11215, A2 => n14420, B1 => n10390, B2 => 
                           n14410, ZN => n14411);
   U1887 : INV_X1 port map( A => n14411, ZN => n2743);
   U1888 : OAI22_X1 port map( A1 => n10088, A2 => n14412, B1 => n10650, B2 => 
                           n14472, ZN => n14413);
   U1889 : INV_X1 port map( A => n14413, ZN => n2915);
   U1890 : OAI22_X1 port map( A1 => n11198, A2 => n14420, B1 => n10366, B2 => 
                           n14414, ZN => n14415);
   U1891 : INV_X1 port map( A => n14415, ZN => n2767);
   U1892 : OAI22_X1 port map( A1 => n11200, A2 => n14420, B1 => n10364, B2 => 
                           n14476, ZN => n14416);
   U1893 : INV_X1 port map( A => n14416, ZN => n2765);
   U1894 : OAI22_X1 port map( A1 => n11203, A2 => n14420, B1 => n10360, B2 => 
                           n14417, ZN => n14418);
   U1895 : INV_X1 port map( A => n14418, ZN => n2741);
   U1896 : OAI22_X1 port map( A1 => n11216, A2 => n14420, B1 => n10389, B2 => 
                           n14419, ZN => n14421);
   U1897 : INV_X1 port map( A => n14421, ZN => n2744);
   U1898 : OAI22_X1 port map( A1 => n11218, A2 => n14423, B1 => n10249, B2 => 
                           n14422, ZN => n14424);
   U1899 : INV_X1 port map( A => n14424, ZN => n2683);
   U1900 : OAI22_X1 port map( A1 => n10092, A2 => n14594, B1 => n10344, B2 => 
                           n14456, ZN => n14425);
   U1901 : INV_X1 port map( A => n14425, ZN => n3487);
   U1902 : OAI22_X1 port map( A1 => n10093, A2 => n14594, B1 => n10343, B2 => 
                           n14450, ZN => n14426);
   U1903 : INV_X1 port map( A => n14426, ZN => n3486);
   U1904 : OAI22_X1 port map( A1 => n10093, A2 => n14488, B1 => n10756, B2 => 
                           n14450, ZN => n14427);
   U1905 : INV_X1 port map( A => n14427, ZN => n2910);
   U1906 : OAI22_X1 port map( A1 => n10093, A2 => n14490, B1 => n10436, B2 => 
                           n14450, ZN => n14428);
   U1907 : INV_X1 port map( A => n14428, ZN => n3006);
   U1908 : OAI22_X1 port map( A1 => n10093, A2 => n14484, B1 => n10817, B2 => 
                           n14450, ZN => n14429);
   U1909 : INV_X1 port map( A => n14429, ZN => n3070);
   U1910 : OAI22_X1 port map( A1 => n10092, A2 => n14488, B1 => n10757, B2 => 
                           n14456, ZN => n14430);
   U1911 : INV_X1 port map( A => n14430, ZN => n2911);
   U1912 : OAI22_X1 port map( A1 => n10092, A2 => n14490, B1 => n10437, B2 => 
                           n14456, ZN => n14431);
   U1913 : INV_X1 port map( A => n14431, ZN => n3007);
   U1914 : OAI22_X1 port map( A1 => n10094, A2 => n14594, B1 => n10342, B2 => 
                           n14454, ZN => n14432);
   U1915 : INV_X1 port map( A => n14432, ZN => n3485);
   U1916 : OAI22_X1 port map( A1 => n10093, A2 => n14599, B1 => n10735, B2 => 
                           n14450, ZN => n14433);
   U1917 : INV_X1 port map( A => n14433, ZN => n3454);
   U1918 : OAI22_X1 port map( A1 => n10094, A2 => n14488, B1 => n10755, B2 => 
                           n14454, ZN => n14434);
   U1919 : INV_X1 port map( A => n14434, ZN => n2909);
   U1920 : OAI22_X1 port map( A1 => n10094, A2 => n14610, B1 => n11078, B2 => 
                           n14454, ZN => n14435);
   U1921 : INV_X1 port map( A => n14435, ZN => n3357);
   U1922 : OAI22_X1 port map( A1 => n10094, A2 => n14619, B1 => n11048, B2 => 
                           n14454, ZN => n14436);
   U1923 : INV_X1 port map( A => n14436, ZN => n3325);
   U1924 : OAI22_X1 port map( A1 => n10094, A2 => n14599, B1 => n10734, B2 => 
                           n14454, ZN => n14437);
   U1925 : INV_X1 port map( A => n14437, ZN => n3453);
   U1926 : OAI22_X1 port map( A1 => n10093, A2 => n14604, B1 => n10705, B2 => 
                           n14450, ZN => n14438);
   U1927 : INV_X1 port map( A => n14438, ZN => n3422);
   U1928 : OAI22_X1 port map( A1 => n10093, A2 => n14619, B1 => n11049, B2 => 
                           n14450, ZN => n14439);
   U1929 : INV_X1 port map( A => n14439, ZN => n3326);
   U1930 : OAI22_X1 port map( A1 => n10093, A2 => n14573, B1 => n11109, B2 => 
                           n14450, ZN => n14440);
   U1931 : INV_X1 port map( A => n14440, ZN => n3390);
   U1932 : OAI22_X1 port map( A1 => n10092, A2 => n14619, B1 => n11050, B2 => 
                           n14456, ZN => n14441);
   U1933 : INV_X1 port map( A => n14441, ZN => n3327);
   U1934 : OAI22_X1 port map( A1 => n10094, A2 => n14591, B1 => n10675, B2 => 
                           n14454, ZN => n14442);
   U1935 : INV_X1 port map( A => n14442, ZN => n3517);
   U1936 : OAI22_X1 port map( A1 => n10094, A2 => n14484, B1 => n10816, B2 => 
                           n14454, ZN => n14443);
   U1937 : INV_X1 port map( A => n14443, ZN => n3069);
   U1938 : OAI22_X1 port map( A1 => n10092, A2 => n14599, B1 => n10736, B2 => 
                           n14456, ZN => n14444);
   U1939 : INV_X1 port map( A => n14444, ZN => n3455);
   U1940 : OAI22_X1 port map( A1 => n10092, A2 => n14484, B1 => n10818, B2 => 
                           n14456, ZN => n14445);
   U1941 : INV_X1 port map( A => n14445, ZN => n3071);
   U1942 : OAI22_X1 port map( A1 => n10094, A2 => n14490, B1 => n10435, B2 => 
                           n14454, ZN => n14446);
   U1943 : INV_X1 port map( A => n14446, ZN => n3005);
   U1944 : OAI22_X1 port map( A1 => n10092, A2 => n14604, B1 => n10706, B2 => 
                           n14456, ZN => n14447);
   U1945 : INV_X1 port map( A => n14447, ZN => n3423);
   U1946 : OAI22_X1 port map( A1 => n10093, A2 => n14591, B1 => n10676, B2 => 
                           n14450, ZN => n14448);
   U1947 : INV_X1 port map( A => n14448, ZN => n3518);
   U1948 : OAI22_X1 port map( A1 => n10094, A2 => n14604, B1 => n10704, B2 => 
                           n14454, ZN => n14449);
   U1949 : INV_X1 port map( A => n14449, ZN => n3421);
   U1950 : OAI22_X1 port map( A1 => n10093, A2 => n14610, B1 => n11079, B2 => 
                           n14450, ZN => n14451);
   U1951 : INV_X1 port map( A => n14451, ZN => n3358);
   U1952 : OAI22_X1 port map( A1 => n10092, A2 => n14610, B1 => n11080, B2 => 
                           n14456, ZN => n14452);
   U1953 : INV_X1 port map( A => n14452, ZN => n3359);
   U1954 : OAI22_X1 port map( A1 => n10092, A2 => n14591, B1 => n10677, B2 => 
                           n14456, ZN => n14453);
   U1955 : INV_X1 port map( A => n14453, ZN => n3519);
   U1956 : OAI22_X1 port map( A1 => n10094, A2 => n14573, B1 => n11108, B2 => 
                           n14454, ZN => n14455);
   U1957 : INV_X1 port map( A => n14455, ZN => n3389);
   U1958 : OAI22_X1 port map( A1 => n10092, A2 => n14573, B1 => n11110, B2 => 
                           n14456, ZN => n14457);
   U1959 : INV_X1 port map( A => n14457, ZN => n3391);
   U1960 : CLKBUF_X1 port map( A => n14458, Z => n14597);
   U1961 : OAI22_X1 port map( A1 => n10144, A2 => n14597, B1 => n10083, B2 => 
                           n14479, ZN => n14459);
   U1962 : INV_X1 port map( A => n14459, ZN => n3560);
   U1963 : CLKBUF_X1 port map( A => n14460, Z => n14601);
   U1964 : OAI22_X1 port map( A1 => n10148, A2 => n14601, B1 => n10079, B2 => 
                           n14479, ZN => n14461);
   U1965 : INV_X1 port map( A => n14461, ZN => n3564);
   U1966 : CLKBUF_X1 port map( A => n14462, Z => n14515);
   U1967 : OAI22_X1 port map( A1 => n10160, A2 => n14515, B1 => n10089, B2 => 
                           n14479, ZN => n14463);
   U1968 : INV_X1 port map( A => n14463, ZN => n3554);
   U1969 : CLKBUF_X1 port map( A => n14464, Z => n14612);
   U1970 : OAI22_X1 port map( A1 => n10159, A2 => n14612, B1 => n10090, B2 => 
                           n14479, ZN => n14465);
   U1971 : INV_X1 port map( A => n14465, ZN => n3553);
   U1972 : CLKBUF_X1 port map( A => n14466, Z => n14616);
   U1973 : OAI22_X1 port map( A1 => n10146, A2 => n14616, B1 => n10081, B2 => 
                           n14479, ZN => n14467);
   U1974 : INV_X1 port map( A => n14467, ZN => n3562);
   U1975 : CLKBUF_X1 port map( A => n14468, Z => n14603);
   U1976 : OAI22_X1 port map( A1 => n10141, A2 => n14603, B1 => n10086, B2 => 
                           n14479, ZN => n14469);
   U1977 : INV_X1 port map( A => n14469, ZN => n3557);
   U1978 : CLKBUF_X1 port map( A => n14470, Z => n14614);
   U1979 : OAI22_X1 port map( A1 => n10143, A2 => n14614, B1 => n10084, B2 => 
                           n14479, ZN => n14471);
   U1980 : INV_X1 port map( A => n14471, ZN => n3559);
   U1981 : CLKBUF_X1 port map( A => n14472, Z => n14510);
   U1982 : OAI22_X1 port map( A1 => n10161, A2 => n14510, B1 => n10088, B2 => 
                           n14479, ZN => n14473);
   U1983 : INV_X1 port map( A => n14473, ZN => n3555);
   U1984 : CLKBUF_X1 port map( A => n14474, Z => n14608);
   U1985 : OAI22_X1 port map( A1 => n10150, A2 => n14608, B1 => n10077, B2 => 
                           n14479, ZN => n14475);
   U1986 : INV_X1 port map( A => n14475, ZN => n3566);
   U1987 : CLKBUF_X1 port map( A => n14476, Z => n14606);
   U1988 : OAI22_X1 port map( A1 => n10149, A2 => n14606, B1 => n10078, B2 => 
                           n14479, ZN => n14477);
   U1989 : INV_X1 port map( A => n14477, ZN => n3565);
   U1990 : CLKBUF_X1 port map( A => n14478, Z => n14588);
   U1991 : OAI22_X1 port map( A1 => n10147, A2 => n14588, B1 => n10080, B2 => 
                           n14479, ZN => n14480);
   U1992 : INV_X1 port map( A => n14480, ZN => n3563);
   U1993 : OAI22_X1 port map( A1 => n10091, A2 => n14599, B1 => n10737, B2 => 
                           n14493, ZN => n14481);
   U1994 : INV_X1 port map( A => n14481, ZN => n3456);
   U1995 : OAI22_X1 port map( A1 => n10091, A2 => n14619, B1 => n11029, B2 => 
                           n14493, ZN => n14482);
   U1996 : INV_X1 port map( A => n14482, ZN => n3328);
   U1997 : OAI22_X1 port map( A1 => n10091, A2 => n14594, B1 => n10345, B2 => 
                           n14493, ZN => n14483);
   U1998 : INV_X1 port map( A => n14483, ZN => n3488);
   U1999 : OAI22_X1 port map( A1 => n10091, A2 => n14484, B1 => n10819, B2 => 
                           n14493, ZN => n14485);
   U2000 : INV_X1 port map( A => n14485, ZN => n3072);
   U2001 : OAI22_X1 port map( A1 => n10091, A2 => n14573, B1 => n11111, B2 => 
                           n14493, ZN => n14486);
   U2002 : INV_X1 port map( A => n14486, ZN => n3392);
   U2003 : OAI22_X1 port map( A1 => n10091, A2 => n14610, B1 => n11081, B2 => 
                           n14493, ZN => n14487);
   U2004 : INV_X1 port map( A => n14487, ZN => n3360);
   U2005 : OAI22_X1 port map( A1 => n10091, A2 => n14488, B1 => n10758, B2 => 
                           n14493, ZN => n14489);
   U2006 : INV_X1 port map( A => n14489, ZN => n2912);
   U2007 : OAI22_X1 port map( A1 => n10091, A2 => n14490, B1 => n10438, B2 => 
                           n14493, ZN => n14491);
   U2008 : INV_X1 port map( A => n14491, ZN => n3008);
   U2009 : OAI22_X1 port map( A1 => n10091, A2 => n14604, B1 => n10707, B2 => 
                           n14493, ZN => n14492);
   U2010 : INV_X1 port map( A => n14492, ZN => n3424);
   U2011 : OAI22_X1 port map( A1 => n10091, A2 => n14591, B1 => n10678, B2 => 
                           n14493, ZN => n14494);
   U2012 : INV_X1 port map( A => n14494, ZN => n3520);
   U2013 : OAI22_X1 port map( A1 => n10088, A2 => n14508, B1 => n11062, B2 => 
                           n14510, ZN => n14495);
   U2014 : INV_X1 port map( A => n14495, ZN => n3363);
   U2015 : OAI22_X1 port map( A1 => n10088, A2 => n14499, B1 => n11032, B2 => 
                           n14510, ZN => n14496);
   U2016 : INV_X1 port map( A => n14496, ZN => n3331);
   U2017 : OAI22_X1 port map( A1 => n10089, A2 => n14505, B1 => n10347, B2 => 
                           n14515, ZN => n14497);
   U2018 : INV_X1 port map( A => n14497, ZN => n3490);
   U2019 : OAI22_X1 port map( A1 => n10088, A2 => n14516, B1 => n10688, B2 => 
                           n14510, ZN => n14498);
   U2020 : INV_X1 port map( A => n14498, ZN => n3427);
   U2021 : OAI22_X1 port map( A1 => n10089, A2 => n14499, B1 => n11031, B2 => 
                           n14515, ZN => n14500);
   U2022 : INV_X1 port map( A => n14500, ZN => n3330);
   U2023 : OAI22_X1 port map( A1 => n10088, A2 => n14502, B1 => n11092, B2 => 
                           n14510, ZN => n14501);
   U2024 : INV_X1 port map( A => n14501, ZN => n3395);
   U2025 : OAI22_X1 port map( A1 => n10089, A2 => n14502, B1 => n11091, B2 => 
                           n14515, ZN => n14503);
   U2026 : INV_X1 port map( A => n14503, ZN => n3394);
   U2027 : OAI22_X1 port map( A1 => n10088, A2 => n14513, B1 => n10681, B2 => 
                           n14510, ZN => n14504);
   U2028 : INV_X1 port map( A => n14504, ZN => n3523);
   U2029 : OAI22_X1 port map( A1 => n10088, A2 => n14505, B1 => n10348, B2 => 
                           n14510, ZN => n14506);
   U2030 : INV_X1 port map( A => n14506, ZN => n3491);
   U2031 : OAI22_X1 port map( A1 => n10089, A2 => n14511, B1 => n10739, B2 => 
                           n14515, ZN => n14507);
   U2032 : INV_X1 port map( A => n14507, ZN => n3458);
   U2033 : OAI22_X1 port map( A1 => n10089, A2 => n14508, B1 => n11061, B2 => 
                           n14515, ZN => n14509);
   U2034 : INV_X1 port map( A => n14509, ZN => n3362);
   U2035 : OAI22_X1 port map( A1 => n10088, A2 => n14511, B1 => n10740, B2 => 
                           n14510, ZN => n14512);
   U2036 : INV_X1 port map( A => n14512, ZN => n3459);
   U2037 : OAI22_X1 port map( A1 => n10089, A2 => n14513, B1 => n10680, B2 => 
                           n14515, ZN => n14514);
   U2038 : INV_X1 port map( A => n14514, ZN => n3522);
   U2039 : OAI22_X1 port map( A1 => n10089, A2 => n14516, B1 => n10709, B2 => 
                           n14515, ZN => n14517);
   U2040 : INV_X1 port map( A => n14517, ZN => n3426);
   U2041 : OAI22_X1 port map( A1 => n10085, A2 => n14604, B1 => n10691, B2 => 
                           n14583, ZN => n14518);
   U2042 : INV_X1 port map( A => n14518, ZN => n3430);
   U2043 : OAI22_X1 port map( A1 => n10083, A2 => n14604, B1 => n10693, B2 => 
                           n14597, ZN => n14519);
   U2044 : INV_X1 port map( A => n14519, ZN => n3432);
   U2045 : OAI22_X1 port map( A1 => n10086, A2 => n14591, B1 => n10661, B2 => 
                           n14603, ZN => n14520);
   U2046 : INV_X1 port map( A => n14520, ZN => n3525);
   U2047 : OAI22_X1 port map( A1 => n10085, A2 => n14591, B1 => n10662, B2 => 
                           n14583, ZN => n14521);
   U2048 : INV_X1 port map( A => n14521, ZN => n3526);
   U2049 : OAI22_X1 port map( A1 => n10083, A2 => n14591, B1 => n10664, B2 => 
                           n14597, ZN => n14522);
   U2050 : INV_X1 port map( A => n14522, ZN => n3528);
   U2051 : OAI22_X1 port map( A1 => n10082, A2 => n14604, B1 => n10694, B2 => 
                           n14618, ZN => n14523);
   U2052 : INV_X1 port map( A => n14523, ZN => n3433);
   U2053 : OAI22_X1 port map( A1 => n10082, A2 => n14591, B1 => n10665, B2 => 
                           n14618, ZN => n14524);
   U2054 : INV_X1 port map( A => n14524, ZN => n3529);
   U2055 : OAI22_X1 port map( A1 => n10085, A2 => n14599, B1 => n10721, B2 => 
                           n14583, ZN => n14525);
   U2056 : INV_X1 port map( A => n14525, ZN => n3462);
   U2057 : OAI22_X1 port map( A1 => n10086, A2 => n14594, B1 => n10350, B2 => 
                           n14603, ZN => n14526);
   U2058 : INV_X1 port map( A => n14526, ZN => n3493);
   U2059 : OAI22_X1 port map( A1 => n10083, A2 => n14599, B1 => n10723, B2 => 
                           n14597, ZN => n14527);
   U2060 : INV_X1 port map( A => n14527, ZN => n3464);
   U2061 : OAI22_X1 port map( A1 => n10082, A2 => n14599, B1 => n10724, B2 => 
                           n14618, ZN => n14528);
   U2062 : INV_X1 port map( A => n14528, ZN => n3465);
   U2063 : OAI22_X1 port map( A1 => n10085, A2 => n14594, B1 => n10329, B2 => 
                           n14583, ZN => n14529);
   U2064 : INV_X1 port map( A => n14529, ZN => n3494);
   U2065 : OAI22_X1 port map( A1 => n10084, A2 => n14599, B1 => n10722, B2 => 
                           n14614, ZN => n14530);
   U2066 : INV_X1 port map( A => n14530, ZN => n3463);
   U2067 : OAI22_X1 port map( A1 => n10077, A2 => n14599, B1 => n10729, B2 => 
                           n14608, ZN => n14531);
   U2068 : INV_X1 port map( A => n14531, ZN => n3470);
   U2069 : OAI22_X1 port map( A1 => n10077, A2 => n14591, B1 => n10670, B2 => 
                           n14608, ZN => n14532);
   U2070 : INV_X1 port map( A => n14532, ZN => n3534);
   U2071 : OAI22_X1 port map( A1 => n10087, A2 => n14619, B1 => n11033, B2 => 
                           n14580, ZN => n14533);
   U2072 : INV_X1 port map( A => n14533, ZN => n3332);
   U2073 : OAI22_X1 port map( A1 => n10087, A2 => n14604, B1 => n10689, B2 => 
                           n14580, ZN => n14534);
   U2074 : INV_X1 port map( A => n14534, ZN => n3428);
   U2075 : OAI22_X1 port map( A1 => n10078, A2 => n14591, B1 => n10669, B2 => 
                           n14606, ZN => n14535);
   U2076 : INV_X1 port map( A => n14535, ZN => n3533);
   U2077 : OAI22_X1 port map( A1 => n10080, A2 => n14591, B1 => n10667, B2 => 
                           n14588, ZN => n14536);
   U2078 : INV_X1 port map( A => n14536, ZN => n3531);
   U2079 : OAI22_X1 port map( A1 => n10078, A2 => n14599, B1 => n10728, B2 => 
                           n14606, ZN => n14537);
   U2080 : INV_X1 port map( A => n14537, ZN => n3469);
   U2081 : OAI22_X1 port map( A1 => n10080, A2 => n14599, B1 => n10726, B2 => 
                           n14588, ZN => n14538);
   U2082 : INV_X1 port map( A => n14538, ZN => n3467);
   U2083 : OAI22_X1 port map( A1 => n10078, A2 => n14604, B1 => n10698, B2 => 
                           n14606, ZN => n14539);
   U2084 : INV_X1 port map( A => n14539, ZN => n3437);
   U2085 : OAI22_X1 port map( A1 => n10080, A2 => n14604, B1 => n10696, B2 => 
                           n14588, ZN => n14540);
   U2086 : INV_X1 port map( A => n14540, ZN => n3435);
   U2087 : OAI22_X1 port map( A1 => n10084, A2 => n14604, B1 => n10692, B2 => 
                           n14614, ZN => n14541);
   U2088 : INV_X1 port map( A => n14541, ZN => n3431);
   U2089 : OAI22_X1 port map( A1 => n10077, A2 => n14604, B1 => n11113, B2 => 
                           n14608, ZN => n14542);
   U2090 : INV_X1 port map( A => n14542, ZN => n3438);
   U2091 : OAI22_X1 port map( A1 => n10087, A2 => n14599, B1 => n10719, B2 => 
                           n14580, ZN => n14543);
   U2092 : INV_X1 port map( A => n14543, ZN => n3460);
   U2093 : OAI22_X1 port map( A1 => n10087, A2 => n14594, B1 => n10349, B2 => 
                           n14580, ZN => n14544);
   U2094 : INV_X1 port map( A => n14544, ZN => n3492);
   U2095 : OAI22_X1 port map( A1 => n10087, A2 => n14591, B1 => n10682, B2 => 
                           n14580, ZN => n14545);
   U2096 : INV_X1 port map( A => n14545, ZN => n3524);
   U2097 : OAI22_X1 port map( A1 => n10080, A2 => n14573, B1 => n11100, B2 => 
                           n14588, ZN => n14546);
   U2098 : INV_X1 port map( A => n14546, ZN => n3403);
   U2099 : OAI22_X1 port map( A1 => n10090, A2 => n14591, B1 => n10679, B2 => 
                           n14612, ZN => n14547);
   U2100 : INV_X1 port map( A => n14547, ZN => n3521);
   U2101 : OAI22_X1 port map( A1 => n10082, A2 => n14573, B1 => n11098, B2 => 
                           n14618, ZN => n14548);
   U2102 : INV_X1 port map( A => n14548, ZN => n3401);
   U2103 : OAI22_X1 port map( A1 => n10090, A2 => n14594, B1 => n10346, B2 => 
                           n14612, ZN => n14549);
   U2104 : INV_X1 port map( A => n14549, ZN => n3489);
   U2105 : OAI22_X1 port map( A1 => n10083, A2 => n14573, B1 => n11097, B2 => 
                           n14597, ZN => n14550);
   U2106 : INV_X1 port map( A => n14550, ZN => n3400);
   U2107 : OAI22_X1 port map( A1 => n10085, A2 => n14573, B1 => n11095, B2 => 
                           n14583, ZN => n14551);
   U2108 : INV_X1 port map( A => n14551, ZN => n3398);
   U2109 : OAI22_X1 port map( A1 => n10090, A2 => n14599, B1 => n10738, B2 => 
                           n14612, ZN => n14552);
   U2110 : INV_X1 port map( A => n14552, ZN => n3457);
   U2111 : OAI22_X1 port map( A1 => n10090, A2 => n14604, B1 => n10708, B2 => 
                           n14612, ZN => n14553);
   U2112 : INV_X1 port map( A => n14553, ZN => n3425);
   U2113 : OAI22_X1 port map( A1 => n10090, A2 => n14573, B1 => n11112, B2 => 
                           n14612, ZN => n14554);
   U2114 : INV_X1 port map( A => n14554, ZN => n3393);
   U2115 : OAI22_X1 port map( A1 => n10081, A2 => n14591, B1 => n10666, B2 => 
                           n14616, ZN => n14555);
   U2116 : INV_X1 port map( A => n14555, ZN => n3530);
   U2117 : OAI22_X1 port map( A1 => n10087, A2 => n14573, B1 => n11093, B2 => 
                           n14580, ZN => n14556);
   U2118 : INV_X1 port map( A => n14556, ZN => n3396);
   U2119 : OAI22_X1 port map( A1 => n10084, A2 => n14591, B1 => n10663, B2 => 
                           n14614, ZN => n14557);
   U2120 : INV_X1 port map( A => n14557, ZN => n3527);
   U2121 : OAI22_X1 port map( A1 => n10084, A2 => n14573, B1 => n11096, B2 => 
                           n14614, ZN => n14558);
   U2122 : INV_X1 port map( A => n14558, ZN => n3399);
   U2123 : OAI22_X1 port map( A1 => n10077, A2 => n14573, B1 => n11083, B2 => 
                           n14608, ZN => n14559);
   U2124 : INV_X1 port map( A => n14559, ZN => n3406);
   U2125 : OAI22_X1 port map( A1 => n10081, A2 => n14599, B1 => n10725, B2 => 
                           n14616, ZN => n14560);
   U2126 : INV_X1 port map( A => n14560, ZN => n3466);
   U2127 : OAI22_X1 port map( A1 => n10078, A2 => n14573, B1 => n11082, B2 => 
                           n14606, ZN => n14561);
   U2128 : INV_X1 port map( A => n14561, ZN => n3405);
   U2129 : OAI22_X1 port map( A1 => n10079, A2 => n14573, B1 => n11101, B2 => 
                           n14601, ZN => n14562);
   U2130 : INV_X1 port map( A => n14562, ZN => n3404);
   U2131 : OAI22_X1 port map( A1 => n10079, A2 => n14604, B1 => n10697, B2 => 
                           n14601, ZN => n14563);
   U2132 : INV_X1 port map( A => n14563, ZN => n3436);
   U2133 : OAI22_X1 port map( A1 => n10079, A2 => n14599, B1 => n10727, B2 => 
                           n14601, ZN => n14564);
   U2134 : INV_X1 port map( A => n14564, ZN => n3468);
   U2135 : OAI22_X1 port map( A1 => n10080, A2 => n14610, B1 => n11070, B2 => 
                           n14588, ZN => n14565);
   U2136 : INV_X1 port map( A => n14565, ZN => n3371);
   U2137 : OAI22_X1 port map( A1 => n10081, A2 => n14604, B1 => n10695, B2 => 
                           n14616, ZN => n14566);
   U2138 : INV_X1 port map( A => n14566, ZN => n3434);
   U2139 : OAI22_X1 port map( A1 => n10081, A2 => n14573, B1 => n11099, B2 => 
                           n14616, ZN => n14567);
   U2140 : INV_X1 port map( A => n14567, ZN => n3402);
   U2141 : OAI22_X1 port map( A1 => n10081, A2 => n14610, B1 => n11069, B2 => 
                           n14616, ZN => n14568);
   U2142 : INV_X1 port map( A => n14568, ZN => n3370);
   U2143 : OAI22_X1 port map( A1 => n10078, A2 => n14610, B1 => n11052, B2 => 
                           n14606, ZN => n14569);
   U2144 : INV_X1 port map( A => n14569, ZN => n3373);
   U2145 : OAI22_X1 port map( A1 => n10082, A2 => n14610, B1 => n11068, B2 => 
                           n14618, ZN => n14570);
   U2146 : INV_X1 port map( A => n14570, ZN => n3369);
   U2147 : OAI22_X1 port map( A1 => n10083, A2 => n14610, B1 => n11067, B2 => 
                           n14597, ZN => n14571);
   U2148 : INV_X1 port map( A => n14571, ZN => n3368);
   U2149 : OAI22_X1 port map( A1 => n10086, A2 => n14619, B1 => n11034, B2 => 
                           n14603, ZN => n14572);
   U2150 : INV_X1 port map( A => n14572, ZN => n3333);
   U2151 : OAI22_X1 port map( A1 => n10086, A2 => n14573, B1 => n11094, B2 => 
                           n14603, ZN => n14574);
   U2152 : INV_X1 port map( A => n14574, ZN => n3397);
   U2153 : OAI22_X1 port map( A1 => n10084, A2 => n14594, B1 => n10330, B2 => 
                           n14614, ZN => n14575);
   U2154 : INV_X1 port map( A => n14575, ZN => n3495);
   U2155 : OAI22_X1 port map( A1 => n10085, A2 => n14610, B1 => n11065, B2 => 
                           n14583, ZN => n14576);
   U2156 : INV_X1 port map( A => n14576, ZN => n3366);
   U2157 : OAI22_X1 port map( A1 => n10083, A2 => n14594, B1 => n10331, B2 => 
                           n14597, ZN => n14577);
   U2158 : INV_X1 port map( A => n14577, ZN => n3496);
   U2159 : OAI22_X1 port map( A1 => n10082, A2 => n14594, B1 => n10332, B2 => 
                           n14618, ZN => n14578);
   U2160 : INV_X1 port map( A => n14578, ZN => n3497);
   U2161 : OAI22_X1 port map( A1 => n10086, A2 => n14610, B1 => n11064, B2 => 
                           n14603, ZN => n14579);
   U2162 : INV_X1 port map( A => n14579, ZN => n3365);
   U2163 : OAI22_X1 port map( A1 => n10087, A2 => n14610, B1 => n11063, B2 => 
                           n14580, ZN => n14581);
   U2164 : INV_X1 port map( A => n14581, ZN => n3364);
   U2165 : OAI22_X1 port map( A1 => n10090, A2 => n14610, B1 => n11060, B2 => 
                           n14612, ZN => n14582);
   U2166 : INV_X1 port map( A => n14582, ZN => n3361);
   U2167 : OAI22_X1 port map( A1 => n10085, A2 => n14619, B1 => n11035, B2 => 
                           n14583, ZN => n14584);
   U2168 : INV_X1 port map( A => n14584, ZN => n3334);
   U2169 : OAI22_X1 port map( A1 => n10077, A2 => n14594, B1 => n10337, B2 => 
                           n14608, ZN => n14585);
   U2170 : INV_X1 port map( A => n14585, ZN => n3502);
   U2171 : OAI22_X1 port map( A1 => n10081, A2 => n14594, B1 => n10333, B2 => 
                           n14616, ZN => n14586);
   U2172 : INV_X1 port map( A => n14586, ZN => n3498);
   U2173 : OAI22_X1 port map( A1 => n10080, A2 => n14619, B1 => n11019, B2 => 
                           n14588, ZN => n14587);
   U2174 : INV_X1 port map( A => n14587, ZN => n3339);
   U2175 : OAI22_X1 port map( A1 => n10080, A2 => n14594, B1 => n10334, B2 => 
                           n14588, ZN => n14589);
   U2176 : INV_X1 port map( A => n14589, ZN => n3499);
   U2177 : OAI22_X1 port map( A1 => n10079, A2 => n14619, B1 => n11020, B2 => 
                           n14601, ZN => n14590);
   U2178 : INV_X1 port map( A => n14590, ZN => n3340);
   U2179 : OAI22_X1 port map( A1 => n10079, A2 => n14591, B1 => n10668, B2 => 
                           n14601, ZN => n14592);
   U2180 : INV_X1 port map( A => n14592, ZN => n3532);
   U2181 : OAI22_X1 port map( A1 => n10079, A2 => n14594, B1 => n10335, B2 => 
                           n14601, ZN => n14593);
   U2182 : INV_X1 port map( A => n14593, ZN => n3500);
   U2183 : OAI22_X1 port map( A1 => n10078, A2 => n14594, B1 => n10336, B2 => 
                           n14606, ZN => n14595);
   U2184 : INV_X1 port map( A => n14595, ZN => n3501);
   U2185 : OAI22_X1 port map( A1 => n10077, A2 => n14610, B1 => n11053, B2 => 
                           n14608, ZN => n14596);
   U2186 : INV_X1 port map( A => n14596, ZN => n3374);
   U2187 : OAI22_X1 port map( A1 => n10083, A2 => n14619, B1 => n11037, B2 => 
                           n14597, ZN => n14598);
   U2188 : INV_X1 port map( A => n14598, ZN => n3336);
   U2189 : OAI22_X1 port map( A1 => n10086, A2 => n14599, B1 => n10720, B2 => 
                           n14603, ZN => n14600);
   U2190 : INV_X1 port map( A => n14600, ZN => n3461);
   U2191 : OAI22_X1 port map( A1 => n10079, A2 => n14610, B1 => n11051, B2 => 
                           n14601, ZN => n14602);
   U2192 : INV_X1 port map( A => n14602, ZN => n3372);
   U2193 : OAI22_X1 port map( A1 => n10086, A2 => n14604, B1 => n10690, B2 => 
                           n14603, ZN => n14605);
   U2194 : INV_X1 port map( A => n14605, ZN => n3429);
   U2195 : OAI22_X1 port map( A1 => n10078, A2 => n14619, B1 => n11021, B2 => 
                           n14606, ZN => n14607);
   U2196 : INV_X1 port map( A => n14607, ZN => n3341);
   U2197 : OAI22_X1 port map( A1 => n10077, A2 => n14619, B1 => n11022, B2 => 
                           n14608, ZN => n14609);
   U2198 : INV_X1 port map( A => n14609, ZN => n3342);
   U2199 : OAI22_X1 port map( A1 => n10084, A2 => n14610, B1 => n11066, B2 => 
                           n14614, ZN => n14611);
   U2200 : INV_X1 port map( A => n14611, ZN => n3367);
   U2201 : OAI22_X1 port map( A1 => n10090, A2 => n14619, B1 => n11030, B2 => 
                           n14612, ZN => n14613);
   U2202 : INV_X1 port map( A => n14613, ZN => n3329);
   U2203 : OAI22_X1 port map( A1 => n10084, A2 => n14619, B1 => n11036, B2 => 
                           n14614, ZN => n14615);
   U2204 : INV_X1 port map( A => n14615, ZN => n3335);
   U2205 : OAI22_X1 port map( A1 => n10081, A2 => n14619, B1 => n11039, B2 => 
                           n14616, ZN => n14617);
   U2206 : INV_X1 port map( A => n14617, ZN => n3338);
   U2207 : OAI22_X1 port map( A1 => n10082, A2 => n14619, B1 => n11038, B2 => 
                           n14618, ZN => n14620);
   U2208 : INV_X1 port map( A => n14620, ZN => n3337);
   U2209 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1),
                           ZN => n14632);
   U2210 : INV_X1 port map( A => ADD_WR(3), ZN => n14621);
   U2211 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => n14621, ZN => 
                           n14628);
   U2212 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n14628, ZN => n14626);
   U2213 : NAND2_X1 port map( A1 => n14632, A2 => n14626, ZN => n3987);
   U2214 : INV_X1 port map( A => ADD_WR(0), ZN => n14622);
   U2215 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n14622, ZN
                           => n14633);
   U2216 : NAND2_X1 port map( A1 => n14626, A2 => n14633, ZN => n3991);
   U2217 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n14622, ZN => n14623);
   U2218 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n14623, ZN => n14634);
   U2219 : NAND2_X1 port map( A1 => n14626, A2 => n14634, ZN => n3994);
   U2220 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n14624);
   U2221 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n14624, ZN => n14635);
   U2222 : NAND2_X1 port map( A1 => n14626, A2 => n14635, ZN => n3997);
   U2223 : INV_X1 port map( A => ADD_WR(2), ZN => n14625);
   U2224 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n14625, ZN
                           => n14636);
   U2225 : NAND2_X1 port map( A1 => n14626, A2 => n14636, ZN => n4000);
   U2226 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n14622, A3 => n14625, ZN =>
                           n14637);
   U2227 : NAND2_X1 port map( A1 => n14626, A2 => n14637, ZN => n4005);
   U2228 : NOR2_X1 port map( A1 => n14625, A2 => n14623, ZN => n14638);
   U2229 : NAND2_X1 port map( A1 => n14626, A2 => n14638, ZN => n4009);
   U2230 : NOR2_X1 port map( A1 => n14625, A2 => n14624, ZN => n14640);
   U2231 : NAND2_X1 port map( A1 => n14626, A2 => n14640, ZN => n4034);
   U2232 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(3), ZN => 
                           n14630);
   U2233 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n14630, ZN => n14627);
   U2234 : NAND2_X1 port map( A1 => n14632, A2 => n14627, ZN => n4039);
   U2235 : NAND2_X1 port map( A1 => n14633, A2 => n14627, ZN => n4043);
   U2236 : NAND2_X1 port map( A1 => n14634, A2 => n14627, ZN => n4046);
   U2237 : NAND2_X1 port map( A1 => n14635, A2 => n14627, ZN => n4049);
   U2238 : NAND2_X1 port map( A1 => n14636, A2 => n14627, ZN => n4052);
   U2239 : NAND2_X1 port map( A1 => n14637, A2 => n14627, ZN => n4055);
   U2240 : NAND2_X1 port map( A1 => n14638, A2 => n14627, ZN => n4059);
   U2241 : NAND2_X1 port map( A1 => n14640, A2 => n14627, ZN => n4063);
   U2242 : INV_X1 port map( A => ADD_WR(4), ZN => n14631);
   U2243 : NOR2_X1 port map( A1 => n14631, A2 => n14628, ZN => n14629);
   U2244 : NAND2_X1 port map( A1 => n14632, A2 => n14629, ZN => n4067);
   U2245 : NAND2_X1 port map( A1 => n14633, A2 => n14629, ZN => n4071);
   U2246 : NAND2_X1 port map( A1 => n14634, A2 => n14629, ZN => n4075);
   U2247 : NAND2_X1 port map( A1 => n14635, A2 => n14629, ZN => n4079);
   U2248 : NAND2_X1 port map( A1 => n14636, A2 => n14629, ZN => n4090);
   U2249 : NAND2_X1 port map( A1 => n14637, A2 => n14629, ZN => n4094);
   U2250 : NAND2_X1 port map( A1 => n14638, A2 => n14629, ZN => n4097);
   U2251 : NAND2_X1 port map( A1 => n14640, A2 => n14629, ZN => n4102);
   U2252 : NOR2_X1 port map( A1 => n14631, A2 => n14630, ZN => n14639);
   U2253 : NAND2_X1 port map( A1 => n14632, A2 => n14639, ZN => n4110);
   U2254 : NAND2_X1 port map( A1 => n14633, A2 => n14639, ZN => n4115);
   U2255 : NAND2_X1 port map( A1 => n14634, A2 => n14639, ZN => n4120);
   U2256 : NAND2_X1 port map( A1 => n14635, A2 => n14639, ZN => n4125);
   U2257 : NAND2_X1 port map( A1 => n14636, A2 => n14639, ZN => n4130);
   U2258 : NAND2_X1 port map( A1 => n14637, A2 => n14639, ZN => n4135);
   U2259 : NAND2_X1 port map( A1 => n14638, A2 => n14639, ZN => n4140);
   U2260 : NAND2_X1 port map( A1 => n14640, A2 => n14639, ZN => n4177);
   U2261 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n3583, ZN => n14650);
   U2262 : INV_X1 port map( A => n3587, ZN => n14643);
   U2263 : NOR2_X1 port map( A1 => n14650, A2 => n14643, ZN => n4906);
   U2264 : INV_X1 port map( A => n3586, ZN => n14648);
   U2265 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n14645)
                           ;
   U2266 : NOR2_X1 port map( A1 => n14648, A2 => n14645, ZN => n4754);
   U2267 : INV_X1 port map( A => n3588, ZN => n14641);
   U2268 : NOR2_X1 port map( A1 => n14645, A2 => n14641, ZN => n4803);
   U2269 : INV_X1 port map( A => n3585, ZN => n14642);
   U2270 : NOR2_X1 port map( A1 => n14645, A2 => n14642, ZN => n4710);
   U2271 : NOR2_X1 port map( A1 => n14650, A2 => n14641, ZN => n4882);
   U2272 : INV_X1 port map( A => n3590, ZN => n14647);
   U2273 : NOR2_X1 port map( A1 => n14645, A2 => n14647, ZN => n4621);
   U2274 : INV_X1 port map( A => n3591, ZN => n14649);
   U2275 : NOR2_X1 port map( A1 => n14645, A2 => n14649, ZN => n4825);
   U2276 : NOR2_X1 port map( A1 => n14650, A2 => n14642, ZN => n4905);
   U2277 : INV_X1 port map( A => n3589, ZN => n14644);
   U2278 : NOR2_X1 port map( A1 => n14650, A2 => n14644, ZN => n4856);
   U2279 : NOR2_X1 port map( A1 => n14643, A2 => n14645, ZN => n4881);
   U2280 : NOR2_X1 port map( A1 => n14645, A2 => n14644, ZN => n4442);
   U2281 : INV_X1 port map( A => n3584, ZN => n14646);
   U2282 : NOR2_X1 port map( A1 => n14645, A2 => n14646, ZN => n4855);
   U2283 : NOR2_X1 port map( A1 => n14650, A2 => n14646, ZN => n4883);
   U2284 : NOR2_X1 port map( A1 => n14650, A2 => n14647, ZN => n4920);
   U2285 : NOR2_X1 port map( A1 => n14650, A2 => n14648, ZN => n4876);
   U2286 : NOR2_X1 port map( A1 => n14650, A2 => n14649, ZN => n4804);
   U2287 : AOI22_X1 port map( A1 => n9398, A2 => n10070, B1 => n9366, B2 => 
                           n11188, ZN => n14654);
   U2288 : AOI22_X1 port map( A1 => n9206, A2 => n10068, B1 => n9302, B2 => 
                           n10063, ZN => n14653);
   U2289 : AOI22_X1 port map( A1 => n9142, A2 => n11190, B1 => n9430, B2 => 
                           n11187, ZN => n14652);
   U2290 : AOI22_X1 port map( A1 => n9078, A2 => n10069, B1 => n9462, B2 => 
                           n10066, ZN => n14651);
   U2291 : NAND4_X1 port map( A1 => n14654, A2 => n14653, A3 => n14652, A4 => 
                           n14651, ZN => n14660);
   U2292 : AOI22_X1 port map( A1 => n9174, A2 => n10065, B1 => n9110, B2 => 
                           n11189, ZN => n14658);
   U2293 : AOI22_X1 port map( A1 => n9494, A2 => n10055, B1 => n9046, B2 => 
                           n11191, ZN => n14657);
   U2294 : AOI22_X1 port map( A1 => n9526, A2 => n10062, B1 => n9238, B2 => 
                           n10064, ZN => n14656);
   U2295 : AOI22_X1 port map( A1 => n9270, A2 => n10060, B1 => n9334, B2 => 
                           n11186, ZN => n14655);
   U2296 : NAND4_X1 port map( A1 => n14658, A2 => n14657, A3 => n14656, A4 => 
                           n14655, ZN => n14659);
   U2297 : NOR2_X1 port map( A1 => n14660, A2 => n14659, ZN => n14672);
   U2298 : NOR3_X1 port map( A1 => n11265, A2 => n11266, A3 => n15182, ZN => 
                           n15112);
   U2299 : CLKBUF_X1 port map( A => n15112, Z => n15157);
   U2300 : AOI22_X1 port map( A1 => n10038, A2 => n11227, B1 => n10006, B2 => 
                           n11181, ZN => n14664);
   U2301 : AOI22_X1 port map( A1 => n9974, A2 => n11226, B1 => n9878, B2 => 
                           n11180, ZN => n14663);
   U2302 : AOI22_X1 port map( A1 => n9910, A2 => n11182, B1 => n9846, B2 => 
                           n11184, ZN => n14662);
   U2303 : AOI22_X1 port map( A1 => n9814, A2 => n11183, B1 => n9942, B2 => 
                           n11185, ZN => n14661);
   U2304 : NAND4_X1 port map( A1 => n14664, A2 => n14663, A3 => n14662, A4 => 
                           n14661, ZN => n14670);
   U2305 : NOR3_X1 port map( A1 => n11266, A2 => n11192, A3 => n15182, ZN => 
                           n14890);
   U2306 : CLKBUF_X1 port map( A => n14890, Z => n15358);
   U2307 : CLKBUF_X1 port map( A => n11226, Z => n15325);
   U2308 : AOI22_X1 port map( A1 => n15325, A2 => n9718, B1 => n9622, B2 => 
                           n11177, ZN => n14668);
   U2309 : AOI22_X1 port map( A1 => n9750, A2 => n11176, B1 => n9558, B2 => 
                           n11179, ZN => n14667);
   U2310 : CLKBUF_X1 port map( A => n11227, Z => n15352);
   U2311 : AOI22_X1 port map( A1 => n15352, A2 => n9782, B1 => n11184, B2 => 
                           n9590, ZN => n14666);
   U2312 : AOI22_X1 port map( A1 => n11185, A2 => n9686, B1 => n9654, B2 => 
                           n11178, ZN => n14665);
   U2313 : NAND4_X1 port map( A1 => n14668, A2 => n14667, A3 => n14666, A4 => 
                           n14665, ZN => n14669);
   U2314 : AOI22_X1 port map( A1 => n15157, A2 => n14670, B1 => n15358, B2 => 
                           n14669, ZN => n14671);
   U2315 : OAI21_X1 port map( B1 => n15182, B2 => n14672, A => n14671, ZN => 
                           OUT2(31));
   U2316 : AOI22_X1 port map( A1 => n10062, A2 => n9525, B1 => n9205, B2 => 
                           n11173, ZN => n14676);
   U2317 : AOI22_X1 port map( A1 => n10055, A2 => n9493, B1 => n11190, B2 => 
                           n9141, ZN => n14675);
   U2318 : AOI22_X1 port map( A1 => n11191, A2 => n9045, B1 => n11189, B2 => 
                           n9109, ZN => n14674);
   U2319 : AOI22_X1 port map( A1 => n9077, A2 => n11174, B1 => n9397, B2 => 
                           n11175, ZN => n14673);
   U2320 : NAND4_X1 port map( A1 => n14676, A2 => n14675, A3 => n14674, A4 => 
                           n14673, ZN => n14682);
   U2321 : AOI22_X1 port map( A1 => n11187, A2 => n9429, B1 => n9173, B2 => 
                           n11172, ZN => n14680);
   U2322 : AOI22_X1 port map( A1 => n10060, A2 => n9269, B1 => n11188, B2 => 
                           n9365, ZN => n14679);
   U2323 : AOI22_X1 port map( A1 => n10064, A2 => n9237, B1 => n9333, B2 => 
                           n10056, ZN => n14678);
   U2324 : AOI22_X1 port map( A1 => n10063, A2 => n9301, B1 => n10066, B2 => 
                           n9461, ZN => n14677);
   U2325 : NAND4_X1 port map( A1 => n14680, A2 => n14679, A3 => n14678, A4 => 
                           n14677, ZN => n14681);
   U2326 : NOR2_X1 port map( A1 => n14682, A2 => n14681, ZN => n14694);
   U2327 : AOI22_X1 port map( A1 => n11177, A2 => n9877, B1 => n9845, B2 => 
                           n11171, ZN => n14686);
   U2328 : AOI22_X1 port map( A1 => n11181, A2 => n10005, B1 => n11182, B2 => 
                           n9909, ZN => n14685);
   U2329 : AOI22_X1 port map( A1 => n15325, A2 => n9973, B1 => n9941, B2 => 
                           n11170, ZN => n14684);
   U2330 : AOI22_X1 port map( A1 => n11227, A2 => n10037, B1 => n11179, B2 => 
                           n9813, ZN => n14683);
   U2331 : NAND4_X1 port map( A1 => n14686, A2 => n14685, A3 => n14684, A4 => 
                           n14683, ZN => n14692);
   U2332 : AOI22_X1 port map( A1 => n11185, A2 => n9685, B1 => n9749, B2 => 
                           n11169, ZN => n14690);
   U2333 : AOI22_X1 port map( A1 => n11184, A2 => n9589, B1 => n11178, B2 => 
                           n9653, ZN => n14689);
   U2334 : AOI22_X1 port map( A1 => n11226, A2 => n9717, B1 => n11183, B2 => 
                           n9557, ZN => n14688);
   U2335 : AOI22_X1 port map( A1 => n15352, A2 => n9781, B1 => n11177, B2 => 
                           n9621, ZN => n14687);
   U2336 : NAND4_X1 port map( A1 => n14690, A2 => n14689, A3 => n14688, A4 => 
                           n14687, ZN => n14691);
   U2337 : AOI22_X1 port map( A1 => n15157, A2 => n14692, B1 => n15358, B2 => 
                           n14691, ZN => n14693);
   U2338 : OAI21_X1 port map( B1 => n15182, B2 => n14694, A => n14693, ZN => 
                           OUT2(30));
   U2339 : AOI22_X1 port map( A1 => n11189, A2 => n9108, B1 => n9460, B2 => 
                           n11168, ZN => n14698);
   U2340 : AOI22_X1 port map( A1 => n10055, A2 => n9492, B1 => n9524, B2 => 
                           n11167, ZN => n14697);
   U2341 : AOI22_X1 port map( A1 => n11186, A2 => n9332, B1 => n9300, B2 => 
                           n11165, ZN => n14696);
   U2342 : AOI22_X1 port map( A1 => n10060, A2 => n9268, B1 => n9236, B2 => 
                           n11166, ZN => n14695);
   U2343 : NAND4_X1 port map( A1 => n14698, A2 => n14697, A3 => n14696, A4 => 
                           n14695, ZN => n14704);
   U2344 : AOI22_X1 port map( A1 => n11190, A2 => n9140, B1 => n9364, B2 => 
                           n10058, ZN => n14702);
   U2345 : AOI22_X1 port map( A1 => n11173, A2 => n9204, B1 => n11175, B2 => 
                           n9396, ZN => n14701);
   U2346 : AOI22_X1 port map( A1 => n11174, A2 => n9076, B1 => n9428, B2 => 
                           n10057, ZN => n14700);
   U2347 : AOI22_X1 port map( A1 => n10065, A2 => n9172, B1 => n9044, B2 => 
                           n10067, ZN => n14699);
   U2348 : NAND4_X1 port map( A1 => n14702, A2 => n14701, A3 => n14700, A4 => 
                           n14699, ZN => n14703);
   U2349 : NOR2_X1 port map( A1 => n14704, A2 => n14703, ZN => n14716);
   U2350 : AOI22_X1 port map( A1 => n11178, A2 => n9908, B1 => n9876, B2 => 
                           n11164, ZN => n14708);
   U2351 : AOI22_X1 port map( A1 => n11176, A2 => n10004, B1 => n11170, B2 => 
                           n9940, ZN => n14707);
   U2352 : AOI22_X1 port map( A1 => n11227, A2 => n10036, B1 => n15325, B2 => 
                           n9972, ZN => n14706);
   U2353 : AOI22_X1 port map( A1 => n11184, A2 => n9844, B1 => n9812, B2 => 
                           n11163, ZN => n14705);
   U2354 : NAND4_X1 port map( A1 => n14708, A2 => n14707, A3 => n14706, A4 => 
                           n14705, ZN => n14714);
   U2355 : AOI22_X1 port map( A1 => n11179, A2 => n9556, B1 => n11169, B2 => 
                           n9748, ZN => n14712);
   U2356 : AOI22_X1 port map( A1 => n15352, A2 => n9780, B1 => n11226, B2 => 
                           n9716, ZN => n14711);
   U2357 : AOI22_X1 port map( A1 => n11184, A2 => n9588, B1 => n11178, B2 => 
                           n9652, ZN => n14710);
   U2358 : AOI22_X1 port map( A1 => n11177, A2 => n9620, B1 => n11170, B2 => 
                           n9684, ZN => n14709);
   U2359 : NAND4_X1 port map( A1 => n14712, A2 => n14711, A3 => n14710, A4 => 
                           n14709, ZN => n14713);
   U2360 : AOI22_X1 port map( A1 => n15157, A2 => n14714, B1 => n15358, B2 => 
                           n14713, ZN => n14715);
   U2361 : OAI21_X1 port map( B1 => n15182, B2 => n14716, A => n14715, ZN => 
                           OUT2(29));
   U2362 : AOI22_X1 port map( A1 => n11165, A2 => n9299, B1 => n9139, B2 => 
                           n10061, ZN => n14720);
   U2363 : AOI22_X1 port map( A1 => n11191, A2 => n9043, B1 => n11173, B2 => 
                           n9203, ZN => n14719);
   U2364 : AOI22_X1 port map( A1 => n10070, A2 => n9395, B1 => n11167, B2 => 
                           n9523, ZN => n14718);
   U2365 : AOI22_X1 port map( A1 => n11186, A2 => n9331, B1 => n10069, B2 => 
                           n9075, ZN => n14717);
   U2366 : NAND4_X1 port map( A1 => n14720, A2 => n14719, A3 => n14718, A4 => 
                           n14717, ZN => n14726);
   U2367 : AOI22_X1 port map( A1 => n11189, A2 => n9107, B1 => n9491, B2 => 
                           n11162, ZN => n14724);
   U2368 : AOI22_X1 port map( A1 => n11172, A2 => n9171, B1 => n11168, B2 => 
                           n9459, ZN => n14723);
   U2369 : AOI22_X1 port map( A1 => n11188, A2 => n9363, B1 => n11166, B2 => 
                           n9235, ZN => n14722);
   U2370 : AOI22_X1 port map( A1 => n10060, A2 => n9267, B1 => n11187, B2 => 
                           n9427, ZN => n14721);
   U2371 : NAND4_X1 port map( A1 => n14724, A2 => n14723, A3 => n14722, A4 => 
                           n14721, ZN => n14725);
   U2372 : NOR2_X1 port map( A1 => n14726, A2 => n14725, ZN => n14738);
   U2373 : AOI22_X1 port map( A1 => n11185, A2 => n9939, B1 => n11177, B2 => 
                           n9875, ZN => n14730);
   U2374 : AOI22_X1 port map( A1 => n11227, A2 => n10035, B1 => n11184, B2 => 
                           n9843, ZN => n14729);
   U2375 : AOI22_X1 port map( A1 => n11226, A2 => n9971, B1 => n11183, B2 => 
                           n9811, ZN => n14728);
   U2376 : AOI22_X1 port map( A1 => n11181, A2 => n10003, B1 => n9907, B2 => 
                           n11161, ZN => n14727);
   U2377 : NAND4_X1 port map( A1 => n14730, A2 => n14729, A3 => n14728, A4 => 
                           n14727, ZN => n14736);
   U2378 : AOI22_X1 port map( A1 => n11183, A2 => n9555, B1 => n11177, B2 => 
                           n9619, ZN => n14734);
   U2379 : AOI22_X1 port map( A1 => n15325, A2 => n9715, B1 => n11170, B2 => 
                           n9683, ZN => n14733);
   U2380 : AOI22_X1 port map( A1 => n11176, A2 => n9747, B1 => n11178, B2 => 
                           n9651, ZN => n14732);
   U2381 : AOI22_X1 port map( A1 => n15352, A2 => n9779, B1 => n11184, B2 => 
                           n9587, ZN => n14731);
   U2382 : NAND4_X1 port map( A1 => n14734, A2 => n14733, A3 => n14732, A4 => 
                           n14731, ZN => n14735);
   U2383 : AOI22_X1 port map( A1 => n15157, A2 => n14736, B1 => n15358, B2 => 
                           n14735, ZN => n14737);
   U2384 : OAI21_X1 port map( B1 => n15182, B2 => n14738, A => n14737, ZN => 
                           OUT2(28));
   U2385 : AOI22_X1 port map( A1 => n11190, A2 => n9138, B1 => n10067, B2 => 
                           n9042, ZN => n14742);
   U2386 : AOI22_X1 port map( A1 => n11186, A2 => n9330, B1 => n11175, B2 => 
                           n9394, ZN => n14741);
   U2387 : AOI22_X1 port map( A1 => n11187, A2 => n9426, B1 => n11165, B2 => 
                           n9298, ZN => n14740);
   U2388 : AOI22_X1 port map( A1 => n11189, A2 => n9106, B1 => n11173, B2 => 
                           n9202, ZN => n14739);
   U2389 : NAND4_X1 port map( A1 => n14742, A2 => n14741, A3 => n14740, A4 => 
                           n14739, ZN => n14748);
   U2390 : AOI22_X1 port map( A1 => n10060, A2 => n9266, B1 => n11162, B2 => 
                           n9490, ZN => n14746);
   U2391 : AOI22_X1 port map( A1 => n10065, A2 => n9170, B1 => n11167, B2 => 
                           n9522, ZN => n14745);
   U2392 : AOI22_X1 port map( A1 => n11174, A2 => n9074, B1 => n11166, B2 => 
                           n9234, ZN => n14744);
   U2393 : AOI22_X1 port map( A1 => n10058, A2 => n9362, B1 => n11168, B2 => 
                           n9458, ZN => n14743);
   U2394 : NAND4_X1 port map( A1 => n14746, A2 => n14745, A3 => n14744, A4 => 
                           n14743, ZN => n14747);
   U2395 : NOR2_X1 port map( A1 => n14748, A2 => n14747, ZN => n14760);
   U2396 : AOI22_X1 port map( A1 => n11177, A2 => n9874, B1 => n11176, B2 => 
                           n10002, ZN => n14752);
   U2397 : AOI22_X1 port map( A1 => n15325, A2 => n9970, B1 => n11178, B2 => 
                           n9906, ZN => n14751);
   U2398 : AOI22_X1 port map( A1 => n11179, A2 => n9810, B1 => n11170, B2 => 
                           n9938, ZN => n14750);
   U2399 : AOI22_X1 port map( A1 => n11227, A2 => n10034, B1 => n9842, B2 => 
                           n11160, ZN => n14749);
   U2400 : NAND4_X1 port map( A1 => n14752, A2 => n14751, A3 => n14750, A4 => 
                           n14749, ZN => n14758);
   U2401 : AOI22_X1 port map( A1 => n11226, A2 => n9714, B1 => n11179, B2 => 
                           n9554, ZN => n14756);
   U2402 : AOI22_X1 port map( A1 => n11176, A2 => n9746, B1 => n11160, B2 => 
                           n9586, ZN => n14755);
   U2403 : AOI22_X1 port map( A1 => n11178, A2 => n9650, B1 => n11170, B2 => 
                           n9682, ZN => n14754);
   U2404 : AOI22_X1 port map( A1 => n15352, A2 => n9778, B1 => n11177, B2 => 
                           n9618, ZN => n14753);
   U2405 : NAND4_X1 port map( A1 => n14756, A2 => n14755, A3 => n14754, A4 => 
                           n14753, ZN => n14757);
   U2406 : AOI22_X1 port map( A1 => n15157, A2 => n14758, B1 => n14890, B2 => 
                           n14757, ZN => n14759);
   U2407 : OAI21_X1 port map( B1 => n15182, B2 => n14760, A => n14759, ZN => 
                           OUT2(27));
   U2408 : AOI22_X1 port map( A1 => n11190, A2 => n9137, B1 => n11165, B2 => 
                           n9297, ZN => n14764);
   U2409 : AOI22_X1 port map( A1 => n11189, A2 => n9105, B1 => n10060, B2 => 
                           n9265, ZN => n14763);
   U2410 : AOI22_X1 port map( A1 => n10056, A2 => n9329, B1 => n10058, B2 => 
                           n9361, ZN => n14762);
   U2411 : AOI22_X1 port map( A1 => n11175, A2 => n9393, B1 => n10057, B2 => 
                           n9425, ZN => n14761);
   U2412 : NAND4_X1 port map( A1 => n14764, A2 => n14763, A3 => n14762, A4 => 
                           n14761, ZN => n14770);
   U2413 : AOI22_X1 port map( A1 => n11167, A2 => n9521, B1 => n11168, B2 => 
                           n9457, ZN => n14768);
   U2414 : AOI22_X1 port map( A1 => n10055, A2 => n9489, B1 => n11173, B2 => 
                           n9201, ZN => n14767);
   U2415 : AOI22_X1 port map( A1 => n11191, A2 => n9041, B1 => n11172, B2 => 
                           n9169, ZN => n14766);
   U2416 : AOI22_X1 port map( A1 => n11174, A2 => n9073, B1 => n11166, B2 => 
                           n9233, ZN => n14765);
   U2417 : NAND4_X1 port map( A1 => n14768, A2 => n14767, A3 => n14766, A4 => 
                           n14765, ZN => n14769);
   U2418 : NOR2_X1 port map( A1 => n14770, A2 => n14769, ZN => n14782);
   U2419 : AOI22_X1 port map( A1 => n11226, A2 => n9969, B1 => n11177, B2 => 
                           n9873, ZN => n14774);
   U2420 : AOI22_X1 port map( A1 => n11227, A2 => n10033, B1 => n11163, B2 => 
                           n9809, ZN => n14773);
   U2421 : AOI22_X1 port map( A1 => n11178, A2 => n9905, B1 => n11169, B2 => 
                           n10001, ZN => n14772);
   U2422 : AOI22_X1 port map( A1 => n11171, A2 => n9841, B1 => n9937, B2 => 
                           n11159, ZN => n14771);
   U2423 : NAND4_X1 port map( A1 => n14774, A2 => n14773, A3 => n14772, A4 => 
                           n14771, ZN => n14780);
   U2424 : AOI22_X1 port map( A1 => n11177, A2 => n9617, B1 => n11159, B2 => 
                           n9681, ZN => n14778);
   U2425 : AOI22_X1 port map( A1 => n11176, A2 => n9745, B1 => n9777, B2 => 
                           n11158, ZN => n14777);
   U2426 : AOI22_X1 port map( A1 => n11161, A2 => n9649, B1 => n11160, B2 => 
                           n9585, ZN => n14776);
   U2427 : AOI22_X1 port map( A1 => n15325, A2 => n9713, B1 => n11163, B2 => 
                           n9553, ZN => n14775);
   U2428 : NAND4_X1 port map( A1 => n14778, A2 => n14777, A3 => n14776, A4 => 
                           n14775, ZN => n14779);
   U2429 : AOI22_X1 port map( A1 => n15157, A2 => n14780, B1 => n14890, B2 => 
                           n14779, ZN => n14781);
   U2430 : OAI21_X1 port map( B1 => n15182, B2 => n14782, A => n14781, ZN => 
                           OUT2(26));
   U2431 : AOI22_X1 port map( A1 => n11175, A2 => n9392, B1 => n10061, B2 => 
                           n9136, ZN => n14786);
   U2432 : AOI22_X1 port map( A1 => n11189, A2 => n9104, B1 => n10069, B2 => 
                           n9072, ZN => n14785);
   U2433 : AOI22_X1 port map( A1 => n10055, A2 => n9488, B1 => n9264, B2 => 
                           n11157, ZN => n14784);
   U2434 : AOI22_X1 port map( A1 => n11191, A2 => n9040, B1 => n11188, B2 => 
                           n9360, ZN => n14783);
   U2435 : NAND4_X1 port map( A1 => n14786, A2 => n14785, A3 => n14784, A4 => 
                           n14783, ZN => n14792);
   U2436 : AOI22_X1 port map( A1 => n11187, A2 => n9424, B1 => n11168, B2 => 
                           n9456, ZN => n14790);
   U2437 : AOI22_X1 port map( A1 => n10065, A2 => n9168, B1 => n11186, B2 => 
                           n9328, ZN => n14789);
   U2438 : AOI22_X1 port map( A1 => n11167, A2 => n9520, B1 => n11166, B2 => 
                           n9232, ZN => n14788);
   U2439 : AOI22_X1 port map( A1 => n11173, A2 => n9200, B1 => n11165, B2 => 
                           n9296, ZN => n14787);
   U2440 : NAND4_X1 port map( A1 => n14790, A2 => n14789, A3 => n14788, A4 => 
                           n14787, ZN => n14791);
   U2441 : NOR2_X1 port map( A1 => n14792, A2 => n14791, ZN => n14804);
   U2442 : AOI22_X1 port map( A1 => n11181, A2 => n10000, B1 => n11163, B2 => 
                           n9808, ZN => n14796);
   U2443 : AOI22_X1 port map( A1 => n11184, A2 => n9840, B1 => n11161, B2 => 
                           n9904, ZN => n14795);
   U2444 : AOI22_X1 port map( A1 => n15352, A2 => n10032, B1 => n11185, B2 => 
                           n9936, ZN => n14794);
   U2445 : AOI22_X1 port map( A1 => n15325, A2 => n9968, B1 => n11180, B2 => 
                           n9872, ZN => n14793);
   U2446 : NAND4_X1 port map( A1 => n14796, A2 => n14795, A3 => n14794, A4 => 
                           n14793, ZN => n14802);
   U2447 : AOI22_X1 port map( A1 => n11180, A2 => n9616, B1 => n11176, B2 => 
                           n9744, ZN => n14800);
   U2448 : AOI22_X1 port map( A1 => n11226, A2 => n9712, B1 => n11163, B2 => 
                           n9552, ZN => n14799);
   U2449 : AOI22_X1 port map( A1 => n15352, A2 => n9776, B1 => n11171, B2 => 
                           n9584, ZN => n14798);
   U2450 : AOI22_X1 port map( A1 => n11178, A2 => n9648, B1 => n11159, B2 => 
                           n9680, ZN => n14797);
   U2451 : NAND4_X1 port map( A1 => n14800, A2 => n14799, A3 => n14798, A4 => 
                           n14797, ZN => n14801);
   U2452 : AOI22_X1 port map( A1 => n15157, A2 => n14802, B1 => n14890, B2 => 
                           n14801, ZN => n14803);
   U2453 : OAI21_X1 port map( B1 => n15182, B2 => n14804, A => n14803, ZN => 
                           OUT2(25));
   U2454 : AOI22_X1 port map( A1 => n10069, A2 => n9071, B1 => n11162, B2 => 
                           n9487, ZN => n14808);
   U2455 : AOI22_X1 port map( A1 => n10065, A2 => n9167, B1 => n10067, B2 => 
                           n9039, ZN => n14807);
   U2456 : AOI22_X1 port map( A1 => n11186, A2 => n9327, B1 => n11166, B2 => 
                           n9231, ZN => n14806);
   U2457 : AOI22_X1 port map( A1 => n11187, A2 => n9423, B1 => n10061, B2 => 
                           n9135, ZN => n14805);
   U2458 : NAND4_X1 port map( A1 => n14808, A2 => n14807, A3 => n14806, A4 => 
                           n14805, ZN => n14814);
   U2459 : AOI22_X1 port map( A1 => n11189, A2 => n9103, B1 => n11175, B2 => 
                           n9391, ZN => n14812);
   U2460 : AOI22_X1 port map( A1 => n11173, A2 => n9199, B1 => n11165, B2 => 
                           n9295, ZN => n14811);
   U2461 : AOI22_X1 port map( A1 => n10060, A2 => n9263, B1 => n11167, B2 => 
                           n9519, ZN => n14810);
   U2462 : AOI22_X1 port map( A1 => n11188, A2 => n9359, B1 => n11168, B2 => 
                           n9455, ZN => n14809);
   U2463 : NAND4_X1 port map( A1 => n14812, A2 => n14811, A3 => n14810, A4 => 
                           n14809, ZN => n14813);
   U2464 : NOR2_X1 port map( A1 => n14814, A2 => n14813, ZN => n14826);
   U2465 : AOI22_X1 port map( A1 => n11170, A2 => n9935, B1 => n11158, B2 => 
                           n10031, ZN => n14818);
   U2466 : AOI22_X1 port map( A1 => n11226, A2 => n9967, B1 => n11164, B2 => 
                           n9871, ZN => n14817);
   U2467 : AOI22_X1 port map( A1 => n11163, A2 => n9807, B1 => n11160, B2 => 
                           n9839, ZN => n14816);
   U2468 : AOI22_X1 port map( A1 => n11176, A2 => n9999, B1 => n11178, B2 => 
                           n9903, ZN => n14815);
   U2469 : NAND4_X1 port map( A1 => n14818, A2 => n14817, A3 => n14816, A4 => 
                           n14815, ZN => n14824);
   U2470 : AOI22_X1 port map( A1 => n11182, A2 => n9647, B1 => n11184, B2 => 
                           n9583, ZN => n14822);
   U2471 : AOI22_X1 port map( A1 => n11176, A2 => n9743, B1 => n9711, B2 => 
                           n11156, ZN => n14821);
   U2472 : AOI22_X1 port map( A1 => n11177, A2 => n9615, B1 => n11163, B2 => 
                           n9551, ZN => n14820);
   U2473 : AOI22_X1 port map( A1 => n15352, A2 => n9775, B1 => n11170, B2 => 
                           n9679, ZN => n14819);
   U2474 : NAND4_X1 port map( A1 => n14822, A2 => n14821, A3 => n14820, A4 => 
                           n14819, ZN => n14823);
   U2475 : AOI22_X1 port map( A1 => n15157, A2 => n14824, B1 => n14890, B2 => 
                           n14823, ZN => n14825);
   U2476 : OAI21_X1 port map( B1 => n15182, B2 => n14826, A => n14825, ZN => 
                           OUT2(24));
   U2477 : AOI22_X1 port map( A1 => n11188, A2 => n9358, B1 => n11168, B2 => 
                           n9454, ZN => n14830);
   U2478 : AOI22_X1 port map( A1 => n11187, A2 => n9422, B1 => n11165, B2 => 
                           n9294, ZN => n14829);
   U2479 : AOI22_X1 port map( A1 => n10065, A2 => n9166, B1 => n11166, B2 => 
                           n9230, ZN => n14828);
   U2480 : AOI22_X1 port map( A1 => n11174, A2 => n9070, B1 => n11175, B2 => 
                           n9390, ZN => n14827);
   U2481 : NAND4_X1 port map( A1 => n14830, A2 => n14829, A3 => n14828, A4 => 
                           n14827, ZN => n14836);
   U2482 : AOI22_X1 port map( A1 => n11173, A2 => n9198, B1 => n11167, B2 => 
                           n9518, ZN => n14834);
   U2483 : AOI22_X1 port map( A1 => n10060, A2 => n9262, B1 => n11162, B2 => 
                           n9486, ZN => n14833);
   U2484 : AOI22_X1 port map( A1 => n11191, A2 => n9038, B1 => n11189, B2 => 
                           n9102, ZN => n14832);
   U2485 : AOI22_X1 port map( A1 => n11186, A2 => n9326, B1 => n11190, B2 => 
                           n9134, ZN => n14831);
   U2486 : NAND4_X1 port map( A1 => n14834, A2 => n14833, A3 => n14832, A4 => 
                           n14831, ZN => n14835);
   U2487 : NOR2_X1 port map( A1 => n14836, A2 => n14835, ZN => n14848);
   U2488 : AOI22_X1 port map( A1 => n11159, A2 => n9934, B1 => n11158, B2 => 
                           n10030, ZN => n14840);
   U2489 : AOI22_X1 port map( A1 => n15325, A2 => n9966, B1 => n11163, B2 => 
                           n9806, ZN => n14839);
   U2490 : AOI22_X1 port map( A1 => n11178, A2 => n9902, B1 => n11160, B2 => 
                           n9838, ZN => n14838);
   U2491 : AOI22_X1 port map( A1 => n11177, A2 => n9870, B1 => n11176, B2 => 
                           n9998, ZN => n14837);
   U2492 : NAND4_X1 port map( A1 => n14840, A2 => n14839, A3 => n14838, A4 => 
                           n14837, ZN => n14846);
   U2493 : AOI22_X1 port map( A1 => n11170, A2 => n9678, B1 => n11164, B2 => 
                           n9614, ZN => n14844);
   U2494 : AOI22_X1 port map( A1 => n11227, A2 => n9774, B1 => n15325, B2 => 
                           n9710, ZN => n14843);
   U2495 : AOI22_X1 port map( A1 => n11178, A2 => n9646, B1 => n11160, B2 => 
                           n9582, ZN => n14842);
   U2496 : AOI22_X1 port map( A1 => n11176, A2 => n9742, B1 => n11163, B2 => 
                           n9550, ZN => n14841);
   U2497 : NAND4_X1 port map( A1 => n14844, A2 => n14843, A3 => n14842, A4 => 
                           n14841, ZN => n14845);
   U2498 : AOI22_X1 port map( A1 => n15157, A2 => n14846, B1 => n14890, B2 => 
                           n14845, ZN => n14847);
   U2499 : OAI21_X1 port map( B1 => n15363, B2 => n14848, A => n14847, ZN => 
                           OUT2(23));
   U2500 : AOI22_X1 port map( A1 => n10065, A2 => n9165, B1 => n11174, B2 => 
                           n9069, ZN => n14852);
   U2501 : AOI22_X1 port map( A1 => n11186, A2 => n9325, B1 => n10070, B2 => 
                           n9389, ZN => n14851);
   U2502 : AOI22_X1 port map( A1 => n11190, A2 => n9133, B1 => n11187, B2 => 
                           n9421, ZN => n14850);
   U2503 : AOI22_X1 port map( A1 => n11189, A2 => n9101, B1 => n11165, B2 => 
                           n9293, ZN => n14849);
   U2504 : NAND4_X1 port map( A1 => n14852, A2 => n14851, A3 => n14850, A4 => 
                           n14849, ZN => n14858);
   U2505 : AOI22_X1 port map( A1 => n11188, A2 => n9357, B1 => n11166, B2 => 
                           n9229, ZN => n14856);
   U2506 : AOI22_X1 port map( A1 => n10060, A2 => n9261, B1 => n11173, B2 => 
                           n9197, ZN => n14855);
   U2507 : AOI22_X1 port map( A1 => n11168, A2 => n9453, B1 => n11162, B2 => 
                           n9485, ZN => n14854);
   U2508 : AOI22_X1 port map( A1 => n10067, A2 => n9037, B1 => n11167, B2 => 
                           n9517, ZN => n14853);
   U2509 : NAND4_X1 port map( A1 => n14856, A2 => n14855, A3 => n14854, A4 => 
                           n14853, ZN => n14857);
   U2510 : NOR2_X1 port map( A1 => n14858, A2 => n14857, ZN => n14870);
   U2511 : AOI22_X1 port map( A1 => n11185, A2 => n9933, B1 => n11163, B2 => 
                           n9805, ZN => n14862);
   U2512 : AOI22_X1 port map( A1 => n15325, A2 => n9965, B1 => n11184, B2 => 
                           n9837, ZN => n14861);
   U2513 : AOI22_X1 port map( A1 => n15352, A2 => n10029, B1 => n11178, B2 => 
                           n9901, ZN => n14860);
   U2514 : AOI22_X1 port map( A1 => n11177, A2 => n9869, B1 => n11176, B2 => 
                           n9997, ZN => n14859);
   U2515 : NAND4_X1 port map( A1 => n14862, A2 => n14861, A3 => n14860, A4 => 
                           n14859, ZN => n14868);
   U2516 : AOI22_X1 port map( A1 => n15352, A2 => n9773, B1 => n11159, B2 => 
                           n9677, ZN => n14866);
   U2517 : AOI22_X1 port map( A1 => n11226, A2 => n9709, B1 => n11160, B2 => 
                           n9581, ZN => n14865);
   U2518 : AOI22_X1 port map( A1 => n11176, A2 => n9741, B1 => n11163, B2 => 
                           n9549, ZN => n14864);
   U2519 : AOI22_X1 port map( A1 => n11177, A2 => n9613, B1 => n11161, B2 => 
                           n9645, ZN => n14863);
   U2520 : NAND4_X1 port map( A1 => n14866, A2 => n14865, A3 => n14864, A4 => 
                           n14863, ZN => n14867);
   U2521 : AOI22_X1 port map( A1 => n15157, A2 => n14868, B1 => n14890, B2 => 
                           n14867, ZN => n14869);
   U2522 : OAI21_X1 port map( B1 => n15363, B2 => n14870, A => n14869, ZN => 
                           OUT2(22));
   U2523 : AOI22_X1 port map( A1 => n11190, A2 => n9132, B1 => n11187, B2 => 
                           n9420, ZN => n14874);
   U2524 : AOI22_X1 port map( A1 => n11167, A2 => n9516, B1 => n11165, B2 => 
                           n9292, ZN => n14873);
   U2525 : AOI22_X1 port map( A1 => n10069, A2 => n9068, B1 => n11166, B2 => 
                           n9228, ZN => n14872);
   U2526 : AOI22_X1 port map( A1 => n11175, A2 => n9388, B1 => n11162, B2 => 
                           n9484, ZN => n14871);
   U2527 : NAND4_X1 port map( A1 => n14874, A2 => n14873, A3 => n14872, A4 => 
                           n14871, ZN => n14880);
   U2528 : AOI22_X1 port map( A1 => n11191, A2 => n9036, B1 => n11189, B2 => 
                           n9100, ZN => n14878);
   U2529 : AOI22_X1 port map( A1 => n11173, A2 => n9196, B1 => n11168, B2 => 
                           n9452, ZN => n14877);
   U2530 : AOI22_X1 port map( A1 => n10065, A2 => n9164, B1 => n10060, B2 => 
                           n9260, ZN => n14876);
   U2531 : AOI22_X1 port map( A1 => n11186, A2 => n9324, B1 => n11188, B2 => 
                           n9356, ZN => n14875);
   U2532 : NAND4_X1 port map( A1 => n14878, A2 => n14877, A3 => n14876, A4 => 
                           n14875, ZN => n14879);
   U2533 : NOR2_X1 port map( A1 => n14880, A2 => n14879, ZN => n14893);
   U2534 : AOI22_X1 port map( A1 => n11184, A2 => n9836, B1 => n11163, B2 => 
                           n9804, ZN => n14884);
   U2535 : AOI22_X1 port map( A1 => n11226, A2 => n9964, B1 => n11158, B2 => 
                           n10028, ZN => n14883);
   U2536 : AOI22_X1 port map( A1 => n11178, A2 => n9900, B1 => n11170, B2 => 
                           n9932, ZN => n14882);
   U2537 : AOI22_X1 port map( A1 => n11180, A2 => n9868, B1 => n11176, B2 => 
                           n9996, ZN => n14881);
   U2538 : NAND4_X1 port map( A1 => n14884, A2 => n14883, A3 => n14882, A4 => 
                           n14881, ZN => n14891);
   U2539 : AOI22_X1 port map( A1 => n11181, A2 => n9740, B1 => n11184, B2 => 
                           n9580, ZN => n14888);
   U2540 : AOI22_X1 port map( A1 => n15325, A2 => n9708, B1 => n11163, B2 => 
                           n9548, ZN => n14887);
   U2541 : AOI22_X1 port map( A1 => n15352, A2 => n9772, B1 => n11170, B2 => 
                           n9676, ZN => n14886);
   U2542 : AOI22_X1 port map( A1 => n11177, A2 => n9612, B1 => n11178, B2 => 
                           n9644, ZN => n14885);
   U2543 : NAND4_X1 port map( A1 => n14888, A2 => n14887, A3 => n14886, A4 => 
                           n14885, ZN => n14889);
   U2544 : AOI22_X1 port map( A1 => n15157, A2 => n14891, B1 => n14890, B2 => 
                           n14889, ZN => n14892);
   U2545 : OAI21_X1 port map( B1 => n15363, B2 => n14893, A => n14892, ZN => 
                           OUT2(21));
   U2546 : AOI22_X1 port map( A1 => n11186, A2 => n9323, B1 => n11172, B2 => 
                           n9163, ZN => n14897);
   U2547 : AOI22_X1 port map( A1 => n10064, A2 => n9227, B1 => n11175, B2 => 
                           n9387, ZN => n14896);
   U2548 : AOI22_X1 port map( A1 => n11190, A2 => n9131, B1 => n11162, B2 => 
                           n9483, ZN => n14895);
   U2549 : AOI22_X1 port map( A1 => n11187, A2 => n9419, B1 => n10067, B2 => 
                           n9035, ZN => n14894);
   U2550 : NAND4_X1 port map( A1 => n14897, A2 => n14896, A3 => n14895, A4 => 
                           n14894, ZN => n14903);
   U2551 : AOI22_X1 port map( A1 => n10060, A2 => n9259, B1 => n11165, B2 => 
                           n9291, ZN => n14901);
   U2552 : AOI22_X1 port map( A1 => n11189, A2 => n9099, B1 => n11167, B2 => 
                           n9515, ZN => n14900);
   U2553 : AOI22_X1 port map( A1 => n10069, A2 => n9067, B1 => n11173, B2 => 
                           n9195, ZN => n14899);
   U2554 : AOI22_X1 port map( A1 => n11188, A2 => n9355, B1 => n11168, B2 => 
                           n9451, ZN => n14898);
   U2555 : NAND4_X1 port map( A1 => n14901, A2 => n14900, A3 => n14899, A4 => 
                           n14898, ZN => n14902);
   U2556 : NOR2_X1 port map( A1 => n14903, A2 => n14902, ZN => n14915);
   U2557 : AOI22_X1 port map( A1 => n11178, A2 => n9899, B1 => n11163, B2 => 
                           n9803, ZN => n14907);
   U2558 : AOI22_X1 port map( A1 => n15325, A2 => n9963, B1 => n11180, B2 => 
                           n9867, ZN => n14906);
   U2559 : AOI22_X1 port map( A1 => n11227, A2 => n10027, B1 => n11185, B2 => 
                           n9931, ZN => n14905);
   U2560 : AOI22_X1 port map( A1 => n11176, A2 => n9995, B1 => n11160, B2 => 
                           n9835, ZN => n14904);
   U2561 : NAND4_X1 port map( A1 => n14907, A2 => n14906, A3 => n14905, A4 => 
                           n14904, ZN => n14913);
   U2562 : AOI22_X1 port map( A1 => n11180, A2 => n9611, B1 => n11185, B2 => 
                           n9675, ZN => n14911);
   U2563 : AOI22_X1 port map( A1 => n11169, A2 => n9739, B1 => n11163, B2 => 
                           n9547, ZN => n14910);
   U2564 : AOI22_X1 port map( A1 => n15352, A2 => n9771, B1 => n11171, B2 => 
                           n9579, ZN => n14909);
   U2565 : AOI22_X1 port map( A1 => n11161, A2 => n9643, B1 => n11156, B2 => 
                           n9707, ZN => n14908);
   U2566 : NAND4_X1 port map( A1 => n14911, A2 => n14910, A3 => n14909, A4 => 
                           n14908, ZN => n14912);
   U2567 : AOI22_X1 port map( A1 => n15157, A2 => n14913, B1 => n15358, B2 => 
                           n14912, ZN => n14914);
   U2568 : OAI21_X1 port map( B1 => n15363, B2 => n14915, A => n14914, ZN => 
                           OUT2(20));
   U2569 : AOI22_X1 port map( A1 => n11191, A2 => n9034, B1 => n11189, B2 => 
                           n9098, ZN => n14919);
   U2570 : AOI22_X1 port map( A1 => n11167, A2 => n9514, B1 => n11165, B2 => 
                           n9290, ZN => n14918);
   U2571 : AOI22_X1 port map( A1 => n11187, A2 => n9418, B1 => n11157, B2 => 
                           n9258, ZN => n14917);
   U2572 : AOI22_X1 port map( A1 => n11186, A2 => n9322, B1 => n10064, B2 => 
                           n9226, ZN => n14916);
   U2573 : NAND4_X1 port map( A1 => n14919, A2 => n14918, A3 => n14917, A4 => 
                           n14916, ZN => n14925);
   U2574 : AOI22_X1 port map( A1 => n11188, A2 => n9354, B1 => n11173, B2 => 
                           n9194, ZN => n14923);
   U2575 : AOI22_X1 port map( A1 => n11190, A2 => n9130, B1 => n11174, B2 => 
                           n9066, ZN => n14922);
   U2576 : AOI22_X1 port map( A1 => n11175, A2 => n9386, B1 => n11168, B2 => 
                           n9450, ZN => n14921);
   U2577 : AOI22_X1 port map( A1 => n10055, A2 => n9482, B1 => n11172, B2 => 
                           n9162, ZN => n14920);
   U2578 : NAND4_X1 port map( A1 => n14923, A2 => n14922, A3 => n14921, A4 => 
                           n14920, ZN => n14924);
   U2579 : NOR2_X1 port map( A1 => n14925, A2 => n14924, ZN => n14937);
   U2580 : AOI22_X1 port map( A1 => n11184, A2 => n9834, B1 => n11183, B2 => 
                           n9802, ZN => n14929);
   U2581 : AOI22_X1 port map( A1 => n11180, A2 => n9866, B1 => n11185, B2 => 
                           n9930, ZN => n14928);
   U2582 : AOI22_X1 port map( A1 => n11227, A2 => n10026, B1 => n11178, B2 => 
                           n9898, ZN => n14927);
   U2583 : AOI22_X1 port map( A1 => n11226, A2 => n9962, B1 => n11176, B2 => 
                           n9994, ZN => n14926);
   U2584 : NAND4_X1 port map( A1 => n14929, A2 => n14928, A3 => n14927, A4 => 
                           n14926, ZN => n14935);
   U2585 : AOI22_X1 port map( A1 => n11180, A2 => n9610, B1 => n11176, B2 => 
                           n9738, ZN => n14933);
   U2586 : AOI22_X1 port map( A1 => n11171, A2 => n9578, B1 => n11161, B2 => 
                           n9642, ZN => n14932);
   U2587 : AOI22_X1 port map( A1 => n11227, A2 => n9770, B1 => n11185, B2 => 
                           n9674, ZN => n14931);
   U2588 : AOI22_X1 port map( A1 => n11226, A2 => n9706, B1 => n11163, B2 => 
                           n9546, ZN => n14930);
   U2589 : NAND4_X1 port map( A1 => n14933, A2 => n14932, A3 => n14931, A4 => 
                           n14930, ZN => n14934);
   U2590 : AOI22_X1 port map( A1 => n15157, A2 => n14935, B1 => n15358, B2 => 
                           n14934, ZN => n14936);
   U2591 : OAI21_X1 port map( B1 => n15363, B2 => n14937, A => n14936, ZN => 
                           OUT2(19));
   U2592 : AOI22_X1 port map( A1 => n11175, A2 => n9385, B1 => n11157, B2 => 
                           n9257, ZN => n14941);
   U2593 : AOI22_X1 port map( A1 => n11186, A2 => n9321, B1 => n11190, B2 => 
                           n9129, ZN => n14940);
   U2594 : AOI22_X1 port map( A1 => n11187, A2 => n9417, B1 => n9097, B2 => 
                           n10059, ZN => n14939);
   U2595 : AOI22_X1 port map( A1 => n11167, A2 => n9513, B1 => n11168, B2 => 
                           n9449, ZN => n14938);
   U2596 : NAND4_X1 port map( A1 => n14941, A2 => n14940, A3 => n14939, A4 => 
                           n14938, ZN => n14947);
   U2597 : AOI22_X1 port map( A1 => n10055, A2 => n9481, B1 => n10065, B2 => 
                           n9161, ZN => n14945);
   U2598 : AOI22_X1 port map( A1 => n11191, A2 => n9033, B1 => n11174, B2 => 
                           n9065, ZN => n14944);
   U2599 : AOI22_X1 port map( A1 => n10064, A2 => n9225, B1 => n11165, B2 => 
                           n9289, ZN => n14943);
   U2600 : AOI22_X1 port map( A1 => n10068, A2 => n9193, B1 => n11188, B2 => 
                           n9353, ZN => n14942);
   U2601 : NAND4_X1 port map( A1 => n14945, A2 => n14944, A3 => n14943, A4 => 
                           n14942, ZN => n14946);
   U2602 : NOR2_X1 port map( A1 => n14947, A2 => n14946, ZN => n14959);
   U2603 : CLKBUF_X1 port map( A => n15112, Z => n15360);
   U2604 : AOI22_X1 port map( A1 => n11178, A2 => n9897, B1 => n11171, B2 => 
                           n9833, ZN => n14951);
   U2605 : AOI22_X1 port map( A1 => n11227, A2 => n10025, B1 => n11226, B2 => 
                           n9961, ZN => n14950);
   U2606 : AOI22_X1 port map( A1 => n11177, A2 => n9865, B1 => n11179, B2 => 
                           n9801, ZN => n14949);
   U2607 : AOI22_X1 port map( A1 => n11181, A2 => n9993, B1 => n11185, B2 => 
                           n9929, ZN => n14948);
   U2608 : NAND4_X1 port map( A1 => n14951, A2 => n14950, A3 => n14949, A4 => 
                           n14948, ZN => n14957);
   U2609 : AOI22_X1 port map( A1 => n15352, A2 => n9769, B1 => n11180, B2 => 
                           n9609, ZN => n14955);
   U2610 : AOI22_X1 port map( A1 => n11161, A2 => n9641, B1 => n11156, B2 => 
                           n9705, ZN => n14954);
   U2611 : AOI22_X1 port map( A1 => n11183, A2 => n9545, B1 => n11169, B2 => 
                           n9737, ZN => n14953);
   U2612 : AOI22_X1 port map( A1 => n11185, A2 => n9673, B1 => n11171, B2 => 
                           n9577, ZN => n14952);
   U2613 : NAND4_X1 port map( A1 => n14955, A2 => n14954, A3 => n14953, A4 => 
                           n14952, ZN => n14956);
   U2614 : AOI22_X1 port map( A1 => n15360, A2 => n14957, B1 => n15358, B2 => 
                           n14956, ZN => n14958);
   U2615 : OAI21_X1 port map( B1 => n15363, B2 => n14959, A => n14958, ZN => 
                           OUT2(18));
   U2616 : AOI22_X1 port map( A1 => n11189, A2 => n9096, B1 => n11157, B2 => 
                           n9256, ZN => n14963);
   U2617 : AOI22_X1 port map( A1 => n11191, A2 => n9032, B1 => n10064, B2 => 
                           n9224, ZN => n14962);
   U2618 : AOI22_X1 port map( A1 => n11190, A2 => n9128, B1 => n11173, B2 => 
                           n9192, ZN => n14961);
   U2619 : AOI22_X1 port map( A1 => n11175, A2 => n9384, B1 => n11167, B2 => 
                           n9512, ZN => n14960);
   U2620 : NAND4_X1 port map( A1 => n14963, A2 => n14962, A3 => n14961, A4 => 
                           n14960, ZN => n14969);
   U2621 : AOI22_X1 port map( A1 => n11188, A2 => n9352, B1 => n11165, B2 => 
                           n9288, ZN => n14967);
   U2622 : AOI22_X1 port map( A1 => n11186, A2 => n9320, B1 => n11162, B2 => 
                           n9480, ZN => n14966);
   U2623 : AOI22_X1 port map( A1 => n11172, A2 => n9160, B1 => n11168, B2 => 
                           n9448, ZN => n14965);
   U2624 : AOI22_X1 port map( A1 => n11174, A2 => n9064, B1 => n10057, B2 => 
                           n9416, ZN => n14964);
   U2625 : NAND4_X1 port map( A1 => n14967, A2 => n14966, A3 => n14965, A4 => 
                           n14964, ZN => n14968);
   U2626 : NOR2_X1 port map( A1 => n14969, A2 => n14968, ZN => n14981);
   U2627 : AOI22_X1 port map( A1 => n11178, A2 => n9896, B1 => n11156, B2 => 
                           n9960, ZN => n14973);
   U2628 : AOI22_X1 port map( A1 => n11184, A2 => n9832, B1 => n11185, B2 => 
                           n9928, ZN => n14972);
   U2629 : AOI22_X1 port map( A1 => n11180, A2 => n9864, B1 => n11169, B2 => 
                           n9992, ZN => n14971);
   U2630 : AOI22_X1 port map( A1 => n11227, A2 => n10024, B1 => n11179, B2 => 
                           n9800, ZN => n14970);
   U2631 : NAND4_X1 port map( A1 => n14973, A2 => n14972, A3 => n14971, A4 => 
                           n14970, ZN => n14979);
   U2632 : AOI22_X1 port map( A1 => n11181, A2 => n9736, B1 => n11179, B2 => 
                           n9544, ZN => n14977);
   U2633 : AOI22_X1 port map( A1 => n11180, A2 => n9608, B1 => n11185, B2 => 
                           n9672, ZN => n14976);
   U2634 : AOI22_X1 port map( A1 => n11227, A2 => n9768, B1 => n11178, B2 => 
                           n9640, ZN => n14975);
   U2635 : AOI22_X1 port map( A1 => n11226, A2 => n9704, B1 => n11171, B2 => 
                           n9576, ZN => n14974);
   U2636 : NAND4_X1 port map( A1 => n14977, A2 => n14976, A3 => n14975, A4 => 
                           n14974, ZN => n14978);
   U2637 : AOI22_X1 port map( A1 => n15360, A2 => n14979, B1 => n15358, B2 => 
                           n14978, ZN => n14980);
   U2638 : OAI21_X1 port map( B1 => n15363, B2 => n14981, A => n14980, ZN => 
                           OUT2(17));
   U2639 : AOI22_X1 port map( A1 => n10058, A2 => n9351, B1 => n11162, B2 => 
                           n9479, ZN => n14985);
   U2640 : AOI22_X1 port map( A1 => n10067, A2 => n9031, B1 => n10061, B2 => 
                           n9127, ZN => n14984);
   U2641 : AOI22_X1 port map( A1 => n10069, A2 => n9063, B1 => n11175, B2 => 
                           n9383, ZN => n14983);
   U2642 : AOI22_X1 port map( A1 => n11186, A2 => n9319, B1 => n11173, B2 => 
                           n9191, ZN => n14982);
   U2643 : NAND4_X1 port map( A1 => n14985, A2 => n14984, A3 => n14983, A4 => 
                           n14982, ZN => n14991);
   U2644 : AOI22_X1 port map( A1 => n11166, A2 => n9223, B1 => n11157, B2 => 
                           n9255, ZN => n14989);
   U2645 : AOI22_X1 port map( A1 => n10063, A2 => n9287, B1 => n11167, B2 => 
                           n9511, ZN => n14988);
   U2646 : AOI22_X1 port map( A1 => n11172, A2 => n9159, B1 => n11168, B2 => 
                           n9447, ZN => n14987);
   U2647 : AOI22_X1 port map( A1 => n11189, A2 => n9095, B1 => n11187, B2 => 
                           n9415, ZN => n14986);
   U2648 : NAND4_X1 port map( A1 => n14989, A2 => n14988, A3 => n14987, A4 => 
                           n14986, ZN => n14990);
   U2649 : NOR2_X1 port map( A1 => n14991, A2 => n14990, ZN => n15003);
   U2650 : AOI22_X1 port map( A1 => n11180, A2 => n9863, B1 => n11160, B2 => 
                           n9831, ZN => n14995);
   U2651 : AOI22_X1 port map( A1 => n15325, A2 => n9959, B1 => n11185, B2 => 
                           n9927, ZN => n14994);
   U2652 : AOI22_X1 port map( A1 => n11227, A2 => n10023, B1 => n11163, B2 => 
                           n9799, ZN => n14993);
   U2653 : AOI22_X1 port map( A1 => n11182, A2 => n9895, B1 => n11169, B2 => 
                           n9991, ZN => n14992);
   U2654 : NAND4_X1 port map( A1 => n14995, A2 => n14994, A3 => n14993, A4 => 
                           n14992, ZN => n15001);
   U2655 : AOI22_X1 port map( A1 => n15352, A2 => n9767, B1 => n11160, B2 => 
                           n9575, ZN => n14999);
   U2656 : AOI22_X1 port map( A1 => n11176, A2 => n9735, B1 => n11159, B2 => 
                           n9671, ZN => n14998);
   U2657 : AOI22_X1 port map( A1 => n11226, A2 => n9703, B1 => n11163, B2 => 
                           n9543, ZN => n14997);
   U2658 : AOI22_X1 port map( A1 => n11180, A2 => n9607, B1 => n11161, B2 => 
                           n9639, ZN => n14996);
   U2659 : NAND4_X1 port map( A1 => n14999, A2 => n14998, A3 => n14997, A4 => 
                           n14996, ZN => n15000);
   U2660 : AOI22_X1 port map( A1 => n15157, A2 => n15001, B1 => n15358, B2 => 
                           n15000, ZN => n15002);
   U2661 : OAI21_X1 port map( B1 => n15363, B2 => n15003, A => n15002, ZN => 
                           OUT2(16));
   U2662 : AOI22_X1 port map( A1 => n11167, A2 => n9510, B1 => n10059, B2 => 
                           n9094, ZN => n15007);
   U2663 : AOI22_X1 port map( A1 => n10065, A2 => n9158, B1 => n11190, B2 => 
                           n9126, ZN => n15006);
   U2664 : AOI22_X1 port map( A1 => n11186, A2 => n9318, B1 => n11175, B2 => 
                           n9382, ZN => n15005);
   U2665 : AOI22_X1 port map( A1 => n11191, A2 => n9030, B1 => n11174, B2 => 
                           n9062, ZN => n15004);
   U2666 : NAND4_X1 port map( A1 => n15007, A2 => n15006, A3 => n15005, A4 => 
                           n15004, ZN => n15013);
   U2667 : AOI22_X1 port map( A1 => n10068, A2 => n9190, B1 => n11168, B2 => 
                           n9446, ZN => n15011);
   U2668 : AOI22_X1 port map( A1 => n11166, A2 => n9222, B1 => n11162, B2 => 
                           n9478, ZN => n15010);
   U2669 : AOI22_X1 port map( A1 => n10063, A2 => n9286, B1 => n10057, B2 => 
                           n9414, ZN => n15009);
   U2670 : AOI22_X1 port map( A1 => n11188, A2 => n9350, B1 => n11157, B2 => 
                           n9254, ZN => n15008);
   U2671 : NAND4_X1 port map( A1 => n15011, A2 => n15010, A3 => n15009, A4 => 
                           n15008, ZN => n15012);
   U2672 : NOR2_X1 port map( A1 => n15013, A2 => n15012, ZN => n15025);
   U2673 : AOI22_X1 port map( A1 => n11227, A2 => n10022, B1 => n11182, B2 => 
                           n9894, ZN => n15017);
   U2674 : AOI22_X1 port map( A1 => n11183, A2 => n9798, B1 => n11185, B2 => 
                           n9926, ZN => n15016);
   U2675 : AOI22_X1 port map( A1 => n11171, A2 => n9830, B1 => n11156, B2 => 
                           n9958, ZN => n15015);
   U2676 : AOI22_X1 port map( A1 => n11177, A2 => n9862, B1 => n11176, B2 => 
                           n9990, ZN => n15014);
   U2677 : NAND4_X1 port map( A1 => n15017, A2 => n15016, A3 => n15015, A4 => 
                           n15014, ZN => n15023);
   U2678 : AOI22_X1 port map( A1 => n11176, A2 => n9734, B1 => n11171, B2 => 
                           n9574, ZN => n15021);
   U2679 : AOI22_X1 port map( A1 => n11226, A2 => n9702, B1 => n11180, B2 => 
                           n9606, ZN => n15020);
   U2680 : AOI22_X1 port map( A1 => n11185, A2 => n9670, B1 => n11161, B2 => 
                           n9638, ZN => n15019);
   U2681 : AOI22_X1 port map( A1 => n11227, A2 => n9766, B1 => n11163, B2 => 
                           n9542, ZN => n15018);
   U2682 : NAND4_X1 port map( A1 => n15021, A2 => n15020, A3 => n15019, A4 => 
                           n15018, ZN => n15022);
   U2683 : AOI22_X1 port map( A1 => n15157, A2 => n15023, B1 => n15358, B2 => 
                           n15022, ZN => n15024);
   U2684 : OAI21_X1 port map( B1 => n15363, B2 => n15025, A => n15024, ZN => 
                           OUT2(15));
   U2685 : AOI22_X1 port map( A1 => n10070, A2 => n9381, B1 => n11173, B2 => 
                           n9189, ZN => n15029);
   U2686 : AOI22_X1 port map( A1 => n11188, A2 => n9349, B1 => n11172, B2 => 
                           n9157, ZN => n15028);
   U2687 : AOI22_X1 port map( A1 => n10069, A2 => n9061, B1 => n11162, B2 => 
                           n9477, ZN => n15027);
   U2688 : AOI22_X1 port map( A1 => n11166, A2 => n9221, B1 => n11165, B2 => 
                           n9285, ZN => n15026);
   U2689 : NAND4_X1 port map( A1 => n15029, A2 => n15028, A3 => n15027, A4 => 
                           n15026, ZN => n15035);
   U2690 : AOI22_X1 port map( A1 => n11189, A2 => n9093, B1 => n10057, B2 => 
                           n9413, ZN => n15033);
   U2691 : AOI22_X1 port map( A1 => n11186, A2 => n9317, B1 => n11157, B2 => 
                           n9253, ZN => n15032);
   U2692 : AOI22_X1 port map( A1 => n10066, A2 => n9445, B1 => n11167, B2 => 
                           n9509, ZN => n15031);
   U2693 : AOI22_X1 port map( A1 => n10067, A2 => n9029, B1 => n10061, B2 => 
                           n9125, ZN => n15030);
   U2694 : NAND4_X1 port map( A1 => n15033, A2 => n15032, A3 => n15031, A4 => 
                           n15030, ZN => n15034);
   U2695 : NOR2_X1 port map( A1 => n15035, A2 => n15034, ZN => n15047);
   U2696 : AOI22_X1 port map( A1 => n11227, A2 => n10021, B1 => n11160, B2 => 
                           n9829, ZN => n15039);
   U2697 : AOI22_X1 port map( A1 => n11170, A2 => n9925, B1 => n11161, B2 => 
                           n9893, ZN => n15038);
   U2698 : AOI22_X1 port map( A1 => n11163, A2 => n9797, B1 => n11156, B2 => 
                           n9957, ZN => n15037);
   U2699 : AOI22_X1 port map( A1 => n11177, A2 => n9861, B1 => n11169, B2 => 
                           n9989, ZN => n15036);
   U2700 : NAND4_X1 port map( A1 => n15039, A2 => n15038, A3 => n15037, A4 => 
                           n15036, ZN => n15045);
   U2701 : AOI22_X1 port map( A1 => n11170, A2 => n9669, B1 => n11161, B2 => 
                           n9637, ZN => n15043);
   U2702 : AOI22_X1 port map( A1 => n11181, A2 => n9733, B1 => n11163, B2 => 
                           n9541, ZN => n15042);
   U2703 : AOI22_X1 port map( A1 => n15352, A2 => n9765, B1 => n11156, B2 => 
                           n9701, ZN => n15041);
   U2704 : AOI22_X1 port map( A1 => n11180, A2 => n9605, B1 => n11171, B2 => 
                           n9573, ZN => n15040);
   U2705 : NAND4_X1 port map( A1 => n15043, A2 => n15042, A3 => n15041, A4 => 
                           n15040, ZN => n15044);
   U2706 : AOI22_X1 port map( A1 => n15157, A2 => n15045, B1 => n15358, B2 => 
                           n15044, ZN => n15046);
   U2707 : OAI21_X1 port map( B1 => n15363, B2 => n15047, A => n15046, ZN => 
                           OUT2(14));
   U2708 : AOI22_X1 port map( A1 => n11157, A2 => n9252, B1 => n10059, B2 => 
                           n9092, ZN => n15051);
   U2709 : AOI22_X1 port map( A1 => n10068, A2 => n9188, B1 => n11174, B2 => 
                           n9060, ZN => n15050);
   U2710 : AOI22_X1 port map( A1 => n11190, A2 => n9124, B1 => n11166, B2 => 
                           n9220, ZN => n15049);
   U2711 : AOI22_X1 port map( A1 => n10056, A2 => n9316, B1 => n11175, B2 => 
                           n9380, ZN => n15048);
   U2712 : NAND4_X1 port map( A1 => n15051, A2 => n15050, A3 => n15049, A4 => 
                           n15048, ZN => n15057);
   U2713 : AOI22_X1 port map( A1 => n10058, A2 => n9348, B1 => n11168, B2 => 
                           n9444, ZN => n15055);
   U2714 : AOI22_X1 port map( A1 => n11187, A2 => n9412, B1 => n11167, B2 => 
                           n9508, ZN => n15054);
   U2715 : AOI22_X1 port map( A1 => n11191, A2 => n9028, B1 => n11165, B2 => 
                           n9284, ZN => n15053);
   U2716 : AOI22_X1 port map( A1 => n10065, A2 => n9156, B1 => n11162, B2 => 
                           n9476, ZN => n15052);
   U2717 : NAND4_X1 port map( A1 => n15055, A2 => n15054, A3 => n15053, A4 => 
                           n15052, ZN => n15056);
   U2718 : NOR2_X1 port map( A1 => n15057, A2 => n15056, ZN => n15069);
   U2719 : AOI22_X1 port map( A1 => n11227, A2 => n10020, B1 => n11161, B2 => 
                           n9892, ZN => n15061);
   U2720 : AOI22_X1 port map( A1 => n11183, A2 => n9796, B1 => n11185, B2 => 
                           n9924, ZN => n15060);
   U2721 : AOI22_X1 port map( A1 => n11169, A2 => n9988, B1 => n11164, B2 => 
                           n9860, ZN => n15059);
   U2722 : AOI22_X1 port map( A1 => n11160, A2 => n9828, B1 => n11156, B2 => 
                           n9956, ZN => n15058);
   U2723 : NAND4_X1 port map( A1 => n15061, A2 => n15060, A3 => n15059, A4 => 
                           n15058, ZN => n15067);
   U2724 : AOI22_X1 port map( A1 => n11183, A2 => n9540, B1 => n11169, B2 => 
                           n9732, ZN => n15065);
   U2725 : AOI22_X1 port map( A1 => n11164, A2 => n9604, B1 => n11160, B2 => 
                           n9572, ZN => n15064);
   U2726 : AOI22_X1 port map( A1 => n11182, A2 => n9636, B1 => n11185, B2 => 
                           n9668, ZN => n15063);
   U2727 : AOI22_X1 port map( A1 => n11227, A2 => n9764, B1 => n11156, B2 => 
                           n9700, ZN => n15062);
   U2728 : NAND4_X1 port map( A1 => n15065, A2 => n15064, A3 => n15063, A4 => 
                           n15062, ZN => n15066);
   U2729 : AOI22_X1 port map( A1 => n15157, A2 => n15067, B1 => n15358, B2 => 
                           n15066, ZN => n15068);
   U2730 : OAI21_X1 port map( B1 => n15363, B2 => n15069, A => n15068, ZN => 
                           OUT2(13));
   U2731 : AOI22_X1 port map( A1 => n11174, A2 => n9059, B1 => n10059, B2 => 
                           n9091, ZN => n15073);
   U2732 : AOI22_X1 port map( A1 => n11162, A2 => n9475, B1 => n11157, B2 => 
                           n9251, ZN => n15072);
   U2733 : AOI22_X1 port map( A1 => n10062, A2 => n9507, B1 => n10063, B2 => 
                           n9283, ZN => n15071);
   U2734 : AOI22_X1 port map( A1 => n10068, A2 => n9187, B1 => n10061, B2 => 
                           n9123, ZN => n15070);
   U2735 : NAND4_X1 port map( A1 => n15073, A2 => n15072, A3 => n15071, A4 => 
                           n15070, ZN => n15079);
   U2736 : AOI22_X1 port map( A1 => n11175, A2 => n9379, B1 => n11168, B2 => 
                           n9443, ZN => n15077);
   U2737 : AOI22_X1 port map( A1 => n11188, A2 => n9347, B1 => n10067, B2 => 
                           n9027, ZN => n15076);
   U2738 : AOI22_X1 port map( A1 => n10065, A2 => n9155, B1 => n11186, B2 => 
                           n9315, ZN => n15075);
   U2739 : AOI22_X1 port map( A1 => n10057, A2 => n9411, B1 => n11166, B2 => 
                           n9219, ZN => n15074);
   U2740 : NAND4_X1 port map( A1 => n15077, A2 => n15076, A3 => n15075, A4 => 
                           n15074, ZN => n15078);
   U2741 : NOR2_X1 port map( A1 => n15079, A2 => n15078, ZN => n15091);
   U2742 : AOI22_X1 port map( A1 => n11182, A2 => n9891, B1 => n11171, B2 => 
                           n9827, ZN => n15083);
   U2743 : AOI22_X1 port map( A1 => n11227, A2 => n10019, B1 => n11183, B2 => 
                           n9795, ZN => n15082);
   U2744 : AOI22_X1 port map( A1 => n11159, A2 => n9923, B1 => n11156, B2 => 
                           n9955, ZN => n15081);
   U2745 : AOI22_X1 port map( A1 => n11181, A2 => n9987, B1 => n11180, B2 => 
                           n9859, ZN => n15080);
   U2746 : NAND4_X1 port map( A1 => n15083, A2 => n15082, A3 => n15081, A4 => 
                           n15080, ZN => n15089);
   U2747 : AOI22_X1 port map( A1 => n11158, A2 => n9763, B1 => n11156, B2 => 
                           n9699, ZN => n15087);
   U2748 : AOI22_X1 port map( A1 => n11183, A2 => n9539, B1 => n11171, B2 => 
                           n9571, ZN => n15086);
   U2749 : AOI22_X1 port map( A1 => n11180, A2 => n9603, B1 => n11182, B2 => 
                           n9635, ZN => n15085);
   U2750 : AOI22_X1 port map( A1 => n11181, A2 => n9731, B1 => n11159, B2 => 
                           n9667, ZN => n15084);
   U2751 : NAND4_X1 port map( A1 => n15087, A2 => n15086, A3 => n15085, A4 => 
                           n15084, ZN => n15088);
   U2752 : AOI22_X1 port map( A1 => n15157, A2 => n15089, B1 => n15358, B2 => 
                           n15088, ZN => n15090);
   U2753 : OAI21_X1 port map( B1 => n15363, B2 => n15091, A => n15090, ZN => 
                           OUT2(12));
   U2754 : AOI22_X1 port map( A1 => n10068, A2 => n9186, B1 => n10063, B2 => 
                           n9282, ZN => n15095);
   U2755 : AOI22_X1 port map( A1 => n10069, A2 => n9058, B1 => n11187, B2 => 
                           n9410, ZN => n15094);
   U2756 : AOI22_X1 port map( A1 => n11175, A2 => n9378, B1 => n11166, B2 => 
                           n9218, ZN => n15093);
   U2757 : AOI22_X1 port map( A1 => n10062, A2 => n9506, B1 => n10061, B2 => 
                           n9122, ZN => n15092);
   U2758 : NAND4_X1 port map( A1 => n15095, A2 => n15094, A3 => n15093, A4 => 
                           n15092, ZN => n15101);
   U2759 : AOI22_X1 port map( A1 => n11172, A2 => n9154, B1 => n10056, B2 => 
                           n9314, ZN => n15099);
   U2760 : AOI22_X1 port map( A1 => n10058, A2 => n9346, B1 => n11157, B2 => 
                           n9250, ZN => n15098);
   U2761 : AOI22_X1 port map( A1 => n10067, A2 => n9026, B1 => n10059, B2 => 
                           n9090, ZN => n15097);
   U2762 : AOI22_X1 port map( A1 => n11168, A2 => n9442, B1 => n11162, B2 => 
                           n9474, ZN => n15096);
   U2763 : NAND4_X1 port map( A1 => n15099, A2 => n15098, A3 => n15097, A4 => 
                           n15096, ZN => n15100);
   U2764 : NOR2_X1 port map( A1 => n15101, A2 => n15100, ZN => n15114);
   U2765 : AOI22_X1 port map( A1 => n11180, A2 => n9858, B1 => n11183, B2 => 
                           n9794, ZN => n15105);
   U2766 : AOI22_X1 port map( A1 => n15352, A2 => n10018, B1 => n11156, B2 => 
                           n9954, ZN => n15104);
   U2767 : AOI22_X1 port map( A1 => n11171, A2 => n9826, B1 => n11159, B2 => 
                           n9922, ZN => n15103);
   U2768 : AOI22_X1 port map( A1 => n11181, A2 => n9986, B1 => n11161, B2 => 
                           n9890, ZN => n15102);
   U2769 : NAND4_X1 port map( A1 => n15105, A2 => n15104, A3 => n15103, A4 => 
                           n15102, ZN => n15111);
   U2770 : AOI22_X1 port map( A1 => n11181, A2 => n9730, B1 => n11180, B2 => 
                           n9602, ZN => n15109);
   U2771 : AOI22_X1 port map( A1 => n11227, A2 => n9762, B1 => n11182, B2 => 
                           n9634, ZN => n15108);
   U2772 : AOI22_X1 port map( A1 => n11183, A2 => n9538, B1 => n11185, B2 => 
                           n9666, ZN => n15107);
   U2773 : AOI22_X1 port map( A1 => n11160, A2 => n9570, B1 => n11156, B2 => 
                           n9698, ZN => n15106);
   U2774 : NAND4_X1 port map( A1 => n15109, A2 => n15108, A3 => n15107, A4 => 
                           n15106, ZN => n15110);
   U2775 : AOI22_X1 port map( A1 => n15112, A2 => n15111, B1 => n15358, B2 => 
                           n15110, ZN => n15113);
   U2776 : OAI21_X1 port map( B1 => n15182, B2 => n15114, A => n15113, ZN => 
                           OUT2(11));
   U2777 : AOI22_X1 port map( A1 => n10066, A2 => n9441, B1 => n10056, B2 => 
                           n9313, ZN => n15118);
   U2778 : AOI22_X1 port map( A1 => n11174, A2 => n9057, B1 => n11157, B2 => 
                           n9249, ZN => n15117);
   U2779 : AOI22_X1 port map( A1 => n11189, A2 => n9089, B1 => n10068, B2 => 
                           n9185, ZN => n15116);
   U2780 : AOI22_X1 port map( A1 => n10063, A2 => n9281, B1 => n10061, B2 => 
                           n9121, ZN => n15115);
   U2781 : NAND4_X1 port map( A1 => n15118, A2 => n15117, A3 => n15116, A4 => 
                           n15115, ZN => n15124);
   U2782 : AOI22_X1 port map( A1 => n10057, A2 => n9409, B1 => n11166, B2 => 
                           n9217, ZN => n15122);
   U2783 : AOI22_X1 port map( A1 => n11172, A2 => n9153, B1 => n11167, B2 => 
                           n9505, ZN => n15121);
   U2784 : AOI22_X1 port map( A1 => n11191, A2 => n9025, B1 => n11175, B2 => 
                           n9377, ZN => n15120);
   U2785 : AOI22_X1 port map( A1 => n11188, A2 => n9345, B1 => n11162, B2 => 
                           n9473, ZN => n15119);
   U2786 : NAND4_X1 port map( A1 => n15122, A2 => n15121, A3 => n15120, A4 => 
                           n15119, ZN => n15123);
   U2787 : NOR2_X1 port map( A1 => n15124, A2 => n15123, ZN => n15136);
   U2788 : AOI22_X1 port map( A1 => n11183, A2 => n9793, B1 => n11164, B2 => 
                           n9857, ZN => n15128);
   U2789 : AOI22_X1 port map( A1 => n15352, A2 => n10017, B1 => n11184, B2 => 
                           n9825, ZN => n15127);
   U2790 : AOI22_X1 port map( A1 => n11181, A2 => n9985, B1 => n11156, B2 => 
                           n9953, ZN => n15126);
   U2791 : AOI22_X1 port map( A1 => n11182, A2 => n9889, B1 => n11159, B2 => 
                           n9921, ZN => n15125);
   U2792 : NAND4_X1 port map( A1 => n15128, A2 => n15127, A3 => n15126, A4 => 
                           n15125, ZN => n15134);
   U2793 : AOI22_X1 port map( A1 => n11164, A2 => n9601, B1 => n11156, B2 => 
                           n9697, ZN => n15132);
   U2794 : AOI22_X1 port map( A1 => n11161, A2 => n9633, B1 => n11159, B2 => 
                           n9665, ZN => n15131);
   U2795 : AOI22_X1 port map( A1 => n11227, A2 => n9761, B1 => n11169, B2 => 
                           n9729, ZN => n15130);
   U2796 : AOI22_X1 port map( A1 => n11184, A2 => n9569, B1 => n11183, B2 => 
                           n9537, ZN => n15129);
   U2797 : NAND4_X1 port map( A1 => n15132, A2 => n15131, A3 => n15130, A4 => 
                           n15129, ZN => n15133);
   U2798 : AOI22_X1 port map( A1 => n15157, A2 => n15134, B1 => n15358, B2 => 
                           n15133, ZN => n15135);
   U2799 : OAI21_X1 port map( B1 => n15182, B2 => n15136, A => n15135, ZN => 
                           OUT2(10));
   U2800 : AOI22_X1 port map( A1 => n10067, A2 => n9024, B1 => n11165, B2 => 
                           n9280, ZN => n15140);
   U2801 : AOI22_X1 port map( A1 => n10066, A2 => n9440, B1 => n11157, B2 => 
                           n9248, ZN => n15139);
   U2802 : AOI22_X1 port map( A1 => n10069, A2 => n9056, B1 => n11162, B2 => 
                           n9472, ZN => n15138);
   U2803 : AOI22_X1 port map( A1 => n10068, A2 => n9184, B1 => n10058, B2 => 
                           n9344, ZN => n15137);
   U2804 : NAND4_X1 port map( A1 => n15140, A2 => n15139, A3 => n15138, A4 => 
                           n15137, ZN => n15146);
   U2805 : AOI22_X1 port map( A1 => n10062, A2 => n9504, B1 => n11172, B2 => 
                           n9152, ZN => n15144);
   U2806 : AOI22_X1 port map( A1 => n11190, A2 => n9120, B1 => n11187, B2 => 
                           n9408, ZN => n15143);
   U2807 : AOI22_X1 port map( A1 => n10070, A2 => n9376, B1 => n10056, B2 => 
                           n9312, ZN => n15142);
   U2808 : AOI22_X1 port map( A1 => n11166, A2 => n9216, B1 => n10059, B2 => 
                           n9088, ZN => n15141);
   U2809 : NAND4_X1 port map( A1 => n15144, A2 => n15143, A3 => n15142, A4 => 
                           n15141, ZN => n15145);
   U2810 : NOR2_X1 port map( A1 => n15146, A2 => n15145, ZN => n15159);
   U2811 : AOI22_X1 port map( A1 => n11169, A2 => n9984, B1 => n11164, B2 => 
                           n9856, ZN => n15150);
   U2812 : AOI22_X1 port map( A1 => n11183, A2 => n9792, B1 => n11159, B2 => 
                           n9920, ZN => n15149);
   U2813 : AOI22_X1 port map( A1 => n11171, A2 => n9824, B1 => n11156, B2 => 
                           n9952, ZN => n15148);
   U2814 : AOI22_X1 port map( A1 => n15352, A2 => n10016, B1 => n11161, B2 => 
                           n9888, ZN => n15147);
   U2815 : NAND4_X1 port map( A1 => n15150, A2 => n15149, A3 => n15148, A4 => 
                           n15147, ZN => n15156);
   U2816 : AOI22_X1 port map( A1 => n11183, A2 => n9536, B1 => n11156, B2 => 
                           n9696, ZN => n15154);
   U2817 : AOI22_X1 port map( A1 => n11180, A2 => n9600, B1 => n11159, B2 => 
                           n9664, ZN => n15153);
   U2818 : AOI22_X1 port map( A1 => n11184, A2 => n9568, B1 => n11158, B2 => 
                           n9760, ZN => n15152);
   U2819 : AOI22_X1 port map( A1 => n11181, A2 => n9728, B1 => n11161, B2 => 
                           n9632, ZN => n15151);
   U2820 : NAND4_X1 port map( A1 => n15154, A2 => n15153, A3 => n15152, A4 => 
                           n15151, ZN => n15155);
   U2821 : AOI22_X1 port map( A1 => n15157, A2 => n15156, B1 => n15358, B2 => 
                           n15155, ZN => n15158);
   U2822 : OAI21_X1 port map( B1 => n15182, B2 => n15159, A => n15158, ZN => 
                           OUT2(9));
   U2823 : AOI22_X1 port map( A1 => n10070, A2 => n9375, B1 => n11167, B2 => 
                           n9503, ZN => n15163);
   U2824 : AOI22_X1 port map( A1 => n10064, A2 => n9215, B1 => n11157, B2 => 
                           n9247, ZN => n15162);
   U2825 : AOI22_X1 port map( A1 => n11186, A2 => n9311, B1 => n11172, B2 => 
                           n9151, ZN => n15161);
   U2826 : AOI22_X1 port map( A1 => n11173, A2 => n9183, B1 => n10067, B2 => 
                           n9023, ZN => n15160);
   U2827 : NAND4_X1 port map( A1 => n15163, A2 => n15162, A3 => n15161, A4 => 
                           n15160, ZN => n15169);
   U2828 : AOI22_X1 port map( A1 => n10055, A2 => n9471, B1 => n11187, B2 => 
                           n9407, ZN => n15167);
   U2829 : AOI22_X1 port map( A1 => n11174, A2 => n9055, B1 => n11168, B2 => 
                           n9439, ZN => n15166);
   U2830 : AOI22_X1 port map( A1 => n10063, A2 => n9279, B1 => n11190, B2 => 
                           n9119, ZN => n15165);
   U2831 : AOI22_X1 port map( A1 => n11188, A2 => n9343, B1 => n10059, B2 => 
                           n9087, ZN => n15164);
   U2832 : NAND4_X1 port map( A1 => n15167, A2 => n15166, A3 => n15165, A4 => 
                           n15164, ZN => n15168);
   U2833 : NOR2_X1 port map( A1 => n15169, A2 => n15168, ZN => n15181);
   U2834 : AOI22_X1 port map( A1 => n11183, A2 => n9791, B1 => n11164, B2 => 
                           n9855, ZN => n15173);
   U2835 : AOI22_X1 port map( A1 => n11227, A2 => n10015, B1 => n11159, B2 => 
                           n9919, ZN => n15172);
   U2836 : AOI22_X1 port map( A1 => n11160, A2 => n9823, B1 => n11156, B2 => 
                           n9951, ZN => n15171);
   U2837 : AOI22_X1 port map( A1 => n11181, A2 => n9983, B1 => n11182, B2 => 
                           n9887, ZN => n15170);
   U2838 : NAND4_X1 port map( A1 => n15173, A2 => n15172, A3 => n15171, A4 => 
                           n15170, ZN => n15179);
   U2839 : AOI22_X1 port map( A1 => n15352, A2 => n9759, B1 => n11185, B2 => 
                           n9663, ZN => n15177);
   U2840 : AOI22_X1 port map( A1 => n15325, A2 => n9695, B1 => n11180, B2 => 
                           n9599, ZN => n15176);
   U2841 : AOI22_X1 port map( A1 => n11183, A2 => n9535, B1 => n11169, B2 => 
                           n9727, ZN => n15175);
   U2842 : AOI22_X1 port map( A1 => n11171, A2 => n9567, B1 => n11161, B2 => 
                           n9631, ZN => n15174);
   U2843 : NAND4_X1 port map( A1 => n15177, A2 => n15176, A3 => n15175, A4 => 
                           n15174, ZN => n15178);
   U2844 : AOI22_X1 port map( A1 => n15360, A2 => n15179, B1 => n15358, B2 => 
                           n15178, ZN => n15180);
   U2845 : OAI21_X1 port map( B1 => n15182, B2 => n15181, A => n15180, ZN => 
                           OUT2(8));
   U2846 : AOI22_X1 port map( A1 => n10068, A2 => n9182, B1 => n11166, B2 => 
                           n9214, ZN => n15186);
   U2847 : AOI22_X1 port map( A1 => n10063, A2 => n9278, B1 => n11188, B2 => 
                           n9342, ZN => n15185);
   U2848 : AOI22_X1 port map( A1 => n10055, A2 => n9470, B1 => n11172, B2 => 
                           n9150, ZN => n15184);
   U2849 : AOI22_X1 port map( A1 => n11191, A2 => n9022, B1 => n10062, B2 => 
                           n9502, ZN => n15183);
   U2850 : NAND4_X1 port map( A1 => n15186, A2 => n15185, A3 => n15184, A4 => 
                           n15183, ZN => n15192);
   U2851 : AOI22_X1 port map( A1 => n11190, A2 => n9118, B1 => n10056, B2 => 
                           n9310, ZN => n15190);
   U2852 : AOI22_X1 port map( A1 => n11189, A2 => n9086, B1 => n10066, B2 => 
                           n9438, ZN => n15189);
   U2853 : AOI22_X1 port map( A1 => n10070, A2 => n9374, B1 => n10057, B2 => 
                           n9406, ZN => n15188);
   U2854 : AOI22_X1 port map( A1 => n11174, A2 => n9054, B1 => n11157, B2 => 
                           n9246, ZN => n15187);
   U2855 : NAND4_X1 port map( A1 => n15190, A2 => n15189, A3 => n15188, A4 => 
                           n15187, ZN => n15191);
   U2856 : NOR2_X1 port map( A1 => n15192, A2 => n15191, ZN => n15204);
   U2857 : AOI22_X1 port map( A1 => n11182, A2 => n9886, B1 => n11179, B2 => 
                           n9790, ZN => n15196);
   U2858 : AOI22_X1 port map( A1 => n11164, A2 => n9854, B1 => n11158, B2 => 
                           n10014, ZN => n15195);
   U2859 : AOI22_X1 port map( A1 => n11181, A2 => n9982, B1 => n11160, B2 => 
                           n9822, ZN => n15194);
   U2860 : AOI22_X1 port map( A1 => n15325, A2 => n9950, B1 => n11185, B2 => 
                           n9918, ZN => n15193);
   U2861 : NAND4_X1 port map( A1 => n15196, A2 => n15195, A3 => n15194, A4 => 
                           n15193, ZN => n15202);
   U2862 : AOI22_X1 port map( A1 => n11169, A2 => n9726, B1 => n11158, B2 => 
                           n9758, ZN => n15200);
   U2863 : AOI22_X1 port map( A1 => n11160, A2 => n9566, B1 => n11159, B2 => 
                           n9662, ZN => n15199);
   U2864 : AOI22_X1 port map( A1 => n11179, A2 => n9534, B1 => n11164, B2 => 
                           n9598, ZN => n15198);
   U2865 : AOI22_X1 port map( A1 => n11226, A2 => n9694, B1 => n11182, B2 => 
                           n9630, ZN => n15197);
   U2866 : NAND4_X1 port map( A1 => n15200, A2 => n15199, A3 => n15198, A4 => 
                           n15197, ZN => n15201);
   U2867 : AOI22_X1 port map( A1 => n15360, A2 => n15202, B1 => n15358, B2 => 
                           n15201, ZN => n15203);
   U2868 : OAI21_X1 port map( B1 => n15363, B2 => n15204, A => n15203, ZN => 
                           OUT2(7));
   U2869 : AOI22_X1 port map( A1 => n10064, A2 => n9213, B1 => n10068, B2 => 
                           n9181, ZN => n15208);
   U2870 : AOI22_X1 port map( A1 => n11190, A2 => n9117, B1 => n11172, B2 => 
                           n9149, ZN => n15207);
   U2871 : AOI22_X1 port map( A1 => n11191, A2 => n9021, B1 => n10069, B2 => 
                           n9053, ZN => n15206);
   U2872 : AOI22_X1 port map( A1 => n11175, A2 => n9373, B1 => n11157, B2 => 
                           n9245, ZN => n15205);
   U2873 : NAND4_X1 port map( A1 => n15208, A2 => n15207, A3 => n15206, A4 => 
                           n15205, ZN => n15214);
   U2874 : AOI22_X1 port map( A1 => n11187, A2 => n9405, B1 => n10056, B2 => 
                           n9309, ZN => n15212);
   U2875 : AOI22_X1 port map( A1 => n10062, A2 => n9501, B1 => n10058, B2 => 
                           n9341, ZN => n15211);
   U2876 : AOI22_X1 port map( A1 => n11189, A2 => n9085, B1 => n11162, B2 => 
                           n9469, ZN => n15210);
   U2877 : AOI22_X1 port map( A1 => n10066, A2 => n9437, B1 => n11165, B2 => 
                           n9277, ZN => n15209);
   U2878 : NAND4_X1 port map( A1 => n15212, A2 => n15211, A3 => n15210, A4 => 
                           n15209, ZN => n15213);
   U2879 : NOR2_X1 port map( A1 => n15214, A2 => n15213, ZN => n15226);
   U2880 : AOI22_X1 port map( A1 => n11184, A2 => n9821, B1 => n11158, B2 => 
                           n10013, ZN => n15218);
   U2881 : AOI22_X1 port map( A1 => n11177, A2 => n9853, B1 => n11159, B2 => 
                           n9917, ZN => n15217);
   U2882 : AOI22_X1 port map( A1 => n11226, A2 => n9949, B1 => n11182, B2 => 
                           n9885, ZN => n15216);
   U2883 : AOI22_X1 port map( A1 => n11181, A2 => n9981, B1 => n11179, B2 => 
                           n9789, ZN => n15215);
   U2884 : NAND4_X1 port map( A1 => n15218, A2 => n15217, A3 => n15216, A4 => 
                           n15215, ZN => n15224);
   U2885 : AOI22_X1 port map( A1 => n15325, A2 => n9693, B1 => n11164, B2 => 
                           n9597, ZN => n15222);
   U2886 : AOI22_X1 port map( A1 => n11160, A2 => n9565, B1 => n11158, B2 => 
                           n9757, ZN => n15221);
   U2887 : AOI22_X1 port map( A1 => n11182, A2 => n9629, B1 => n11170, B2 => 
                           n9661, ZN => n15220);
   U2888 : AOI22_X1 port map( A1 => n11181, A2 => n9725, B1 => n11179, B2 => 
                           n9533, ZN => n15219);
   U2889 : NAND4_X1 port map( A1 => n15222, A2 => n15221, A3 => n15220, A4 => 
                           n15219, ZN => n15223);
   U2890 : AOI22_X1 port map( A1 => n15360, A2 => n15224, B1 => n15358, B2 => 
                           n15223, ZN => n15225);
   U2891 : OAI21_X1 port map( B1 => n15363, B2 => n15226, A => n15225, ZN => 
                           OUT2(6));
   U2892 : AOI22_X1 port map( A1 => n11186, A2 => n9308, B1 => n11165, B2 => 
                           n9276, ZN => n15230);
   U2893 : AOI22_X1 port map( A1 => n11174, A2 => n9052, B1 => n11157, B2 => 
                           n9244, ZN => n15229);
   U2894 : AOI22_X1 port map( A1 => n10066, A2 => n9436, B1 => n10059, B2 => 
                           n9084, ZN => n15228);
   U2895 : AOI22_X1 port map( A1 => n10055, A2 => n9468, B1 => n10058, B2 => 
                           n9340, ZN => n15227);
   U2896 : NAND4_X1 port map( A1 => n15230, A2 => n15229, A3 => n15228, A4 => 
                           n15227, ZN => n15236);
   U2897 : AOI22_X1 port map( A1 => n11191, A2 => n9020, B1 => n10062, B2 => 
                           n9500, ZN => n15234);
   U2898 : AOI22_X1 port map( A1 => n10070, A2 => n9372, B1 => n10061, B2 => 
                           n9116, ZN => n15233);
   U2899 : AOI22_X1 port map( A1 => n10064, A2 => n9212, B1 => n11172, B2 => 
                           n9148, ZN => n15232);
   U2900 : AOI22_X1 port map( A1 => n11187, A2 => n9404, B1 => n11173, B2 => 
                           n9180, ZN => n15231);
   U2901 : NAND4_X1 port map( A1 => n15234, A2 => n15233, A3 => n15232, A4 => 
                           n15231, ZN => n15235);
   U2902 : NOR2_X1 port map( A1 => n15236, A2 => n15235, ZN => n15248);
   U2903 : AOI22_X1 port map( A1 => n11161, A2 => n9884, B1 => n11158, B2 => 
                           n10012, ZN => n15240);
   U2904 : AOI22_X1 port map( A1 => n11169, A2 => n9980, B1 => n11164, B2 => 
                           n9852, ZN => n15239);
   U2905 : AOI22_X1 port map( A1 => n11179, A2 => n9788, B1 => n11160, B2 => 
                           n9820, ZN => n15238);
   U2906 : AOI22_X1 port map( A1 => n15325, A2 => n9948, B1 => n11159, B2 => 
                           n9916, ZN => n15237);
   U2907 : NAND4_X1 port map( A1 => n15240, A2 => n15239, A3 => n15238, A4 => 
                           n15237, ZN => n15246);
   U2908 : AOI22_X1 port map( A1 => n11184, A2 => n9564, B1 => n11170, B2 => 
                           n9660, ZN => n15244);
   U2909 : AOI22_X1 port map( A1 => n11164, A2 => n9596, B1 => n11158, B2 => 
                           n9756, ZN => n15243);
   U2910 : AOI22_X1 port map( A1 => n11226, A2 => n9692, B1 => n11179, B2 => 
                           n9532, ZN => n15242);
   U2911 : AOI22_X1 port map( A1 => n11176, A2 => n9724, B1 => n11161, B2 => 
                           n9628, ZN => n15241);
   U2912 : NAND4_X1 port map( A1 => n15244, A2 => n15243, A3 => n15242, A4 => 
                           n15241, ZN => n15245);
   U2913 : AOI22_X1 port map( A1 => n15360, A2 => n15246, B1 => n15358, B2 => 
                           n15245, ZN => n15247);
   U2914 : OAI21_X1 port map( B1 => n15363, B2 => n15248, A => n15247, ZN => 
                           OUT2(5));
   U2915 : AOI22_X1 port map( A1 => n10064, A2 => n9211, B1 => n10059, B2 => 
                           n9083, ZN => n15252);
   U2916 : AOI22_X1 port map( A1 => n10062, A2 => n9499, B1 => n11174, B2 => 
                           n9051, ZN => n15251);
   U2917 : AOI22_X1 port map( A1 => n11191, A2 => n9019, B1 => n11165, B2 => 
                           n9275, ZN => n15250);
   U2918 : AOI22_X1 port map( A1 => n10056, A2 => n9307, B1 => n10058, B2 => 
                           n9339, ZN => n15249);
   U2919 : NAND4_X1 port map( A1 => n15252, A2 => n15251, A3 => n15250, A4 => 
                           n15249, ZN => n15258);
   U2920 : AOI22_X1 port map( A1 => n10055, A2 => n9467, B1 => n11157, B2 => 
                           n9243, ZN => n15256);
   U2921 : AOI22_X1 port map( A1 => n10068, A2 => n9179, B1 => n10066, B2 => 
                           n9435, ZN => n15255);
   U2922 : AOI22_X1 port map( A1 => n11187, A2 => n9403, B1 => n11172, B2 => 
                           n9147, ZN => n15254);
   U2923 : AOI22_X1 port map( A1 => n11190, A2 => n9115, B1 => n11175, B2 => 
                           n9371, ZN => n15253);
   U2924 : NAND4_X1 port map( A1 => n15256, A2 => n15255, A3 => n15254, A4 => 
                           n15253, ZN => n15257);
   U2925 : NOR2_X1 port map( A1 => n15258, A2 => n15257, ZN => n15270);
   U2926 : AOI22_X1 port map( A1 => n11181, A2 => n9979, B1 => n11158, B2 => 
                           n10011, ZN => n15262);
   U2927 : AOI22_X1 port map( A1 => n11182, A2 => n9883, B1 => n11164, B2 => 
                           n9851, ZN => n15261);
   U2928 : AOI22_X1 port map( A1 => n11171, A2 => n9819, B1 => n11159, B2 => 
                           n9915, ZN => n15260);
   U2929 : AOI22_X1 port map( A1 => n11226, A2 => n9947, B1 => n11179, B2 => 
                           n9787, ZN => n15259);
   U2930 : NAND4_X1 port map( A1 => n15262, A2 => n15261, A3 => n15260, A4 => 
                           n15259, ZN => n15268);
   U2931 : AOI22_X1 port map( A1 => n11164, A2 => n9595, B1 => n11160, B2 => 
                           n9563, ZN => n15266);
   U2932 : AOI22_X1 port map( A1 => n11176, A2 => n9723, B1 => n11158, B2 => 
                           n9755, ZN => n15265);
   U2933 : AOI22_X1 port map( A1 => n11226, A2 => n9691, B1 => n11178, B2 => 
                           n9627, ZN => n15264);
   U2934 : AOI22_X1 port map( A1 => n11179, A2 => n9531, B1 => n11170, B2 => 
                           n9659, ZN => n15263);
   U2935 : NAND4_X1 port map( A1 => n15266, A2 => n15265, A3 => n15264, A4 => 
                           n15263, ZN => n15267);
   U2936 : AOI22_X1 port map( A1 => n15360, A2 => n15268, B1 => n15358, B2 => 
                           n15267, ZN => n15269);
   U2937 : OAI21_X1 port map( B1 => n15363, B2 => n15270, A => n15269, ZN => 
                           OUT2(4));
   U2938 : AOI22_X1 port map( A1 => n11186, A2 => n9306, B1 => n11162, B2 => 
                           n9466, ZN => n15274);
   U2939 : AOI22_X1 port map( A1 => n10063, A2 => n9274, B1 => n10070, B2 => 
                           n9370, ZN => n15273);
   U2940 : AOI22_X1 port map( A1 => n10066, A2 => n9434, B1 => n10057, B2 => 
                           n9402, ZN => n15272);
   U2941 : AOI22_X1 port map( A1 => n11188, A2 => n9338, B1 => n11173, B2 => 
                           n9178, ZN => n15271);
   U2942 : NAND4_X1 port map( A1 => n15274, A2 => n15273, A3 => n15272, A4 => 
                           n15271, ZN => n15280);
   U2943 : AOI22_X1 port map( A1 => n11172, A2 => n9146, B1 => n11157, B2 => 
                           n9242, ZN => n15278);
   U2944 : AOI22_X1 port map( A1 => n11190, A2 => n9114, B1 => n10059, B2 => 
                           n9082, ZN => n15277);
   U2945 : AOI22_X1 port map( A1 => n10062, A2 => n9498, B1 => n10064, B2 => 
                           n9210, ZN => n15276);
   U2946 : AOI22_X1 port map( A1 => n11191, A2 => n9018, B1 => n11174, B2 => 
                           n9050, ZN => n15275);
   U2947 : NAND4_X1 port map( A1 => n15278, A2 => n15277, A3 => n15276, A4 => 
                           n15275, ZN => n15279);
   U2948 : NOR2_X1 port map( A1 => n15280, A2 => n15279, ZN => n15292);
   U2949 : AOI22_X1 port map( A1 => n15325, A2 => n9946, B1 => n11164, B2 => 
                           n9850, ZN => n15284);
   U2950 : AOI22_X1 port map( A1 => n11182, A2 => n9882, B1 => n11179, B2 => 
                           n9786, ZN => n15283);
   U2951 : AOI22_X1 port map( A1 => n11171, A2 => n9818, B1 => n11169, B2 => 
                           n9978, ZN => n15282);
   U2952 : AOI22_X1 port map( A1 => n11170, A2 => n9914, B1 => n11158, B2 => 
                           n10010, ZN => n15281);
   U2953 : NAND4_X1 port map( A1 => n15284, A2 => n15283, A3 => n15282, A4 => 
                           n15281, ZN => n15290);
   U2954 : AOI22_X1 port map( A1 => n11182, A2 => n9626, B1 => n11169, B2 => 
                           n9722, ZN => n15288);
   U2955 : AOI22_X1 port map( A1 => n11177, A2 => n9594, B1 => n11170, B2 => 
                           n9658, ZN => n15287);
   U2956 : AOI22_X1 port map( A1 => n11226, A2 => n9690, B1 => n11158, B2 => 
                           n9754, ZN => n15286);
   U2957 : AOI22_X1 port map( A1 => n11179, A2 => n9530, B1 => n11171, B2 => 
                           n9562, ZN => n15285);
   U2958 : NAND4_X1 port map( A1 => n15288, A2 => n15287, A3 => n15286, A4 => 
                           n15285, ZN => n15289);
   U2959 : AOI22_X1 port map( A1 => n15360, A2 => n15290, B1 => n15358, B2 => 
                           n15289, ZN => n15291);
   U2960 : OAI21_X1 port map( B1 => n15363, B2 => n15292, A => n15291, ZN => 
                           OUT2(3));
   U2961 : AOI22_X1 port map( A1 => n11187, A2 => n9401, B1 => n11157, B2 => 
                           n9241, ZN => n15296);
   U2962 : AOI22_X1 port map( A1 => n10056, A2 => n9305, B1 => n11174, B2 => 
                           n9049, ZN => n15295);
   U2963 : AOI22_X1 port map( A1 => n11191, A2 => n9017, B1 => n10061, B2 => 
                           n9113, ZN => n15294);
   U2964 : AOI22_X1 port map( A1 => n11162, A2 => n9465, B1 => n10059, B2 => 
                           n9081, ZN => n15293);
   U2965 : NAND4_X1 port map( A1 => n15296, A2 => n15295, A3 => n15294, A4 => 
                           n15293, ZN => n15302);
   U2966 : AOI22_X1 port map( A1 => n10062, A2 => n9497, B1 => n11165, B2 => 
                           n9273, ZN => n15300);
   U2967 : AOI22_X1 port map( A1 => n11175, A2 => n9369, B1 => n11166, B2 => 
                           n9209, ZN => n15299);
   U2968 : AOI22_X1 port map( A1 => n11188, A2 => n9337, B1 => n10066, B2 => 
                           n9433, ZN => n15298);
   U2969 : AOI22_X1 port map( A1 => n11172, A2 => n9145, B1 => n11173, B2 => 
                           n9177, ZN => n15297);
   U2970 : NAND4_X1 port map( A1 => n15300, A2 => n15299, A3 => n15298, A4 => 
                           n15297, ZN => n15301);
   U2971 : NOR2_X1 port map( A1 => n15302, A2 => n15301, ZN => n15314);
   U2972 : AOI22_X1 port map( A1 => n11171, A2 => n9817, B1 => n11161, B2 => 
                           n9881, ZN => n15306);
   U2973 : AOI22_X1 port map( A1 => n11170, A2 => n9913, B1 => n11158, B2 => 
                           n10009, ZN => n15305);
   U2974 : AOI22_X1 port map( A1 => n11179, A2 => n9785, B1 => n11169, B2 => 
                           n9977, ZN => n15304);
   U2975 : AOI22_X1 port map( A1 => n15325, A2 => n9945, B1 => n11164, B2 => 
                           n9849, ZN => n15303);
   U2976 : NAND4_X1 port map( A1 => n15306, A2 => n15305, A3 => n15304, A4 => 
                           n15303, ZN => n15312);
   U2977 : AOI22_X1 port map( A1 => n11184, A2 => n9561, B1 => n11170, B2 => 
                           n9657, ZN => n15310);
   U2978 : AOI22_X1 port map( A1 => n11179, A2 => n9529, B1 => n11158, B2 => 
                           n9753, ZN => n15309);
   U2979 : AOI22_X1 port map( A1 => n11226, A2 => n9689, B1 => n11161, B2 => 
                           n9625, ZN => n15308);
   U2980 : AOI22_X1 port map( A1 => n11169, A2 => n9721, B1 => n11164, B2 => 
                           n9593, ZN => n15307);
   U2981 : NAND4_X1 port map( A1 => n15310, A2 => n15309, A3 => n15308, A4 => 
                           n15307, ZN => n15311);
   U2982 : AOI22_X1 port map( A1 => n15360, A2 => n15312, B1 => n15358, B2 => 
                           n15311, ZN => n15313);
   U2983 : OAI21_X1 port map( B1 => n15363, B2 => n15314, A => n15313, ZN => 
                           OUT2(2));
   U2984 : AOI22_X1 port map( A1 => n10066, A2 => n9432, B1 => n11173, B2 => 
                           n9176, ZN => n15318);
   U2985 : AOI22_X1 port map( A1 => n10056, A2 => n9304, B1 => n11157, B2 => 
                           n9240, ZN => n15317);
   U2986 : AOI22_X1 port map( A1 => n11174, A2 => n9048, B1 => n11167, B2 => 
                           n9496, ZN => n15316);
   U2987 : AOI22_X1 port map( A1 => n11189, A2 => n9080, B1 => n10057, B2 => 
                           n9400, ZN => n15315);
   U2988 : NAND4_X1 port map( A1 => n15318, A2 => n15317, A3 => n15316, A4 => 
                           n15315, ZN => n15324);
   U2989 : AOI22_X1 port map( A1 => n10063, A2 => n9272, B1 => n11166, B2 => 
                           n9208, ZN => n15322);
   U2990 : AOI22_X1 port map( A1 => n10058, A2 => n9336, B1 => n10061, B2 => 
                           n9112, ZN => n15321);
   U2991 : AOI22_X1 port map( A1 => n11172, A2 => n9144, B1 => n11162, B2 => 
                           n9464, ZN => n15320);
   U2992 : AOI22_X1 port map( A1 => n11191, A2 => n9016, B1 => n10070, B2 => 
                           n9368, ZN => n15319);
   U2993 : NAND4_X1 port map( A1 => n15322, A2 => n15321, A3 => n15320, A4 => 
                           n15319, ZN => n15323);
   U2994 : NOR2_X1 port map( A1 => n15324, A2 => n15323, ZN => n15337);
   U2995 : AOI22_X1 port map( A1 => n11171, A2 => n9816, B1 => n11170, B2 => 
                           n9912, ZN => n15329);
   U2996 : AOI22_X1 port map( A1 => n11183, A2 => n9784, B1 => n11158, B2 => 
                           n10008, ZN => n15328);
   U2997 : AOI22_X1 port map( A1 => n15325, A2 => n9944, B1 => n11164, B2 => 
                           n9848, ZN => n15327);
   U2998 : AOI22_X1 port map( A1 => n11182, A2 => n9880, B1 => n11169, B2 => 
                           n9976, ZN => n15326);
   U2999 : NAND4_X1 port map( A1 => n15329, A2 => n15328, A3 => n15327, A4 => 
                           n15326, ZN => n15335);
   U3000 : AOI22_X1 port map( A1 => n11181, A2 => n9720, B1 => n11179, B2 => 
                           n9528, ZN => n15333);
   U3001 : AOI22_X1 port map( A1 => n11227, A2 => n9752, B1 => n11160, B2 => 
                           n9560, ZN => n15332);
   U3002 : AOI22_X1 port map( A1 => n11182, A2 => n9624, B1 => n11156, B2 => 
                           n9688, ZN => n15331);
   U3003 : AOI22_X1 port map( A1 => n11164, A2 => n9592, B1 => n11159, B2 => 
                           n9656, ZN => n15330);
   U3004 : NAND4_X1 port map( A1 => n15333, A2 => n15332, A3 => n15331, A4 => 
                           n15330, ZN => n15334);
   U3005 : AOI22_X1 port map( A1 => n15360, A2 => n15335, B1 => n15358, B2 => 
                           n15334, ZN => n15336);
   U3006 : OAI21_X1 port map( B1 => n15363, B2 => n15337, A => n15336, ZN => 
                           OUT2(1));
   U3007 : AOI22_X1 port map( A1 => n10070, A2 => n9367, B1 => n11166, B2 => 
                           n9207, ZN => n15341);
   U3008 : AOI22_X1 port map( A1 => n11188, A2 => n9335, B1 => n11162, B2 => 
                           n9463, ZN => n15340);
   U3009 : AOI22_X1 port map( A1 => n11186, A2 => n9303, B1 => n11190, B2 => 
                           n9111, ZN => n15339);
   U3010 : AOI22_X1 port map( A1 => n11189, A2 => n9079, B1 => n11174, B2 => 
                           n9047, ZN => n15338);
   U3011 : NAND4_X1 port map( A1 => n15341, A2 => n15340, A3 => n15339, A4 => 
                           n15338, ZN => n15347);
   U3012 : AOI22_X1 port map( A1 => n10063, A2 => n9271, B1 => n11167, B2 => 
                           n9495, ZN => n15345);
   U3013 : AOI22_X1 port map( A1 => n11172, A2 => n9143, B1 => n11168, B2 => 
                           n9431, ZN => n15344);
   U3014 : AOI22_X1 port map( A1 => n11191, A2 => n9015, B1 => n11157, B2 => 
                           n9239, ZN => n15343);
   U3015 : AOI22_X1 port map( A1 => n11173, A2 => n9175, B1 => n10057, B2 => 
                           n9399, ZN => n15342);
   U3016 : NAND4_X1 port map( A1 => n15345, A2 => n15344, A3 => n15343, A4 => 
                           n15342, ZN => n15346);
   U3017 : NOR2_X1 port map( A1 => n15347, A2 => n15346, ZN => n15362);
   U3018 : AOI22_X1 port map( A1 => n11181, A2 => n9975, B1 => n11184, B2 => 
                           n9815, ZN => n15351);
   U3019 : AOI22_X1 port map( A1 => n11226, A2 => n9943, B1 => n11158, B2 => 
                           n10007, ZN => n15350);
   U3020 : AOI22_X1 port map( A1 => n11182, A2 => n9879, B1 => n11164, B2 => 
                           n9847, ZN => n15349);
   U3021 : AOI22_X1 port map( A1 => n11179, A2 => n9783, B1 => n11170, B2 => 
                           n9911, ZN => n15348);
   U3022 : NAND4_X1 port map( A1 => n15351, A2 => n15350, A3 => n15349, A4 => 
                           n15348, ZN => n15359);
   U3023 : AOI22_X1 port map( A1 => n11182, A2 => n9623, B1 => n11183, B2 => 
                           n9527, ZN => n15356);
   U3024 : AOI22_X1 port map( A1 => n11171, A2 => n9559, B1 => n11159, B2 => 
                           n9655, ZN => n15355);
   U3025 : AOI22_X1 port map( A1 => n11169, A2 => n9719, B1 => n11156, B2 => 
                           n9687, ZN => n15354);
   U3026 : AOI22_X1 port map( A1 => n15352, A2 => n9751, B1 => n11177, B2 => 
                           n9591, ZN => n15353);
   U3027 : NAND4_X1 port map( A1 => n15356, A2 => n15355, A3 => n15354, A4 => 
                           n15353, ZN => n15357);
   U3028 : AOI22_X1 port map( A1 => n15360, A2 => n15359, B1 => n15358, B2 => 
                           n15357, ZN => n15361);
   U3029 : OAI21_X1 port map( B1 => n15363, B2 => n15362, A => n15361, ZN => 
                           OUT2(0));
   U3030 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n15373)
                           ;
   U3031 : INV_X1 port map( A => n3579, ZN => n15364);
   U3032 : NOR2_X1 port map( A1 => n15373, A2 => n15364, ZN => n5699);
   U3033 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n3574, ZN => n15369);
   U3034 : INV_X1 port map( A => n3578, ZN => n15366);
   U3035 : NOR2_X1 port map( A1 => n15369, A2 => n15366, ZN => n5599);
   U3036 : NOR2_X1 port map( A1 => n15364, A2 => n15369, ZN => n5700);
   U3037 : INV_X1 port map( A => n3580, ZN => n15365);
   U3038 : NOR2_X1 port map( A1 => n15373, A2 => n15365, ZN => n5688);
   U3039 : INV_X1 port map( A => n3581, ZN => n15371);
   U3040 : NOR2_X1 port map( A1 => n15369, A2 => n15371, ZN => n5654);
   U3041 : INV_X1 port map( A => n3582, ZN => n15367);
   U3042 : NOR2_X1 port map( A1 => n15369, A2 => n15367, ZN => n5697);
   U3043 : INV_X1 port map( A => n3577, ZN => n15370);
   U3044 : NOR2_X1 port map( A1 => n15369, A2 => n15370, ZN => n5686);
   U3045 : NOR2_X1 port map( A1 => n15369, A2 => n15365, ZN => n5645);
   U3046 : NOR2_X1 port map( A1 => n15373, A2 => n15366, ZN => n5648);
   U3047 : NOR2_X1 port map( A1 => n15373, A2 => n15367, ZN => n5624);
   U3048 : INV_X1 port map( A => n3576, ZN => n15368);
   U3049 : NOR2_X1 port map( A1 => n15369, A2 => n15368, ZN => n5594);
   U3050 : NOR2_X1 port map( A1 => n15373, A2 => n15368, ZN => n5696);
   U3051 : INV_X1 port map( A => n3575, ZN => n15372);
   U3052 : NOR2_X1 port map( A1 => n15369, A2 => n15372, ZN => n5570);
   U3053 : NOR2_X1 port map( A1 => n15373, A2 => n15370, ZN => n5694);
   U3054 : NOR2_X1 port map( A1 => n15373, A2 => n15371, ZN => n5655);
   U3055 : NOR2_X1 port map( A1 => n15373, A2 => n15372, ZN => n5625);
   U3056 : AOI22_X1 port map( A1 => n9110, A2 => n10040, B1 => n9462, B2 => 
                           n11151, ZN => n15377);
   U3057 : AOI22_X1 port map( A1 => n9174, A2 => n10041, B1 => n9526, B2 => 
                           n10052, ZN => n15376);
   U3058 : AOI22_X1 port map( A1 => n9238, A2 => n10039, B1 => n9206, B2 => 
                           n11153, ZN => n15375);
   U3059 : AOI22_X1 port map( A1 => n9494, A2 => n10042, B1 => n9334, B2 => 
                           n10044, ZN => n15374);
   U3060 : NAND4_X1 port map( A1 => n15377, A2 => n15376, A3 => n15375, A4 => 
                           n15374, ZN => n15383);
   U3061 : AOI22_X1 port map( A1 => n9046, A2 => n11150, B1 => n9430, B2 => 
                           n10048, ZN => n15381);
   U3062 : AOI22_X1 port map( A1 => n9270, A2 => n10054, B1 => n9398, B2 => 
                           n11154, ZN => n15380);
   U3063 : AOI22_X1 port map( A1 => n9078, A2 => n11149, B1 => n9142, B2 => 
                           n10046, ZN => n15379);
   U3064 : AOI22_X1 port map( A1 => n9302, A2 => n11152, B1 => n9366, B2 => 
                           n10050, ZN => n15378);
   U3065 : NAND4_X1 port map( A1 => n15381, A2 => n15380, A3 => n15379, A4 => 
                           n15378, ZN => n15382);
   U3066 : NOR2_X1 port map( A1 => n15383, A2 => n15382, ZN => n15395);
   U3067 : NOR3_X1 port map( A1 => n11267, A2 => n11268, A3 => n15905, ZN => 
                           n15835);
   U3068 : CLKBUF_X1 port map( A => n15835, Z => n15880);
   U3069 : AOI22_X1 port map( A1 => n10006, A2 => n11228, B1 => n9910, B2 => 
                           n11148, ZN => n15387);
   U3070 : AOI22_X1 port map( A1 => n9878, A2 => n11229, B1 => n9942, B2 => 
                           n11232, ZN => n15386);
   U3071 : CLKBUF_X1 port map( A => n11231, Z => n16072);
   U3072 : AOI22_X1 port map( A1 => n10038, A2 => n16072, B1 => n9846, B2 => 
                           n11147, ZN => n15385);
   U3073 : CLKBUF_X1 port map( A => n11230, Z => n16048);
   U3074 : AOI22_X1 port map( A1 => n9974, A2 => n16048, B1 => n9814, B2 => 
                           n11225, ZN => n15384);
   U3075 : NAND4_X1 port map( A1 => n15387, A2 => n15386, A3 => n15385, A4 => 
                           n15384, ZN => n15393);
   U3076 : NOR3_X1 port map( A1 => n11268, A2 => n11155, A3 => n15905, ZN => 
                           n15613);
   U3077 : CLKBUF_X1 port map( A => n15613, Z => n16085);
   U3078 : CLKBUF_X1 port map( A => n11225, Z => n16077);
   U3079 : CLKBUF_X1 port map( A => n11232, Z => n16079);
   U3080 : AOI22_X1 port map( A1 => n9558, A2 => n16077, B1 => n9686, B2 => 
                           n16079, ZN => n15391);
   U3081 : AOI22_X1 port map( A1 => n9622, A2 => n11229, B1 => n9782, B2 => 
                           n11146, ZN => n15390);
   U3082 : AOI22_X1 port map( A1 => n9750, A2 => n11228, B1 => n9654, B2 => 
                           n11144, ZN => n15389);
   U3083 : AOI22_X1 port map( A1 => n9718, A2 => n11230, B1 => n9590, B2 => 
                           n11145, ZN => n15388);
   U3084 : NAND4_X1 port map( A1 => n15391, A2 => n15390, A3 => n15389, A4 => 
                           n15388, ZN => n15392);
   U3085 : AOI22_X1 port map( A1 => n15880, A2 => n15393, B1 => n16085, B2 => 
                           n15392, ZN => n15394);
   U3086 : OAI21_X1 port map( B1 => n15905, B2 => n15395, A => n15394, ZN => 
                           OUT1(31));
   U3087 : AOI22_X1 port map( A1 => n9493, A2 => n10042, B1 => n9045, B2 => 
                           n11150, ZN => n15399);
   U3088 : AOI22_X1 port map( A1 => n9525, A2 => n11136, B1 => n9109, B2 => 
                           n11142, ZN => n15398);
   U3089 : AOI22_X1 port map( A1 => n9461, A2 => n11151, B1 => n9237, B2 => 
                           n11143, ZN => n15397);
   U3090 : AOI22_X1 port map( A1 => n9173, A2 => n11140, B1 => n9333, B2 => 
                           n11138, ZN => n15396);
   U3091 : NAND4_X1 port map( A1 => n15399, A2 => n15398, A3 => n15397, A4 => 
                           n15396, ZN => n15405);
   U3092 : AOI22_X1 port map( A1 => n9365, A2 => n11139, B1 => n9429, B2 => 
                           n11141, ZN => n15403);
   U3093 : AOI22_X1 port map( A1 => n9269, A2 => n10054, B1 => n9077, B2 => 
                           n10043, ZN => n15402);
   U3094 : AOI22_X1 port map( A1 => n9141, A2 => n11137, B1 => n9205, B2 => 
                           n10051, ZN => n15401);
   U3095 : AOI22_X1 port map( A1 => n9301, A2 => n11152, B1 => n9397, B2 => 
                           n11154, ZN => n15400);
   U3096 : NAND4_X1 port map( A1 => n15403, A2 => n15402, A3 => n15401, A4 => 
                           n15400, ZN => n15404);
   U3097 : NOR2_X1 port map( A1 => n15405, A2 => n15404, ZN => n15417);
   U3098 : CLKBUF_X1 port map( A => n11228, Z => n16053);
   U3099 : AOI22_X1 port map( A1 => n10005, A2 => n16053, B1 => n9909, B2 => 
                           n11148, ZN => n15409);
   U3100 : AOI22_X1 port map( A1 => n9845, A2 => n11147, B1 => n9941, B2 => 
                           n11135, ZN => n15408);
   U3101 : AOI22_X1 port map( A1 => n9877, A2 => n11229, B1 => n10037, B2 => 
                           n11146, ZN => n15407);
   U3102 : AOI22_X1 port map( A1 => n9973, A2 => n16048, B1 => n9813, B2 => 
                           n11225, ZN => n15406);
   U3103 : NAND4_X1 port map( A1 => n15409, A2 => n15408, A3 => n15407, A4 => 
                           n15406, ZN => n15415);
   U3104 : AOI22_X1 port map( A1 => n9685, A2 => n11135, B1 => n9653, B2 => 
                           n11148, ZN => n15413);
   U3105 : AOI22_X1 port map( A1 => n9749, A2 => n11228, B1 => n9589, B2 => 
                           n11147, ZN => n15412);
   U3106 : AOI22_X1 port map( A1 => n9557, A2 => n11134, B1 => n9781, B2 => 
                           n11231, ZN => n15411);
   U3107 : AOI22_X1 port map( A1 => n9717, A2 => n11230, B1 => n9621, B2 => 
                           n11229, ZN => n15410);
   U3108 : NAND4_X1 port map( A1 => n15413, A2 => n15412, A3 => n15411, A4 => 
                           n15410, ZN => n15414);
   U3109 : AOI22_X1 port map( A1 => n15880, A2 => n15415, B1 => n16085, B2 => 
                           n15414, ZN => n15416);
   U3110 : OAI21_X1 port map( B1 => n15905, B2 => n15417, A => n15416, ZN => 
                           OUT1(30));
   U3111 : AOI22_X1 port map( A1 => n9396, A2 => n11154, B1 => n9076, B2 => 
                           n11149, ZN => n15421);
   U3112 : AOI22_X1 port map( A1 => n9364, A2 => n11139, B1 => n9460, B2 => 
                           n11151, ZN => n15420);
   U3113 : AOI22_X1 port map( A1 => n9492, A2 => n11133, B1 => n9108, B2 => 
                           n11142, ZN => n15419);
   U3114 : AOI22_X1 port map( A1 => n9236, A2 => n11143, B1 => n9300, B2 => 
                           n10049, ZN => n15418);
   U3115 : NAND4_X1 port map( A1 => n15421, A2 => n15420, A3 => n15419, A4 => 
                           n15418, ZN => n15427);
   U3116 : AOI22_X1 port map( A1 => n9044, A2 => n11150, B1 => n9332, B2 => 
                           n11138, ZN => n15425);
   U3117 : AOI22_X1 port map( A1 => n9204, A2 => n11153, B1 => n9524, B2 => 
                           n11136, ZN => n15424);
   U3118 : AOI22_X1 port map( A1 => n9428, A2 => n11141, B1 => n9268, B2 => 
                           n11132, ZN => n15423);
   U3119 : AOI22_X1 port map( A1 => n9140, A2 => n11137, B1 => n9172, B2 => 
                           n10041, ZN => n15422);
   U3120 : NAND4_X1 port map( A1 => n15425, A2 => n15424, A3 => n15423, A4 => 
                           n15422, ZN => n15426);
   U3121 : NOR2_X1 port map( A1 => n15427, A2 => n15426, ZN => n15439);
   U3122 : AOI22_X1 port map( A1 => n9972, A2 => n16048, B1 => n9844, B2 => 
                           n11145, ZN => n15431);
   U3123 : AOI22_X1 port map( A1 => n9876, A2 => n11131, B1 => n9940, B2 => 
                           n11232, ZN => n15430);
   U3124 : AOI22_X1 port map( A1 => n10036, A2 => n16072, B1 => n9812, B2 => 
                           n16077, ZN => n15429);
   U3125 : AOI22_X1 port map( A1 => n9908, A2 => n11148, B1 => n10004, B2 => 
                           n11130, ZN => n15428);
   U3126 : NAND4_X1 port map( A1 => n15431, A2 => n15430, A3 => n15429, A4 => 
                           n15428, ZN => n15437);
   U3127 : AOI22_X1 port map( A1 => n9748, A2 => n11130, B1 => n9716, B2 => 
                           n11129, ZN => n15435);
   U3128 : AOI22_X1 port map( A1 => n9780, A2 => n11231, B1 => n9652, B2 => 
                           n11144, ZN => n15434);
   U3129 : AOI22_X1 port map( A1 => n9556, A2 => n11134, B1 => n9620, B2 => 
                           n11229, ZN => n15433);
   U3130 : AOI22_X1 port map( A1 => n9588, A2 => n11147, B1 => n9684, B2 => 
                           n16079, ZN => n15432);
   U3131 : NAND4_X1 port map( A1 => n15435, A2 => n15434, A3 => n15433, A4 => 
                           n15432, ZN => n15436);
   U3132 : AOI22_X1 port map( A1 => n15880, A2 => n15437, B1 => n16085, B2 => 
                           n15436, ZN => n15438);
   U3133 : OAI21_X1 port map( B1 => n15905, B2 => n15439, A => n15438, ZN => 
                           OUT1(29));
   U3134 : AOI22_X1 port map( A1 => n9395, A2 => n10053, B1 => n9523, B2 => 
                           n11136, ZN => n15443);
   U3135 : AOI22_X1 port map( A1 => n9235, A2 => n11143, B1 => n9299, B2 => 
                           n10049, ZN => n15442);
   U3136 : AOI22_X1 port map( A1 => n9427, A2 => n11141, B1 => n9363, B2 => 
                           n11139, ZN => n15441);
   U3137 : AOI22_X1 port map( A1 => n9043, A2 => n11150, B1 => n9331, B2 => 
                           n11138, ZN => n15440);
   U3138 : NAND4_X1 port map( A1 => n15443, A2 => n15442, A3 => n15441, A4 => 
                           n15440, ZN => n15449);
   U3139 : AOI22_X1 port map( A1 => n9171, A2 => n10041, B1 => n9491, B2 => 
                           n10042, ZN => n15447);
   U3140 : AOI22_X1 port map( A1 => n9459, A2 => n11151, B1 => n9075, B2 => 
                           n10043, ZN => n15446);
   U3141 : AOI22_X1 port map( A1 => n9203, A2 => n11153, B1 => n9139, B2 => 
                           n11137, ZN => n15445);
   U3142 : AOI22_X1 port map( A1 => n9107, A2 => n11142, B1 => n9267, B2 => 
                           n10054, ZN => n15444);
   U3143 : NAND4_X1 port map( A1 => n15447, A2 => n15446, A3 => n15445, A4 => 
                           n15444, ZN => n15448);
   U3144 : NOR2_X1 port map( A1 => n15449, A2 => n15448, ZN => n15461);
   U3145 : AOI22_X1 port map( A1 => n10035, A2 => n11231, B1 => n9907, B2 => 
                           n11128, ZN => n15453);
   U3146 : AOI22_X1 port map( A1 => n9939, A2 => n11232, B1 => n9811, B2 => 
                           n16077, ZN => n15452);
   U3147 : CLKBUF_X1 port map( A => n11229, Z => n16078);
   U3148 : AOI22_X1 port map( A1 => n9875, A2 => n16078, B1 => n9971, B2 => 
                           n16048, ZN => n15451);
   U3149 : AOI22_X1 port map( A1 => n9843, A2 => n11147, B1 => n10003, B2 => 
                           n11130, ZN => n15450);
   U3150 : NAND4_X1 port map( A1 => n15453, A2 => n15452, A3 => n15451, A4 => 
                           n15450, ZN => n15459);
   U3151 : AOI22_X1 port map( A1 => n9555, A2 => n11225, B1 => n9587, B2 => 
                           n11147, ZN => n15457);
   U3152 : AOI22_X1 port map( A1 => n9715, A2 => n11230, B1 => n9683, B2 => 
                           n11232, ZN => n15456);
   U3153 : AOI22_X1 port map( A1 => n9619, A2 => n11229, B1 => n9779, B2 => 
                           n11146, ZN => n15455);
   U3154 : AOI22_X1 port map( A1 => n9747, A2 => n16053, B1 => n9651, B2 => 
                           n11144, ZN => n15454);
   U3155 : NAND4_X1 port map( A1 => n15457, A2 => n15456, A3 => n15455, A4 => 
                           n15454, ZN => n15458);
   U3156 : AOI22_X1 port map( A1 => n15880, A2 => n15459, B1 => n16085, B2 => 
                           n15458, ZN => n15460);
   U3157 : OAI21_X1 port map( B1 => n15905, B2 => n15461, A => n15460, ZN => 
                           OUT1(28));
   U3158 : AOI22_X1 port map( A1 => n9522, A2 => n11136, B1 => n9234, B2 => 
                           n11143, ZN => n15465);
   U3159 : AOI22_X1 port map( A1 => n9042, A2 => n11150, B1 => n9138, B2 => 
                           n11137, ZN => n15464);
   U3160 : AOI22_X1 port map( A1 => n9426, A2 => n11141, B1 => n9298, B2 => 
                           n10049, ZN => n15463);
   U3161 : AOI22_X1 port map( A1 => n9330, A2 => n11138, B1 => n9202, B2 => 
                           n11153, ZN => n15462);
   U3162 : NAND4_X1 port map( A1 => n15465, A2 => n15464, A3 => n15463, A4 => 
                           n15462, ZN => n15471);
   U3163 : AOI22_X1 port map( A1 => n9170, A2 => n10041, B1 => n9362, B2 => 
                           n11139, ZN => n15469);
   U3164 : AOI22_X1 port map( A1 => n9458, A2 => n11151, B1 => n9394, B2 => 
                           n11154, ZN => n15468);
   U3165 : AOI22_X1 port map( A1 => n9074, A2 => n11149, B1 => n9106, B2 => 
                           n10040, ZN => n15467);
   U3166 : AOI22_X1 port map( A1 => n9266, A2 => n10054, B1 => n9490, B2 => 
                           n11133, ZN => n15466);
   U3167 : NAND4_X1 port map( A1 => n15469, A2 => n15468, A3 => n15467, A4 => 
                           n15466, ZN => n15470);
   U3168 : NOR2_X1 port map( A1 => n15471, A2 => n15470, ZN => n15483);
   U3169 : AOI22_X1 port map( A1 => n10002, A2 => n11228, B1 => n9938, B2 => 
                           n11135, ZN => n15475);
   U3170 : AOI22_X1 port map( A1 => n9906, A2 => n11144, B1 => n10034, B2 => 
                           n11231, ZN => n15474);
   U3171 : AOI22_X1 port map( A1 => n9970, A2 => n16048, B1 => n9842, B2 => 
                           n11127, ZN => n15473);
   U3172 : AOI22_X1 port map( A1 => n9874, A2 => n11131, B1 => n9810, B2 => 
                           n16077, ZN => n15472);
   U3173 : NAND4_X1 port map( A1 => n15475, A2 => n15474, A3 => n15473, A4 => 
                           n15472, ZN => n15481);
   U3174 : AOI22_X1 port map( A1 => n9746, A2 => n11130, B1 => n9650, B2 => 
                           n11128, ZN => n15479);
   U3175 : AOI22_X1 port map( A1 => n9618, A2 => n11131, B1 => n9778, B2 => 
                           n16072, ZN => n15478);
   U3176 : AOI22_X1 port map( A1 => n9554, A2 => n11225, B1 => n9714, B2 => 
                           n11230, ZN => n15477);
   U3177 : AOI22_X1 port map( A1 => n9586, A2 => n11147, B1 => n9682, B2 => 
                           n11232, ZN => n15476);
   U3178 : NAND4_X1 port map( A1 => n15479, A2 => n15478, A3 => n15477, A4 => 
                           n15476, ZN => n15480);
   U3179 : AOI22_X1 port map( A1 => n15880, A2 => n15481, B1 => n15613, B2 => 
                           n15480, ZN => n15482);
   U3180 : OAI21_X1 port map( B1 => n15905, B2 => n15483, A => n15482, ZN => 
                           OUT1(27));
   U3181 : AOI22_X1 port map( A1 => n9201, A2 => n11153, B1 => n9297, B2 => 
                           n11152, ZN => n15487);
   U3182 : AOI22_X1 port map( A1 => n9489, A2 => n10042, B1 => n9041, B2 => 
                           n11150, ZN => n15486);
   U3183 : AOI22_X1 port map( A1 => n9169, A2 => n10041, B1 => n9361, B2 => 
                           n11139, ZN => n15485);
   U3184 : AOI22_X1 port map( A1 => n9521, A2 => n11136, B1 => n9425, B2 => 
                           n11141, ZN => n15484);
   U3185 : NAND4_X1 port map( A1 => n15487, A2 => n15486, A3 => n15485, A4 => 
                           n15484, ZN => n15493);
   U3186 : AOI22_X1 port map( A1 => n9073, A2 => n10043, B1 => n9393, B2 => 
                           n11154, ZN => n15491);
   U3187 : AOI22_X1 port map( A1 => n9265, A2 => n10054, B1 => n9137, B2 => 
                           n11137, ZN => n15490);
   U3188 : AOI22_X1 port map( A1 => n9233, A2 => n11143, B1 => n9105, B2 => 
                           n11142, ZN => n15489);
   U3189 : AOI22_X1 port map( A1 => n9457, A2 => n11151, B1 => n9329, B2 => 
                           n10044, ZN => n15488);
   U3190 : NAND4_X1 port map( A1 => n15491, A2 => n15490, A3 => n15489, A4 => 
                           n15488, ZN => n15492);
   U3191 : NOR2_X1 port map( A1 => n15493, A2 => n15492, ZN => n15505);
   U3192 : AOI22_X1 port map( A1 => n9873, A2 => n11131, B1 => n9841, B2 => 
                           n11147, ZN => n15497);
   U3193 : AOI22_X1 port map( A1 => n10033, A2 => n11231, B1 => n9937, B2 => 
                           n11232, ZN => n15496);
   U3194 : AOI22_X1 port map( A1 => n9969, A2 => n11230, B1 => n9809, B2 => 
                           n11225, ZN => n15495);
   U3195 : AOI22_X1 port map( A1 => n10001, A2 => n11130, B1 => n9905, B2 => 
                           n11128, ZN => n15494);
   U3196 : NAND4_X1 port map( A1 => n15497, A2 => n15496, A3 => n15495, A4 => 
                           n15494, ZN => n15503);
   U3197 : AOI22_X1 port map( A1 => n9777, A2 => n11231, B1 => n9649, B2 => 
                           n11144, ZN => n15501);
   U3198 : AOI22_X1 port map( A1 => n9585, A2 => n11127, B1 => n9713, B2 => 
                           n16048, ZN => n15500);
   U3199 : AOI22_X1 port map( A1 => n9617, A2 => n16078, B1 => n9745, B2 => 
                           n11130, ZN => n15499);
   U3200 : AOI22_X1 port map( A1 => n9681, A2 => n16079, B1 => n9553, B2 => 
                           n11134, ZN => n15498);
   U3201 : NAND4_X1 port map( A1 => n15501, A2 => n15500, A3 => n15499, A4 => 
                           n15498, ZN => n15502);
   U3202 : AOI22_X1 port map( A1 => n15880, A2 => n15503, B1 => n15613, B2 => 
                           n15502, ZN => n15504);
   U3203 : OAI21_X1 port map( B1 => n15905, B2 => n15505, A => n15504, ZN => 
                           OUT1(26));
   U3204 : AOI22_X1 port map( A1 => n9168, A2 => n11140, B1 => n9200, B2 => 
                           n11153, ZN => n15509);
   U3205 : AOI22_X1 port map( A1 => n9456, A2 => n11151, B1 => n9488, B2 => 
                           n10042, ZN => n15508);
   U3206 : AOI22_X1 port map( A1 => n9296, A2 => n11152, B1 => n9136, B2 => 
                           n11137, ZN => n15507);
   U3207 : AOI22_X1 port map( A1 => n9520, A2 => n11136, B1 => n9040, B2 => 
                           n11150, ZN => n15506);
   U3208 : NAND4_X1 port map( A1 => n15509, A2 => n15508, A3 => n15507, A4 => 
                           n15506, ZN => n15515);
   U3209 : AOI22_X1 port map( A1 => n9328, A2 => n10044, B1 => n9392, B2 => 
                           n11154, ZN => n15513);
   U3210 : AOI22_X1 port map( A1 => n9232, A2 => n11143, B1 => n9072, B2 => 
                           n10043, ZN => n15512);
   U3211 : AOI22_X1 port map( A1 => n9424, A2 => n11141, B1 => n9264, B2 => 
                           n11132, ZN => n15511);
   U3212 : AOI22_X1 port map( A1 => n9104, A2 => n11142, B1 => n9360, B2 => 
                           n11139, ZN => n15510);
   U3213 : NAND4_X1 port map( A1 => n15513, A2 => n15512, A3 => n15511, A4 => 
                           n15510, ZN => n15514);
   U3214 : NOR2_X1 port map( A1 => n15515, A2 => n15514, ZN => n15527);
   U3215 : AOI22_X1 port map( A1 => n9904, A2 => n11128, B1 => n9936, B2 => 
                           n16079, ZN => n15519);
   U3216 : AOI22_X1 port map( A1 => n10000, A2 => n11228, B1 => n9968, B2 => 
                           n11230, ZN => n15518);
   U3217 : AOI22_X1 port map( A1 => n9840, A2 => n11127, B1 => n10032, B2 => 
                           n11231, ZN => n15517);
   U3218 : AOI22_X1 port map( A1 => n9808, A2 => n16077, B1 => n9872, B2 => 
                           n11131, ZN => n15516);
   U3219 : NAND4_X1 port map( A1 => n15519, A2 => n15518, A3 => n15517, A4 => 
                           n15516, ZN => n15525);
   U3220 : AOI22_X1 port map( A1 => n9712, A2 => n16048, B1 => n9552, B2 => 
                           n11225, ZN => n15523);
   U3221 : AOI22_X1 port map( A1 => n9616, A2 => n11131, B1 => n9648, B2 => 
                           n11128, ZN => n15522);
   U3222 : AOI22_X1 port map( A1 => n9776, A2 => n16072, B1 => n9680, B2 => 
                           n11135, ZN => n15521);
   U3223 : AOI22_X1 port map( A1 => n9744, A2 => n16053, B1 => n9584, B2 => 
                           n11145, ZN => n15520);
   U3224 : NAND4_X1 port map( A1 => n15523, A2 => n15522, A3 => n15521, A4 => 
                           n15520, ZN => n15524);
   U3225 : AOI22_X1 port map( A1 => n15880, A2 => n15525, B1 => n15613, B2 => 
                           n15524, ZN => n15526);
   U3226 : OAI21_X1 port map( B1 => n15905, B2 => n15527, A => n15526, ZN => 
                           OUT1(25));
   U3227 : AOI22_X1 port map( A1 => n9199, A2 => n11153, B1 => n9455, B2 => 
                           n11151, ZN => n15531);
   U3228 : AOI22_X1 port map( A1 => n9103, A2 => n11142, B1 => n9487, B2 => 
                           n11133, ZN => n15530);
   U3229 : AOI22_X1 port map( A1 => n9039, A2 => n11150, B1 => n9327, B2 => 
                           n11138, ZN => n15529);
   U3230 : AOI22_X1 port map( A1 => n9295, A2 => n11152, B1 => n9071, B2 => 
                           n10043, ZN => n15528);
   U3231 : NAND4_X1 port map( A1 => n15531, A2 => n15530, A3 => n15529, A4 => 
                           n15528, ZN => n15537);
   U3232 : AOI22_X1 port map( A1 => n9359, A2 => n11139, B1 => n9167, B2 => 
                           n11140, ZN => n15535);
   U3233 : AOI22_X1 port map( A1 => n9135, A2 => n11137, B1 => n9231, B2 => 
                           n11143, ZN => n15534);
   U3234 : AOI22_X1 port map( A1 => n9391, A2 => n10053, B1 => n9519, B2 => 
                           n10052, ZN => n15533);
   U3235 : AOI22_X1 port map( A1 => n9263, A2 => n11132, B1 => n9423, B2 => 
                           n11141, ZN => n15532);
   U3236 : NAND4_X1 port map( A1 => n15535, A2 => n15534, A3 => n15533, A4 => 
                           n15532, ZN => n15536);
   U3237 : NOR2_X1 port map( A1 => n15537, A2 => n15536, ZN => n15549);
   U3238 : AOI22_X1 port map( A1 => n10031, A2 => n11146, B1 => n9935, B2 => 
                           n11232, ZN => n15541);
   U3239 : AOI22_X1 port map( A1 => n9999, A2 => n16053, B1 => n9903, B2 => 
                           n11144, ZN => n15540);
   U3240 : AOI22_X1 port map( A1 => n9871, A2 => n11131, B1 => n9839, B2 => 
                           n11127, ZN => n15539);
   U3241 : AOI22_X1 port map( A1 => n9967, A2 => n11129, B1 => n9807, B2 => 
                           n11225, ZN => n15538);
   U3242 : NAND4_X1 port map( A1 => n15541, A2 => n15540, A3 => n15539, A4 => 
                           n15538, ZN => n15547);
   U3243 : AOI22_X1 port map( A1 => n9583, A2 => n11127, B1 => n9679, B2 => 
                           n16079, ZN => n15545);
   U3244 : AOI22_X1 port map( A1 => n9647, A2 => n11144, B1 => n9743, B2 => 
                           n11130, ZN => n15544);
   U3245 : AOI22_X1 port map( A1 => n9551, A2 => n11134, B1 => n9775, B2 => 
                           n11231, ZN => n15543);
   U3246 : AOI22_X1 port map( A1 => n9711, A2 => n11230, B1 => n9615, B2 => 
                           n11131, ZN => n15542);
   U3247 : NAND4_X1 port map( A1 => n15545, A2 => n15544, A3 => n15543, A4 => 
                           n15542, ZN => n15546);
   U3248 : AOI22_X1 port map( A1 => n15880, A2 => n15547, B1 => n15613, B2 => 
                           n15546, ZN => n15548);
   U3249 : OAI21_X1 port map( B1 => n15905, B2 => n15549, A => n15548, ZN => 
                           OUT1(24));
   U3250 : AOI22_X1 port map( A1 => n9390, A2 => n11154, B1 => n9070, B2 => 
                           n11149, ZN => n15553);
   U3251 : AOI22_X1 port map( A1 => n9038, A2 => n11150, B1 => n9102, B2 => 
                           n11142, ZN => n15552);
   U3252 : AOI22_X1 port map( A1 => n9422, A2 => n11141, B1 => n9230, B2 => 
                           n11143, ZN => n15551);
   U3253 : AOI22_X1 port map( A1 => n9134, A2 => n11137, B1 => n9166, B2 => 
                           n11140, ZN => n15550);
   U3254 : NAND4_X1 port map( A1 => n15553, A2 => n15552, A3 => n15551, A4 => 
                           n15550, ZN => n15559);
   U3255 : AOI22_X1 port map( A1 => n9486, A2 => n11133, B1 => n9326, B2 => 
                           n11138, ZN => n15557);
   U3256 : AOI22_X1 port map( A1 => n9262, A2 => n11132, B1 => n9518, B2 => 
                           n10052, ZN => n15556);
   U3257 : AOI22_X1 port map( A1 => n9294, A2 => n11152, B1 => n9454, B2 => 
                           n10047, ZN => n15555);
   U3258 : AOI22_X1 port map( A1 => n9198, A2 => n11153, B1 => n9358, B2 => 
                           n11139, ZN => n15554);
   U3259 : NAND4_X1 port map( A1 => n15557, A2 => n15556, A3 => n15555, A4 => 
                           n15554, ZN => n15558);
   U3260 : NOR2_X1 port map( A1 => n15559, A2 => n15558, ZN => n15571);
   U3261 : AOI22_X1 port map( A1 => n9838, A2 => n11127, B1 => n9998, B2 => 
                           n16053, ZN => n15563);
   U3262 : AOI22_X1 port map( A1 => n10030, A2 => n16072, B1 => n9966, B2 => 
                           n16048, ZN => n15562);
   U3263 : AOI22_X1 port map( A1 => n9806, A2 => n16077, B1 => n9870, B2 => 
                           n16078, ZN => n15561);
   U3264 : AOI22_X1 port map( A1 => n9934, A2 => n11232, B1 => n9902, B2 => 
                           n11144, ZN => n15560);
   U3265 : NAND4_X1 port map( A1 => n15563, A2 => n15562, A3 => n15561, A4 => 
                           n15560, ZN => n15569);
   U3266 : AOI22_X1 port map( A1 => n9646, A2 => n11128, B1 => n9582, B2 => 
                           n11145, ZN => n15567);
   U3267 : AOI22_X1 port map( A1 => n9678, A2 => n16079, B1 => n9742, B2 => 
                           n16053, ZN => n15566);
   U3268 : AOI22_X1 port map( A1 => n9774, A2 => n16072, B1 => n9710, B2 => 
                           n11230, ZN => n15565);
   U3269 : AOI22_X1 port map( A1 => n9614, A2 => n11229, B1 => n9550, B2 => 
                           n11134, ZN => n15564);
   U3270 : NAND4_X1 port map( A1 => n15567, A2 => n15566, A3 => n15565, A4 => 
                           n15564, ZN => n15568);
   U3271 : AOI22_X1 port map( A1 => n15880, A2 => n15569, B1 => n15613, B2 => 
                           n15568, ZN => n15570);
   U3272 : OAI21_X1 port map( B1 => n16090, B2 => n15571, A => n15570, ZN => 
                           OUT1(23));
   U3273 : AOI22_X1 port map( A1 => n9453, A2 => n10047, B1 => n9165, B2 => 
                           n11140, ZN => n15575);
   U3274 : AOI22_X1 port map( A1 => n9229, A2 => n10039, B1 => n9517, B2 => 
                           n10052, ZN => n15574);
   U3275 : AOI22_X1 port map( A1 => n9037, A2 => n11150, B1 => n9389, B2 => 
                           n11154, ZN => n15573);
   U3276 : AOI22_X1 port map( A1 => n9325, A2 => n11138, B1 => n9293, B2 => 
                           n11152, ZN => n15572);
   U3277 : NAND4_X1 port map( A1 => n15575, A2 => n15574, A3 => n15573, A4 => 
                           n15572, ZN => n15581);
   U3278 : AOI22_X1 port map( A1 => n9197, A2 => n11153, B1 => n9101, B2 => 
                           n11142, ZN => n15579);
   U3279 : AOI22_X1 port map( A1 => n9357, A2 => n11139, B1 => n9069, B2 => 
                           n11149, ZN => n15578);
   U3280 : AOI22_X1 port map( A1 => n9261, A2 => n10054, B1 => n9133, B2 => 
                           n11137, ZN => n15577);
   U3281 : AOI22_X1 port map( A1 => n9485, A2 => n11133, B1 => n9421, B2 => 
                           n11141, ZN => n15576);
   U3282 : NAND4_X1 port map( A1 => n15579, A2 => n15578, A3 => n15577, A4 => 
                           n15576, ZN => n15580);
   U3283 : NOR2_X1 port map( A1 => n15581, A2 => n15580, ZN => n15593);
   U3284 : AOI22_X1 port map( A1 => n9933, A2 => n11232, B1 => n9965, B2 => 
                           n16048, ZN => n15585);
   U3285 : AOI22_X1 port map( A1 => n9901, A2 => n11148, B1 => n9997, B2 => 
                           n11130, ZN => n15584);
   U3286 : AOI22_X1 port map( A1 => n9837, A2 => n11127, B1 => n9869, B2 => 
                           n11131, ZN => n15583);
   U3287 : AOI22_X1 port map( A1 => n9805, A2 => n11134, B1 => n10029, B2 => 
                           n11146, ZN => n15582);
   U3288 : NAND4_X1 port map( A1 => n15585, A2 => n15584, A3 => n15583, A4 => 
                           n15582, ZN => n15591);
   U3289 : AOI22_X1 port map( A1 => n9741, A2 => n16053, B1 => n9645, B2 => 
                           n11128, ZN => n15589);
   U3290 : AOI22_X1 port map( A1 => n9709, A2 => n16048, B1 => n9549, B2 => 
                           n11225, ZN => n15588);
   U3291 : AOI22_X1 port map( A1 => n9581, A2 => n11127, B1 => n9613, B2 => 
                           n11229, ZN => n15587);
   U3292 : AOI22_X1 port map( A1 => n9773, A2 => n16072, B1 => n9677, B2 => 
                           n11232, ZN => n15586);
   U3293 : NAND4_X1 port map( A1 => n15589, A2 => n15588, A3 => n15587, A4 => 
                           n15586, ZN => n15590);
   U3294 : AOI22_X1 port map( A1 => n15880, A2 => n15591, B1 => n15613, B2 => 
                           n15590, ZN => n15592);
   U3295 : OAI21_X1 port map( B1 => n16090, B2 => n15593, A => n15592, ZN => 
                           OUT1(22));
   U3296 : AOI22_X1 port map( A1 => n9036, A2 => n10045, B1 => n9100, B2 => 
                           n10040, ZN => n15597);
   U3297 : AOI22_X1 port map( A1 => n9324, A2 => n11138, B1 => n9132, B2 => 
                           n11137, ZN => n15596);
   U3298 : AOI22_X1 port map( A1 => n9356, A2 => n11139, B1 => n9260, B2 => 
                           n11132, ZN => n15595);
   U3299 : AOI22_X1 port map( A1 => n9292, A2 => n10049, B1 => n9228, B2 => 
                           n11143, ZN => n15594);
   U3300 : NAND4_X1 port map( A1 => n15597, A2 => n15596, A3 => n15595, A4 => 
                           n15594, ZN => n15603);
   U3301 : AOI22_X1 port map( A1 => n9164, A2 => n10041, B1 => n9484, B2 => 
                           n11133, ZN => n15601);
   U3302 : AOI22_X1 port map( A1 => n9196, A2 => n11153, B1 => n9420, B2 => 
                           n11141, ZN => n15600);
   U3303 : AOI22_X1 port map( A1 => n9452, A2 => n11151, B1 => n9388, B2 => 
                           n11154, ZN => n15599);
   U3304 : AOI22_X1 port map( A1 => n9516, A2 => n11136, B1 => n9068, B2 => 
                           n11149, ZN => n15598);
   U3305 : NAND4_X1 port map( A1 => n15601, A2 => n15600, A3 => n15599, A4 => 
                           n15598, ZN => n15602);
   U3306 : NOR2_X1 port map( A1 => n15603, A2 => n15602, ZN => n15616);
   U3307 : AOI22_X1 port map( A1 => n10028, A2 => n11231, B1 => n9868, B2 => 
                           n11131, ZN => n15607);
   U3308 : AOI22_X1 port map( A1 => n9804, A2 => n16077, B1 => n9996, B2 => 
                           n11228, ZN => n15606);
   U3309 : AOI22_X1 port map( A1 => n9964, A2 => n11230, B1 => n9932, B2 => 
                           n16079, ZN => n15605);
   U3310 : AOI22_X1 port map( A1 => n9836, A2 => n11145, B1 => n9900, B2 => 
                           n11128, ZN => n15604);
   U3311 : NAND4_X1 port map( A1 => n15607, A2 => n15606, A3 => n15605, A4 => 
                           n15604, ZN => n15614);
   U3312 : AOI22_X1 port map( A1 => n9676, A2 => n16079, B1 => n9612, B2 => 
                           n11131, ZN => n15611);
   U3313 : AOI22_X1 port map( A1 => n9708, A2 => n16048, B1 => n9772, B2 => 
                           n16072, ZN => n15610);
   U3314 : AOI22_X1 port map( A1 => n9580, A2 => n11127, B1 => n9644, B2 => 
                           n11128, ZN => n15609);
   U3315 : AOI22_X1 port map( A1 => n9740, A2 => n11228, B1 => n9548, B2 => 
                           n16077, ZN => n15608);
   U3316 : NAND4_X1 port map( A1 => n15611, A2 => n15610, A3 => n15609, A4 => 
                           n15608, ZN => n15612);
   U3317 : AOI22_X1 port map( A1 => n15880, A2 => n15614, B1 => n15613, B2 => 
                           n15612, ZN => n15615);
   U3318 : OAI21_X1 port map( B1 => n16090, B2 => n15616, A => n15615, ZN => 
                           OUT1(21));
   U3319 : AOI22_X1 port map( A1 => n9451, A2 => n10047, B1 => n9323, B2 => 
                           n11138, ZN => n15620);
   U3320 : AOI22_X1 port map( A1 => n9355, A2 => n11139, B1 => n9227, B2 => 
                           n11143, ZN => n15619);
   U3321 : AOI22_X1 port map( A1 => n9099, A2 => n11142, B1 => n9419, B2 => 
                           n11141, ZN => n15618);
   U3322 : AOI22_X1 port map( A1 => n9131, A2 => n11137, B1 => n9483, B2 => 
                           n11133, ZN => n15617);
   U3323 : NAND4_X1 port map( A1 => n15620, A2 => n15619, A3 => n15618, A4 => 
                           n15617, ZN => n15626);
   U3324 : AOI22_X1 port map( A1 => n9195, A2 => n11153, B1 => n9035, B2 => 
                           n11150, ZN => n15624);
   U3325 : AOI22_X1 port map( A1 => n9515, A2 => n11136, B1 => n9067, B2 => 
                           n11149, ZN => n15623);
   U3326 : AOI22_X1 port map( A1 => n9259, A2 => n11132, B1 => n9387, B2 => 
                           n10053, ZN => n15622);
   U3327 : AOI22_X1 port map( A1 => n9291, A2 => n11152, B1 => n9163, B2 => 
                           n11140, ZN => n15621);
   U3328 : NAND4_X1 port map( A1 => n15624, A2 => n15623, A3 => n15622, A4 => 
                           n15621, ZN => n15625);
   U3329 : NOR2_X1 port map( A1 => n15626, A2 => n15625, ZN => n15638);
   U3330 : AOI22_X1 port map( A1 => n9899, A2 => n11128, B1 => n9867, B2 => 
                           n11131, ZN => n15630);
   U3331 : AOI22_X1 port map( A1 => n9963, A2 => n11230, B1 => n9835, B2 => 
                           n11127, ZN => n15629);
   U3332 : AOI22_X1 port map( A1 => n10027, A2 => n11231, B1 => n9931, B2 => 
                           n11232, ZN => n15628);
   U3333 : AOI22_X1 port map( A1 => n9803, A2 => n11225, B1 => n9995, B2 => 
                           n11130, ZN => n15627);
   U3334 : NAND4_X1 port map( A1 => n15630, A2 => n15629, A3 => n15628, A4 => 
                           n15627, ZN => n15636);
   U3335 : AOI22_X1 port map( A1 => n9675, A2 => n11232, B1 => n9771, B2 => 
                           n11231, ZN => n15634);
   U3336 : AOI22_X1 port map( A1 => n9547, A2 => n11225, B1 => n9707, B2 => 
                           n11230, ZN => n15633);
   U3337 : AOI22_X1 port map( A1 => n9611, A2 => n11131, B1 => n9643, B2 => 
                           n11128, ZN => n15632);
   U3338 : AOI22_X1 port map( A1 => n9739, A2 => n11228, B1 => n9579, B2 => 
                           n11127, ZN => n15631);
   U3339 : NAND4_X1 port map( A1 => n15634, A2 => n15633, A3 => n15632, A4 => 
                           n15631, ZN => n15635);
   U3340 : AOI22_X1 port map( A1 => n15880, A2 => n15636, B1 => n16085, B2 => 
                           n15635, ZN => n15637);
   U3341 : OAI21_X1 port map( B1 => n16090, B2 => n15638, A => n15637, ZN => 
                           OUT1(20));
   U3342 : AOI22_X1 port map( A1 => n9130, A2 => n11137, B1 => n9258, B2 => 
                           n11132, ZN => n15642);
   U3343 : AOI22_X1 port map( A1 => n9066, A2 => n11149, B1 => n9322, B2 => 
                           n10044, ZN => n15641);
   U3344 : AOI22_X1 port map( A1 => n9450, A2 => n11151, B1 => n9034, B2 => 
                           n11150, ZN => n15640);
   U3345 : AOI22_X1 port map( A1 => n9354, A2 => n11139, B1 => n9162, B2 => 
                           n11140, ZN => n15639);
   U3346 : NAND4_X1 port map( A1 => n15642, A2 => n15641, A3 => n15640, A4 => 
                           n15639, ZN => n15648);
   U3347 : AOI22_X1 port map( A1 => n9386, A2 => n11154, B1 => n9290, B2 => 
                           n11152, ZN => n15646);
   U3348 : AOI22_X1 port map( A1 => n9226, A2 => n11143, B1 => n9418, B2 => 
                           n10048, ZN => n15645);
   U3349 : AOI22_X1 port map( A1 => n9482, A2 => n10042, B1 => n9514, B2 => 
                           n11136, ZN => n15644);
   U3350 : AOI22_X1 port map( A1 => n9194, A2 => n11153, B1 => n9098, B2 => 
                           n11142, ZN => n15643);
   U3351 : NAND4_X1 port map( A1 => n15646, A2 => n15645, A3 => n15644, A4 => 
                           n15643, ZN => n15647);
   U3352 : NOR2_X1 port map( A1 => n15648, A2 => n15647, ZN => n15660);
   U3353 : AOI22_X1 port map( A1 => n9962, A2 => n11129, B1 => n9994, B2 => 
                           n11228, ZN => n15652);
   U3354 : AOI22_X1 port map( A1 => n9866, A2 => n11229, B1 => n10026, B2 => 
                           n11146, ZN => n15651);
   U3355 : AOI22_X1 port map( A1 => n9802, A2 => n11225, B1 => n9834, B2 => 
                           n11127, ZN => n15650);
   U3356 : AOI22_X1 port map( A1 => n9930, A2 => n16079, B1 => n9898, B2 => 
                           n11128, ZN => n15649);
   U3357 : NAND4_X1 port map( A1 => n15652, A2 => n15651, A3 => n15650, A4 => 
                           n15649, ZN => n15658);
   U3358 : AOI22_X1 port map( A1 => n9642, A2 => n11148, B1 => n9546, B2 => 
                           n11134, ZN => n15656);
   U3359 : AOI22_X1 port map( A1 => n9738, A2 => n11228, B1 => n9706, B2 => 
                           n11230, ZN => n15655);
   U3360 : AOI22_X1 port map( A1 => n9578, A2 => n11127, B1 => n9770, B2 => 
                           n16072, ZN => n15654);
   U3361 : AOI22_X1 port map( A1 => n9610, A2 => n11131, B1 => n9674, B2 => 
                           n11232, ZN => n15653);
   U3362 : NAND4_X1 port map( A1 => n15656, A2 => n15655, A3 => n15654, A4 => 
                           n15653, ZN => n15657);
   U3363 : AOI22_X1 port map( A1 => n15880, A2 => n15658, B1 => n16085, B2 => 
                           n15657, ZN => n15659);
   U3364 : OAI21_X1 port map( B1 => n16090, B2 => n15660, A => n15659, ZN => 
                           OUT1(19));
   U3365 : AOI22_X1 port map( A1 => n9193, A2 => n10051, B1 => n9289, B2 => 
                           n10049, ZN => n15664);
   U3366 : AOI22_X1 port map( A1 => n9353, A2 => n10050, B1 => n9321, B2 => 
                           n11138, ZN => n15663);
   U3367 : AOI22_X1 port map( A1 => n9513, A2 => n11136, B1 => n9097, B2 => 
                           n11142, ZN => n15662);
   U3368 : AOI22_X1 port map( A1 => n9161, A2 => n10041, B1 => n9257, B2 => 
                           n11132, ZN => n15661);
   U3369 : NAND4_X1 port map( A1 => n15664, A2 => n15663, A3 => n15662, A4 => 
                           n15661, ZN => n15670);
   U3370 : AOI22_X1 port map( A1 => n9065, A2 => n11149, B1 => n9225, B2 => 
                           n11143, ZN => n15668);
   U3371 : AOI22_X1 port map( A1 => n9033, A2 => n10045, B1 => n9417, B2 => 
                           n11141, ZN => n15667);
   U3372 : AOI22_X1 port map( A1 => n9481, A2 => n10042, B1 => n9385, B2 => 
                           n11154, ZN => n15666);
   U3373 : AOI22_X1 port map( A1 => n9129, A2 => n11137, B1 => n9449, B2 => 
                           n10047, ZN => n15665);
   U3374 : NAND4_X1 port map( A1 => n15668, A2 => n15667, A3 => n15666, A4 => 
                           n15665, ZN => n15669);
   U3375 : NOR2_X1 port map( A1 => n15670, A2 => n15669, ZN => n15682);
   U3376 : CLKBUF_X1 port map( A => n15835, Z => n16087);
   U3377 : AOI22_X1 port map( A1 => n9897, A2 => n11128, B1 => n9961, B2 => 
                           n11230, ZN => n15674);
   U3378 : AOI22_X1 port map( A1 => n9833, A2 => n11145, B1 => n9865, B2 => 
                           n16078, ZN => n15673);
   U3379 : AOI22_X1 port map( A1 => n10025, A2 => n11231, B1 => n9993, B2 => 
                           n16053, ZN => n15672);
   U3380 : AOI22_X1 port map( A1 => n9801, A2 => n11134, B1 => n9929, B2 => 
                           n16079, ZN => n15671);
   U3381 : NAND4_X1 port map( A1 => n15674, A2 => n15673, A3 => n15672, A4 => 
                           n15671, ZN => n15680);
   U3382 : AOI22_X1 port map( A1 => n9705, A2 => n16048, B1 => n9577, B2 => 
                           n11145, ZN => n15678);
   U3383 : AOI22_X1 port map( A1 => n9545, A2 => n16077, B1 => n9673, B2 => 
                           n11232, ZN => n15677);
   U3384 : AOI22_X1 port map( A1 => n9609, A2 => n11229, B1 => n9641, B2 => 
                           n11128, ZN => n15676);
   U3385 : AOI22_X1 port map( A1 => n9769, A2 => n11231, B1 => n9737, B2 => 
                           n11130, ZN => n15675);
   U3386 : NAND4_X1 port map( A1 => n15678, A2 => n15677, A3 => n15676, A4 => 
                           n15675, ZN => n15679);
   U3387 : AOI22_X1 port map( A1 => n16087, A2 => n15680, B1 => n16085, B2 => 
                           n15679, ZN => n15681);
   U3388 : OAI21_X1 port map( B1 => n16090, B2 => n15682, A => n15681, ZN => 
                           OUT1(18));
   U3389 : AOI22_X1 port map( A1 => n9288, A2 => n10049, B1 => n9512, B2 => 
                           n11136, ZN => n15686);
   U3390 : AOI22_X1 port map( A1 => n9416, A2 => n10048, B1 => n9192, B2 => 
                           n11153, ZN => n15685);
   U3391 : AOI22_X1 port map( A1 => n9256, A2 => n11132, B1 => n9096, B2 => 
                           n10040, ZN => n15684);
   U3392 : AOI22_X1 port map( A1 => n9352, A2 => n11139, B1 => n9160, B2 => 
                           n11140, ZN => n15683);
   U3393 : NAND4_X1 port map( A1 => n15686, A2 => n15685, A3 => n15684, A4 => 
                           n15683, ZN => n15692);
   U3394 : AOI22_X1 port map( A1 => n9480, A2 => n11133, B1 => n9320, B2 => 
                           n11138, ZN => n15690);
   U3395 : AOI22_X1 port map( A1 => n9448, A2 => n10047, B1 => n9384, B2 => 
                           n11154, ZN => n15689);
   U3396 : AOI22_X1 port map( A1 => n9064, A2 => n11149, B1 => n9032, B2 => 
                           n10045, ZN => n15688);
   U3397 : AOI22_X1 port map( A1 => n9224, A2 => n10039, B1 => n9128, B2 => 
                           n10046, ZN => n15687);
   U3398 : NAND4_X1 port map( A1 => n15690, A2 => n15689, A3 => n15688, A4 => 
                           n15687, ZN => n15691);
   U3399 : NOR2_X1 port map( A1 => n15692, A2 => n15691, ZN => n15704);
   U3400 : AOI22_X1 port map( A1 => n9960, A2 => n11230, B1 => n9832, B2 => 
                           n11145, ZN => n15696);
   U3401 : AOI22_X1 port map( A1 => n9928, A2 => n11232, B1 => n9800, B2 => 
                           n16077, ZN => n15695);
   U3402 : AOI22_X1 port map( A1 => n9896, A2 => n11144, B1 => n10024, B2 => 
                           n11146, ZN => n15694);
   U3403 : AOI22_X1 port map( A1 => n9992, A2 => n16053, B1 => n9864, B2 => 
                           n11131, ZN => n15693);
   U3404 : NAND4_X1 port map( A1 => n15696, A2 => n15695, A3 => n15694, A4 => 
                           n15693, ZN => n15702);
   U3405 : AOI22_X1 port map( A1 => n9672, A2 => n11135, B1 => n9640, B2 => 
                           n11148, ZN => n15700);
   U3406 : AOI22_X1 port map( A1 => n9608, A2 => n16078, B1 => n9768, B2 => 
                           n11231, ZN => n15699);
   U3407 : AOI22_X1 port map( A1 => n9736, A2 => n16053, B1 => n9704, B2 => 
                           n16048, ZN => n15698);
   U3408 : AOI22_X1 port map( A1 => n9544, A2 => n11134, B1 => n9576, B2 => 
                           n11127, ZN => n15697);
   U3409 : NAND4_X1 port map( A1 => n15700, A2 => n15699, A3 => n15698, A4 => 
                           n15697, ZN => n15701);
   U3410 : AOI22_X1 port map( A1 => n16087, A2 => n15702, B1 => n16085, B2 => 
                           n15701, ZN => n15703);
   U3411 : OAI21_X1 port map( B1 => n16090, B2 => n15704, A => n15703, ZN => 
                           OUT1(17));
   U3412 : AOI22_X1 port map( A1 => n9159, A2 => n11140, B1 => n9031, B2 => 
                           n10045, ZN => n15708);
   U3413 : AOI22_X1 port map( A1 => n9319, A2 => n11138, B1 => n9383, B2 => 
                           n10053, ZN => n15707);
   U3414 : AOI22_X1 port map( A1 => n9511, A2 => n10052, B1 => n9095, B2 => 
                           n10040, ZN => n15706);
   U3415 : AOI22_X1 port map( A1 => n9255, A2 => n11132, B1 => n9191, B2 => 
                           n11153, ZN => n15705);
   U3416 : NAND4_X1 port map( A1 => n15708, A2 => n15707, A3 => n15706, A4 => 
                           n15705, ZN => n15714);
   U3417 : AOI22_X1 port map( A1 => n9223, A2 => n11143, B1 => n9351, B2 => 
                           n10050, ZN => n15712);
   U3418 : AOI22_X1 port map( A1 => n9415, A2 => n11141, B1 => n9063, B2 => 
                           n11149, ZN => n15711);
   U3419 : AOI22_X1 port map( A1 => n9447, A2 => n11151, B1 => n9479, B2 => 
                           n11133, ZN => n15710);
   U3420 : AOI22_X1 port map( A1 => n9287, A2 => n11152, B1 => n9127, B2 => 
                           n10046, ZN => n15709);
   U3421 : NAND4_X1 port map( A1 => n15712, A2 => n15711, A3 => n15710, A4 => 
                           n15709, ZN => n15713);
   U3422 : NOR2_X1 port map( A1 => n15714, A2 => n15713, ZN => n15726);
   U3423 : AOI22_X1 port map( A1 => n10023, A2 => n16072, B1 => n9895, B2 => 
                           n11128, ZN => n15718);
   U3424 : AOI22_X1 port map( A1 => n9831, A2 => n11127, B1 => n9799, B2 => 
                           n11225, ZN => n15717);
   U3425 : AOI22_X1 port map( A1 => n9927, A2 => n16079, B1 => n9991, B2 => 
                           n11228, ZN => n15716);
   U3426 : AOI22_X1 port map( A1 => n9863, A2 => n16078, B1 => n9959, B2 => 
                           n16048, ZN => n15715);
   U3427 : NAND4_X1 port map( A1 => n15718, A2 => n15717, A3 => n15716, A4 => 
                           n15715, ZN => n15724);
   U3428 : AOI22_X1 port map( A1 => n9767, A2 => n11146, B1 => n9543, B2 => 
                           n11225, ZN => n15722);
   U3429 : AOI22_X1 port map( A1 => n9703, A2 => n11129, B1 => n9639, B2 => 
                           n11128, ZN => n15721);
   U3430 : AOI22_X1 port map( A1 => n9575, A2 => n11145, B1 => n9735, B2 => 
                           n16053, ZN => n15720);
   U3431 : AOI22_X1 port map( A1 => n9671, A2 => n11232, B1 => n9607, B2 => 
                           n11229, ZN => n15719);
   U3432 : NAND4_X1 port map( A1 => n15722, A2 => n15721, A3 => n15720, A4 => 
                           n15719, ZN => n15723);
   U3433 : AOI22_X1 port map( A1 => n15880, A2 => n15724, B1 => n16085, B2 => 
                           n15723, ZN => n15725);
   U3434 : OAI21_X1 port map( B1 => n16090, B2 => n15726, A => n15725, ZN => 
                           OUT1(16));
   U3435 : AOI22_X1 port map( A1 => n9414, A2 => n10048, B1 => n9382, B2 => 
                           n10053, ZN => n15730);
   U3436 : AOI22_X1 port map( A1 => n9254, A2 => n11132, B1 => n9030, B2 => 
                           n10045, ZN => n15729);
   U3437 : AOI22_X1 port map( A1 => n9446, A2 => n10047, B1 => n9062, B2 => 
                           n10043, ZN => n15728);
   U3438 : AOI22_X1 port map( A1 => n9190, A2 => n11153, B1 => n9318, B2 => 
                           n10044, ZN => n15727);
   U3439 : NAND4_X1 port map( A1 => n15730, A2 => n15729, A3 => n15728, A4 => 
                           n15727, ZN => n15736);
   U3440 : AOI22_X1 port map( A1 => n9350, A2 => n11139, B1 => n9126, B2 => 
                           n10046, ZN => n15734);
   U3441 : AOI22_X1 port map( A1 => n9222, A2 => n11143, B1 => n9286, B2 => 
                           n11152, ZN => n15733);
   U3442 : AOI22_X1 port map( A1 => n9478, A2 => n11133, B1 => n9158, B2 => 
                           n11140, ZN => n15732);
   U3443 : AOI22_X1 port map( A1 => n9510, A2 => n11136, B1 => n9094, B2 => 
                           n11142, ZN => n15731);
   U3444 : NAND4_X1 port map( A1 => n15734, A2 => n15733, A3 => n15732, A4 => 
                           n15731, ZN => n15735);
   U3445 : NOR2_X1 port map( A1 => n15736, A2 => n15735, ZN => n15748);
   U3446 : AOI22_X1 port map( A1 => n9894, A2 => n11148, B1 => n9862, B2 => 
                           n11131, ZN => n15740);
   U3447 : AOI22_X1 port map( A1 => n9798, A2 => n11134, B1 => n9830, B2 => 
                           n11127, ZN => n15739);
   U3448 : AOI22_X1 port map( A1 => n10022, A2 => n11146, B1 => n9990, B2 => 
                           n11130, ZN => n15738);
   U3449 : AOI22_X1 port map( A1 => n9926, A2 => n11135, B1 => n9958, B2 => 
                           n11129, ZN => n15737);
   U3450 : NAND4_X1 port map( A1 => n15740, A2 => n15739, A3 => n15738, A4 => 
                           n15737, ZN => n15746);
   U3451 : AOI22_X1 port map( A1 => n9606, A2 => n11229, B1 => n9542, B2 => 
                           n11225, ZN => n15744);
   U3452 : AOI22_X1 port map( A1 => n9574, A2 => n11127, B1 => n9766, B2 => 
                           n11231, ZN => n15743);
   U3453 : AOI22_X1 port map( A1 => n9734, A2 => n11228, B1 => n9702, B2 => 
                           n16048, ZN => n15742);
   U3454 : AOI22_X1 port map( A1 => n9670, A2 => n16079, B1 => n9638, B2 => 
                           n11144, ZN => n15741);
   U3455 : NAND4_X1 port map( A1 => n15744, A2 => n15743, A3 => n15742, A4 => 
                           n15741, ZN => n15745);
   U3456 : AOI22_X1 port map( A1 => n15880, A2 => n15746, B1 => n16085, B2 => 
                           n15745, ZN => n15747);
   U3457 : OAI21_X1 port map( B1 => n16090, B2 => n15748, A => n15747, ZN => 
                           OUT1(15));
   U3458 : AOI22_X1 port map( A1 => n9029, A2 => n10045, B1 => n9381, B2 => 
                           n11154, ZN => n15752);
   U3459 : AOI22_X1 port map( A1 => n9253, A2 => n10054, B1 => n9413, B2 => 
                           n10048, ZN => n15751);
   U3460 : AOI22_X1 port map( A1 => n9445, A2 => n11151, B1 => n9285, B2 => 
                           n11152, ZN => n15750);
   U3461 : AOI22_X1 port map( A1 => n9509, A2 => n11136, B1 => n9477, B2 => 
                           n11133, ZN => n15749);
   U3462 : NAND4_X1 port map( A1 => n15752, A2 => n15751, A3 => n15750, A4 => 
                           n15749, ZN => n15758);
   U3463 : AOI22_X1 port map( A1 => n9317, A2 => n10044, B1 => n9061, B2 => 
                           n11149, ZN => n15756);
   U3464 : AOI22_X1 port map( A1 => n9093, A2 => n10040, B1 => n9189, B2 => 
                           n11153, ZN => n15755);
   U3465 : AOI22_X1 port map( A1 => n9125, A2 => n10046, B1 => n9221, B2 => 
                           n11143, ZN => n15754);
   U3466 : AOI22_X1 port map( A1 => n9349, A2 => n11139, B1 => n9157, B2 => 
                           n11140, ZN => n15753);
   U3467 : NAND4_X1 port map( A1 => n15756, A2 => n15755, A3 => n15754, A4 => 
                           n15753, ZN => n15757);
   U3468 : NOR2_X1 port map( A1 => n15758, A2 => n15757, ZN => n15770);
   U3469 : AOI22_X1 port map( A1 => n9925, A2 => n11232, B1 => n9989, B2 => 
                           n11228, ZN => n15762);
   U3470 : AOI22_X1 port map( A1 => n9957, A2 => n11129, B1 => n9797, B2 => 
                           n11134, ZN => n15761);
   U3471 : AOI22_X1 port map( A1 => n10021, A2 => n11146, B1 => n9861, B2 => 
                           n11229, ZN => n15760);
   U3472 : AOI22_X1 port map( A1 => n9829, A2 => n11145, B1 => n9893, B2 => 
                           n11144, ZN => n15759);
   U3473 : NAND4_X1 port map( A1 => n15762, A2 => n15761, A3 => n15760, A4 => 
                           n15759, ZN => n15768);
   U3474 : AOI22_X1 port map( A1 => n9733, A2 => n11228, B1 => n9573, B2 => 
                           n11145, ZN => n15766);
   U3475 : AOI22_X1 port map( A1 => n9669, A2 => n11135, B1 => n9637, B2 => 
                           n11144, ZN => n15765);
   U3476 : AOI22_X1 port map( A1 => n9765, A2 => n11146, B1 => n9605, B2 => 
                           n11229, ZN => n15764);
   U3477 : AOI22_X1 port map( A1 => n9541, A2 => n11134, B1 => n9701, B2 => 
                           n11129, ZN => n15763);
   U3478 : NAND4_X1 port map( A1 => n15766, A2 => n15765, A3 => n15764, A4 => 
                           n15763, ZN => n15767);
   U3479 : AOI22_X1 port map( A1 => n15880, A2 => n15768, B1 => n16085, B2 => 
                           n15767, ZN => n15769);
   U3480 : OAI21_X1 port map( B1 => n16090, B2 => n15770, A => n15769, ZN => 
                           OUT1(14));
   U3481 : AOI22_X1 port map( A1 => n9092, A2 => n10040, B1 => n9220, B2 => 
                           n10039, ZN => n15774);
   U3482 : AOI22_X1 port map( A1 => n9380, A2 => n11154, B1 => n9124, B2 => 
                           n10046, ZN => n15773);
   U3483 : AOI22_X1 port map( A1 => n9476, A2 => n11133, B1 => n9028, B2 => 
                           n10045, ZN => n15772);
   U3484 : AOI22_X1 port map( A1 => n9156, A2 => n11140, B1 => n9060, B2 => 
                           n11149, ZN => n15771);
   U3485 : NAND4_X1 port map( A1 => n15774, A2 => n15773, A3 => n15772, A4 => 
                           n15771, ZN => n15780);
   U3486 : AOI22_X1 port map( A1 => n9412, A2 => n11141, B1 => n9444, B2 => 
                           n10047, ZN => n15778);
   U3487 : AOI22_X1 port map( A1 => n9348, A2 => n10050, B1 => n9316, B2 => 
                           n11138, ZN => n15777);
   U3488 : AOI22_X1 port map( A1 => n9284, A2 => n11152, B1 => n9188, B2 => 
                           n10051, ZN => n15776);
   U3489 : AOI22_X1 port map( A1 => n9508, A2 => n11136, B1 => n9252, B2 => 
                           n11132, ZN => n15775);
   U3490 : NAND4_X1 port map( A1 => n15778, A2 => n15777, A3 => n15776, A4 => 
                           n15775, ZN => n15779);
   U3491 : NOR2_X1 port map( A1 => n15780, A2 => n15779, ZN => n15792);
   U3492 : AOI22_X1 port map( A1 => n9892, A2 => n11144, B1 => n9796, B2 => 
                           n16077, ZN => n15784);
   U3493 : AOI22_X1 port map( A1 => n10020, A2 => n16072, B1 => n9988, B2 => 
                           n11228, ZN => n15783);
   U3494 : AOI22_X1 port map( A1 => n9924, A2 => n11135, B1 => n9828, B2 => 
                           n11147, ZN => n15782);
   U3495 : AOI22_X1 port map( A1 => n9860, A2 => n11131, B1 => n9956, B2 => 
                           n16048, ZN => n15781);
   U3496 : NAND4_X1 port map( A1 => n15784, A2 => n15783, A3 => n15782, A4 => 
                           n15781, ZN => n15790);
   U3497 : AOI22_X1 port map( A1 => n9604, A2 => n16078, B1 => n9668, B2 => 
                           n11232, ZN => n15788);
   U3498 : AOI22_X1 port map( A1 => n9540, A2 => n16077, B1 => n9572, B2 => 
                           n11127, ZN => n15787);
   U3499 : AOI22_X1 port map( A1 => n9764, A2 => n11231, B1 => n9700, B2 => 
                           n11230, ZN => n15786);
   U3500 : AOI22_X1 port map( A1 => n9732, A2 => n11228, B1 => n9636, B2 => 
                           n11144, ZN => n15785);
   U3501 : NAND4_X1 port map( A1 => n15788, A2 => n15787, A3 => n15786, A4 => 
                           n15785, ZN => n15789);
   U3502 : AOI22_X1 port map( A1 => n15880, A2 => n15790, B1 => n16085, B2 => 
                           n15789, ZN => n15791);
   U3503 : OAI21_X1 port map( B1 => n16090, B2 => n15792, A => n15791, ZN => 
                           OUT1(13));
   U3504 : AOI22_X1 port map( A1 => n9219, A2 => n11143, B1 => n9283, B2 => 
                           n11152, ZN => n15796);
   U3505 : AOI22_X1 port map( A1 => n9027, A2 => n11150, B1 => n9091, B2 => 
                           n10040, ZN => n15795);
   U3506 : AOI22_X1 port map( A1 => n9155, A2 => n11140, B1 => n9315, B2 => 
                           n11138, ZN => n15794);
   U3507 : AOI22_X1 port map( A1 => n9475, A2 => n11133, B1 => n9059, B2 => 
                           n11149, ZN => n15793);
   U3508 : NAND4_X1 port map( A1 => n15796, A2 => n15795, A3 => n15794, A4 => 
                           n15793, ZN => n15802);
   U3509 : AOI22_X1 port map( A1 => n9443, A2 => n11151, B1 => n9123, B2 => 
                           n10046, ZN => n15800);
   U3510 : AOI22_X1 port map( A1 => n9347, A2 => n10050, B1 => n9251, B2 => 
                           n10054, ZN => n15799);
   U3511 : AOI22_X1 port map( A1 => n9379, A2 => n11154, B1 => n9187, B2 => 
                           n10051, ZN => n15798);
   U3512 : AOI22_X1 port map( A1 => n9411, A2 => n10048, B1 => n9507, B2 => 
                           n11136, ZN => n15797);
   U3513 : NAND4_X1 port map( A1 => n15800, A2 => n15799, A3 => n15798, A4 => 
                           n15797, ZN => n15801);
   U3514 : NOR2_X1 port map( A1 => n15802, A2 => n15801, ZN => n15814);
   U3515 : AOI22_X1 port map( A1 => n9891, A2 => n11148, B1 => n9795, B2 => 
                           n11134, ZN => n15806);
   U3516 : AOI22_X1 port map( A1 => n9859, A2 => n11131, B1 => n9987, B2 => 
                           n11228, ZN => n15805);
   U3517 : AOI22_X1 port map( A1 => n9955, A2 => n11129, B1 => n9923, B2 => 
                           n16079, ZN => n15804);
   U3518 : AOI22_X1 port map( A1 => n9827, A2 => n11127, B1 => n10019, B2 => 
                           n11146, ZN => n15803);
   U3519 : NAND4_X1 port map( A1 => n15806, A2 => n15805, A3 => n15804, A4 => 
                           n15803, ZN => n15812);
   U3520 : AOI22_X1 port map( A1 => n9763, A2 => n16072, B1 => n9667, B2 => 
                           n11135, ZN => n15810);
   U3521 : AOI22_X1 port map( A1 => n9539, A2 => n16077, B1 => n9635, B2 => 
                           n11144, ZN => n15809);
   U3522 : AOI22_X1 port map( A1 => n9699, A2 => n11230, B1 => n9731, B2 => 
                           n11228, ZN => n15808);
   U3523 : AOI22_X1 port map( A1 => n9571, A2 => n11145, B1 => n9603, B2 => 
                           n11229, ZN => n15807);
   U3524 : NAND4_X1 port map( A1 => n15810, A2 => n15809, A3 => n15808, A4 => 
                           n15807, ZN => n15811);
   U3525 : AOI22_X1 port map( A1 => n15880, A2 => n15812, B1 => n16085, B2 => 
                           n15811, ZN => n15813);
   U3526 : OAI21_X1 port map( B1 => n16090, B2 => n15814, A => n15813, ZN => 
                           OUT1(12));
   U3527 : AOI22_X1 port map( A1 => n9090, A2 => n11142, B1 => n9186, B2 => 
                           n11153, ZN => n15818);
   U3528 : AOI22_X1 port map( A1 => n9282, A2 => n10049, B1 => n9218, B2 => 
                           n11143, ZN => n15817);
   U3529 : AOI22_X1 port map( A1 => n9154, A2 => n10041, B1 => n9378, B2 => 
                           n11154, ZN => n15816);
   U3530 : AOI22_X1 port map( A1 => n9314, A2 => n10044, B1 => n9122, B2 => 
                           n11137, ZN => n15815);
   U3531 : NAND4_X1 port map( A1 => n15818, A2 => n15817, A3 => n15816, A4 => 
                           n15815, ZN => n15824);
   U3532 : AOI22_X1 port map( A1 => n9442, A2 => n10047, B1 => n9410, B2 => 
                           n10048, ZN => n15822);
   U3533 : AOI22_X1 port map( A1 => n9250, A2 => n11132, B1 => n9026, B2 => 
                           n11150, ZN => n15821);
   U3534 : AOI22_X1 port map( A1 => n9346, A2 => n11139, B1 => n9058, B2 => 
                           n11149, ZN => n15820);
   U3535 : AOI22_X1 port map( A1 => n9474, A2 => n11133, B1 => n9506, B2 => 
                           n11136, ZN => n15819);
   U3536 : NAND4_X1 port map( A1 => n15822, A2 => n15821, A3 => n15820, A4 => 
                           n15819, ZN => n15823);
   U3537 : NOR2_X1 port map( A1 => n15824, A2 => n15823, ZN => n15837);
   U3538 : AOI22_X1 port map( A1 => n10018, A2 => n11231, B1 => n9890, B2 => 
                           n11144, ZN => n15828);
   U3539 : AOI22_X1 port map( A1 => n9826, A2 => n11145, B1 => n9986, B2 => 
                           n16053, ZN => n15827);
   U3540 : AOI22_X1 port map( A1 => n9858, A2 => n11229, B1 => n9922, B2 => 
                           n11232, ZN => n15826);
   U3541 : AOI22_X1 port map( A1 => n9794, A2 => n11134, B1 => n9954, B2 => 
                           n11230, ZN => n15825);
   U3542 : NAND4_X1 port map( A1 => n15828, A2 => n15827, A3 => n15826, A4 => 
                           n15825, ZN => n15834);
   U3543 : AOI22_X1 port map( A1 => n9730, A2 => n16053, B1 => n9634, B2 => 
                           n11144, ZN => n15832);
   U3544 : AOI22_X1 port map( A1 => n9602, A2 => n16078, B1 => n9538, B2 => 
                           n11225, ZN => n15831);
   U3545 : AOI22_X1 port map( A1 => n9698, A2 => n11129, B1 => n9570, B2 => 
                           n11145, ZN => n15830);
   U3546 : AOI22_X1 port map( A1 => n9762, A2 => n11146, B1 => n9666, B2 => 
                           n16079, ZN => n15829);
   U3547 : NAND4_X1 port map( A1 => n15832, A2 => n15831, A3 => n15830, A4 => 
                           n15829, ZN => n15833);
   U3548 : AOI22_X1 port map( A1 => n15835, A2 => n15834, B1 => n16085, B2 => 
                           n15833, ZN => n15836);
   U3549 : OAI21_X1 port map( B1 => n15905, B2 => n15837, A => n15836, ZN => 
                           OUT1(11));
   U3550 : AOI22_X1 port map( A1 => n9377, A2 => n10053, B1 => n9089, B2 => 
                           n11142, ZN => n15841);
   U3551 : AOI22_X1 port map( A1 => n9345, A2 => n11139, B1 => n9025, B2 => 
                           n11150, ZN => n15840);
   U3552 : AOI22_X1 port map( A1 => n9281, A2 => n11152, B1 => n9185, B2 => 
                           n11153, ZN => n15839);
   U3553 : AOI22_X1 port map( A1 => n9473, A2 => n11133, B1 => n9249, B2 => 
                           n10054, ZN => n15838);
   U3554 : NAND4_X1 port map( A1 => n15841, A2 => n15840, A3 => n15839, A4 => 
                           n15838, ZN => n15847);
   U3555 : AOI22_X1 port map( A1 => n9505, A2 => n11136, B1 => n9441, B2 => 
                           n11151, ZN => n15845);
   U3556 : AOI22_X1 port map( A1 => n9057, A2 => n11149, B1 => n9121, B2 => 
                           n10046, ZN => n15844);
   U3557 : AOI22_X1 port map( A1 => n9153, A2 => n11140, B1 => n9217, B2 => 
                           n10039, ZN => n15843);
   U3558 : AOI22_X1 port map( A1 => n9409, A2 => n10048, B1 => n9313, B2 => 
                           n11138, ZN => n15842);
   U3559 : NAND4_X1 port map( A1 => n15845, A2 => n15844, A3 => n15843, A4 => 
                           n15842, ZN => n15846);
   U3560 : NOR2_X1 port map( A1 => n15847, A2 => n15846, ZN => n15859);
   U3561 : AOI22_X1 port map( A1 => n9857, A2 => n16078, B1 => n10017, B2 => 
                           n11146, ZN => n15851);
   U3562 : AOI22_X1 port map( A1 => n9793, A2 => n11225, B1 => n9985, B2 => 
                           n11228, ZN => n15850);
   U3563 : AOI22_X1 port map( A1 => n9953, A2 => n11129, B1 => n9889, B2 => 
                           n11148, ZN => n15849);
   U3564 : AOI22_X1 port map( A1 => n9825, A2 => n11145, B1 => n9921, B2 => 
                           n11232, ZN => n15848);
   U3565 : NAND4_X1 port map( A1 => n15851, A2 => n15850, A3 => n15849, A4 => 
                           n15848, ZN => n15857);
   U3566 : AOI22_X1 port map( A1 => n9697, A2 => n11230, B1 => n9761, B2 => 
                           n11146, ZN => n15855);
   U3567 : AOI22_X1 port map( A1 => n9633, A2 => n11128, B1 => n9729, B2 => 
                           n11228, ZN => n15854);
   U3568 : AOI22_X1 port map( A1 => n9665, A2 => n11135, B1 => n9537, B2 => 
                           n11134, ZN => n15853);
   U3569 : AOI22_X1 port map( A1 => n9601, A2 => n11229, B1 => n9569, B2 => 
                           n11145, ZN => n15852);
   U3570 : NAND4_X1 port map( A1 => n15855, A2 => n15854, A3 => n15853, A4 => 
                           n15852, ZN => n15856);
   U3571 : AOI22_X1 port map( A1 => n15880, A2 => n15857, B1 => n16085, B2 => 
                           n15856, ZN => n15858);
   U3572 : OAI21_X1 port map( B1 => n15905, B2 => n15859, A => n15858, ZN => 
                           OUT1(10));
   U3573 : AOI22_X1 port map( A1 => n9376, A2 => n11154, B1 => n9344, B2 => 
                           n10050, ZN => n15863);
   U3574 : AOI22_X1 port map( A1 => n9152, A2 => n11140, B1 => n9440, B2 => 
                           n11151, ZN => n15862);
   U3575 : AOI22_X1 port map( A1 => n9120, A2 => n10046, B1 => n9248, B2 => 
                           n11132, ZN => n15861);
   U3576 : AOI22_X1 port map( A1 => n9408, A2 => n10048, B1 => n9504, B2 => 
                           n11136, ZN => n15860);
   U3577 : NAND4_X1 port map( A1 => n15863, A2 => n15862, A3 => n15861, A4 => 
                           n15860, ZN => n15869);
   U3578 : AOI22_X1 port map( A1 => n9088, A2 => n11142, B1 => n9280, B2 => 
                           n11152, ZN => n15867);
   U3579 : AOI22_X1 port map( A1 => n9024, A2 => n11150, B1 => n9184, B2 => 
                           n11153, ZN => n15866);
   U3580 : AOI22_X1 port map( A1 => n9216, A2 => n11143, B1 => n9472, B2 => 
                           n10042, ZN => n15865);
   U3581 : AOI22_X1 port map( A1 => n9312, A2 => n10044, B1 => n9056, B2 => 
                           n11149, ZN => n15864);
   U3582 : NAND4_X1 port map( A1 => n15867, A2 => n15866, A3 => n15865, A4 => 
                           n15864, ZN => n15868);
   U3583 : NOR2_X1 port map( A1 => n15869, A2 => n15868, ZN => n15882);
   U3584 : AOI22_X1 port map( A1 => n9984, A2 => n16053, B1 => n9888, B2 => 
                           n11144, ZN => n15873);
   U3585 : AOI22_X1 port map( A1 => n9792, A2 => n11225, B1 => n9824, B2 => 
                           n11145, ZN => n15872);
   U3586 : AOI22_X1 port map( A1 => n9856, A2 => n11229, B1 => n9952, B2 => 
                           n11230, ZN => n15871);
   U3587 : AOI22_X1 port map( A1 => n9920, A2 => n16079, B1 => n10016, B2 => 
                           n11146, ZN => n15870);
   U3588 : NAND4_X1 port map( A1 => n15873, A2 => n15872, A3 => n15871, A4 => 
                           n15870, ZN => n15879);
   U3589 : AOI22_X1 port map( A1 => n9600, A2 => n11229, B1 => n9568, B2 => 
                           n11147, ZN => n15877);
   U3590 : AOI22_X1 port map( A1 => n9536, A2 => n16077, B1 => n9760, B2 => 
                           n11146, ZN => n15876);
   U3591 : AOI22_X1 port map( A1 => n9664, A2 => n11135, B1 => n9728, B2 => 
                           n11228, ZN => n15875);
   U3592 : AOI22_X1 port map( A1 => n9696, A2 => n11230, B1 => n9632, B2 => 
                           n11144, ZN => n15874);
   U3593 : NAND4_X1 port map( A1 => n15877, A2 => n15876, A3 => n15875, A4 => 
                           n15874, ZN => n15878);
   U3594 : AOI22_X1 port map( A1 => n15880, A2 => n15879, B1 => n16085, B2 => 
                           n15878, ZN => n15881);
   U3595 : OAI21_X1 port map( B1 => n15905, B2 => n15882, A => n15881, ZN => 
                           OUT1(9));
   U3596 : AOI22_X1 port map( A1 => n9087, A2 => n11142, B1 => n9247, B2 => 
                           n11132, ZN => n15886);
   U3597 : AOI22_X1 port map( A1 => n9055, A2 => n11149, B1 => n9151, B2 => 
                           n11140, ZN => n15885);
   U3598 : AOI22_X1 port map( A1 => n9023, A2 => n11150, B1 => n9183, B2 => 
                           n10051, ZN => n15884);
   U3599 : AOI22_X1 port map( A1 => n9343, A2 => n11139, B1 => n9311, B2 => 
                           n11138, ZN => n15883);
   U3600 : NAND4_X1 port map( A1 => n15886, A2 => n15885, A3 => n15884, A4 => 
                           n15883, ZN => n15892);
   U3601 : AOI22_X1 port map( A1 => n9407, A2 => n11141, B1 => n9471, B2 => 
                           n11133, ZN => n15890);
   U3602 : AOI22_X1 port map( A1 => n9215, A2 => n10039, B1 => n9503, B2 => 
                           n10052, ZN => n15889);
   U3603 : AOI22_X1 port map( A1 => n9119, A2 => n10046, B1 => n9279, B2 => 
                           n11152, ZN => n15888);
   U3604 : AOI22_X1 port map( A1 => n9439, A2 => n11151, B1 => n9375, B2 => 
                           n10053, ZN => n15887);
   U3605 : NAND4_X1 port map( A1 => n15890, A2 => n15889, A3 => n15888, A4 => 
                           n15887, ZN => n15891);
   U3606 : NOR2_X1 port map( A1 => n15892, A2 => n15891, ZN => n15904);
   U3607 : AOI22_X1 port map( A1 => n9855, A2 => n11131, B1 => n9983, B2 => 
                           n16053, ZN => n15896);
   U3608 : AOI22_X1 port map( A1 => n9791, A2 => n11134, B1 => n10015, B2 => 
                           n11231, ZN => n15895);
   U3609 : AOI22_X1 port map( A1 => n9823, A2 => n11145, B1 => n9887, B2 => 
                           n11144, ZN => n15894);
   U3610 : AOI22_X1 port map( A1 => n9919, A2 => n11135, B1 => n9951, B2 => 
                           n11129, ZN => n15893);
   U3611 : NAND4_X1 port map( A1 => n15896, A2 => n15895, A3 => n15894, A4 => 
                           n15893, ZN => n15902);
   U3612 : AOI22_X1 port map( A1 => n9727, A2 => n11130, B1 => n9535, B2 => 
                           n11225, ZN => n15900);
   U3613 : AOI22_X1 port map( A1 => n9599, A2 => n16078, B1 => n9695, B2 => 
                           n11230, ZN => n15899);
   U3614 : AOI22_X1 port map( A1 => n9663, A2 => n11135, B1 => n9567, B2 => 
                           n11145, ZN => n15898);
   U3615 : AOI22_X1 port map( A1 => n9759, A2 => n11146, B1 => n9631, B2 => 
                           n11148, ZN => n15897);
   U3616 : NAND4_X1 port map( A1 => n15900, A2 => n15899, A3 => n15898, A4 => 
                           n15897, ZN => n15901);
   U3617 : AOI22_X1 port map( A1 => n16087, A2 => n15902, B1 => n16085, B2 => 
                           n15901, ZN => n15903);
   U3618 : OAI21_X1 port map( B1 => n15905, B2 => n15904, A => n15903, ZN => 
                           OUT1(8));
   U3619 : AOI22_X1 port map( A1 => n9086, A2 => n11142, B1 => n9246, B2 => 
                           n11132, ZN => n15909);
   U3620 : AOI22_X1 port map( A1 => n9054, A2 => n11149, B1 => n9406, B2 => 
                           n11141, ZN => n15908);
   U3621 : AOI22_X1 port map( A1 => n9438, A2 => n11151, B1 => n9374, B2 => 
                           n10053, ZN => n15907);
   U3622 : AOI22_X1 port map( A1 => n9118, A2 => n11137, B1 => n9278, B2 => 
                           n11152, ZN => n15906);
   U3623 : NAND4_X1 port map( A1 => n15909, A2 => n15908, A3 => n15907, A4 => 
                           n15906, ZN => n15915);
   U3624 : AOI22_X1 port map( A1 => n9310, A2 => n10044, B1 => n9182, B2 => 
                           n10051, ZN => n15913);
   U3625 : AOI22_X1 port map( A1 => n9342, A2 => n10050, B1 => n9150, B2 => 
                           n11140, ZN => n15912);
   U3626 : AOI22_X1 port map( A1 => n9502, A2 => n10052, B1 => n9470, B2 => 
                           n10042, ZN => n15911);
   U3627 : AOI22_X1 port map( A1 => n9214, A2 => n10039, B1 => n9022, B2 => 
                           n11150, ZN => n15910);
   U3628 : NAND4_X1 port map( A1 => n15913, A2 => n15912, A3 => n15911, A4 => 
                           n15910, ZN => n15914);
   U3629 : NOR2_X1 port map( A1 => n15915, A2 => n15914, ZN => n15927);
   U3630 : AOI22_X1 port map( A1 => n9790, A2 => n16077, B1 => n9918, B2 => 
                           n16079, ZN => n15919);
   U3631 : AOI22_X1 port map( A1 => n9982, A2 => n11130, B1 => n9950, B2 => 
                           n11129, ZN => n15918);
   U3632 : AOI22_X1 port map( A1 => n9886, A2 => n11148, B1 => n9822, B2 => 
                           n11147, ZN => n15917);
   U3633 : AOI22_X1 port map( A1 => n9854, A2 => n11229, B1 => n10014, B2 => 
                           n11231, ZN => n15916);
   U3634 : NAND4_X1 port map( A1 => n15919, A2 => n15918, A3 => n15917, A4 => 
                           n15916, ZN => n15925);
   U3635 : AOI22_X1 port map( A1 => n9662, A2 => n11232, B1 => n9630, B2 => 
                           n11128, ZN => n15923);
   U3636 : AOI22_X1 port map( A1 => n9534, A2 => n16077, B1 => n9694, B2 => 
                           n11129, ZN => n15922);
   U3637 : AOI22_X1 port map( A1 => n9758, A2 => n11231, B1 => n9598, B2 => 
                           n16078, ZN => n15921);
   U3638 : AOI22_X1 port map( A1 => n9726, A2 => n16053, B1 => n9566, B2 => 
                           n11147, ZN => n15920);
   U3639 : NAND4_X1 port map( A1 => n15923, A2 => n15922, A3 => n15921, A4 => 
                           n15920, ZN => n15924);
   U3640 : AOI22_X1 port map( A1 => n16087, A2 => n15925, B1 => n16085, B2 => 
                           n15924, ZN => n15926);
   U3641 : OAI21_X1 port map( B1 => n16090, B2 => n15927, A => n15926, ZN => 
                           OUT1(7));
   U3642 : AOI22_X1 port map( A1 => n9277, A2 => n11152, B1 => n9181, B2 => 
                           n10051, ZN => n15931);
   U3643 : AOI22_X1 port map( A1 => n9469, A2 => n11133, B1 => n9149, B2 => 
                           n10041, ZN => n15930);
   U3644 : AOI22_X1 port map( A1 => n9085, A2 => n10040, B1 => n9021, B2 => 
                           n10045, ZN => n15929);
   U3645 : AOI22_X1 port map( A1 => n9405, A2 => n11141, B1 => n9309, B2 => 
                           n11138, ZN => n15928);
   U3646 : NAND4_X1 port map( A1 => n15931, A2 => n15930, A3 => n15929, A4 => 
                           n15928, ZN => n15937);
   U3647 : AOI22_X1 port map( A1 => n9341, A2 => n11139, B1 => n9213, B2 => 
                           n10039, ZN => n15935);
   U3648 : AOI22_X1 port map( A1 => n9501, A2 => n11136, B1 => n9245, B2 => 
                           n11132, ZN => n15934);
   U3649 : AOI22_X1 port map( A1 => n9117, A2 => n11137, B1 => n9053, B2 => 
                           n10043, ZN => n15933);
   U3650 : AOI22_X1 port map( A1 => n9437, A2 => n10047, B1 => n9373, B2 => 
                           n11154, ZN => n15932);
   U3651 : NAND4_X1 port map( A1 => n15935, A2 => n15934, A3 => n15933, A4 => 
                           n15932, ZN => n15936);
   U3652 : NOR2_X1 port map( A1 => n15937, A2 => n15936, ZN => n15949);
   U3653 : AOI22_X1 port map( A1 => n9821, A2 => n11145, B1 => n9885, B2 => 
                           n11148, ZN => n15941);
   U3654 : AOI22_X1 port map( A1 => n9853, A2 => n16078, B1 => n9981, B2 => 
                           n11130, ZN => n15940);
   U3655 : AOI22_X1 port map( A1 => n9917, A2 => n11135, B1 => n9949, B2 => 
                           n16048, ZN => n15939);
   U3656 : AOI22_X1 port map( A1 => n10013, A2 => n11231, B1 => n9789, B2 => 
                           n11225, ZN => n15938);
   U3657 : NAND4_X1 port map( A1 => n15941, A2 => n15940, A3 => n15939, A4 => 
                           n15938, ZN => n15947);
   U3658 : AOI22_X1 port map( A1 => n9597, A2 => n11229, B1 => n9725, B2 => 
                           n11228, ZN => n15945);
   U3659 : AOI22_X1 port map( A1 => n9693, A2 => n11129, B1 => n9629, B2 => 
                           n11148, ZN => n15944);
   U3660 : AOI22_X1 port map( A1 => n9661, A2 => n11232, B1 => n9533, B2 => 
                           n11225, ZN => n15943);
   U3661 : AOI22_X1 port map( A1 => n9565, A2 => n11147, B1 => n9757, B2 => 
                           n11231, ZN => n15942);
   U3662 : NAND4_X1 port map( A1 => n15945, A2 => n15944, A3 => n15943, A4 => 
                           n15942, ZN => n15946);
   U3663 : AOI22_X1 port map( A1 => n16087, A2 => n15947, B1 => n16085, B2 => 
                           n15946, ZN => n15948);
   U3664 : OAI21_X1 port map( B1 => n16090, B2 => n15949, A => n15948, ZN => 
                           OUT1(6));
   U3665 : AOI22_X1 port map( A1 => n9340, A2 => n10050, B1 => n9468, B2 => 
                           n10042, ZN => n15953);
   U3666 : AOI22_X1 port map( A1 => n9116, A2 => n11137, B1 => n9436, B2 => 
                           n10047, ZN => n15952);
   U3667 : AOI22_X1 port map( A1 => n9500, A2 => n10052, B1 => n9084, B2 => 
                           n11142, ZN => n15951);
   U3668 : AOI22_X1 port map( A1 => n9404, A2 => n11141, B1 => n9244, B2 => 
                           n11132, ZN => n15950);
   U3669 : NAND4_X1 port map( A1 => n15953, A2 => n15952, A3 => n15951, A4 => 
                           n15950, ZN => n15959);
   U3670 : AOI22_X1 port map( A1 => n9020, A2 => n10045, B1 => n9212, B2 => 
                           n10039, ZN => n15957);
   U3671 : AOI22_X1 port map( A1 => n9148, A2 => n11140, B1 => n9052, B2 => 
                           n10043, ZN => n15956);
   U3672 : AOI22_X1 port map( A1 => n9180, A2 => n11153, B1 => n9308, B2 => 
                           n11138, ZN => n15955);
   U3673 : AOI22_X1 port map( A1 => n9372, A2 => n10053, B1 => n9276, B2 => 
                           n10049, ZN => n15954);
   U3674 : NAND4_X1 port map( A1 => n15957, A2 => n15956, A3 => n15955, A4 => 
                           n15954, ZN => n15958);
   U3675 : NOR2_X1 port map( A1 => n15959, A2 => n15958, ZN => n15971);
   U3676 : AOI22_X1 port map( A1 => n10012, A2 => n11231, B1 => n9980, B2 => 
                           n16053, ZN => n15963);
   U3677 : AOI22_X1 port map( A1 => n9820, A2 => n11147, B1 => n9948, B2 => 
                           n11129, ZN => n15962);
   U3678 : AOI22_X1 port map( A1 => n9852, A2 => n11229, B1 => n9916, B2 => 
                           n11232, ZN => n15961);
   U3679 : AOI22_X1 port map( A1 => n9884, A2 => n11148, B1 => n9788, B2 => 
                           n16077, ZN => n15960);
   U3680 : NAND4_X1 port map( A1 => n15963, A2 => n15962, A3 => n15961, A4 => 
                           n15960, ZN => n15969);
   U3681 : AOI22_X1 port map( A1 => n9596, A2 => n16078, B1 => n9692, B2 => 
                           n11129, ZN => n15967);
   U3682 : AOI22_X1 port map( A1 => n9564, A2 => n11147, B1 => n9628, B2 => 
                           n11128, ZN => n15966);
   U3683 : AOI22_X1 port map( A1 => n9660, A2 => n11135, B1 => n9756, B2 => 
                           n16072, ZN => n15965);
   U3684 : AOI22_X1 port map( A1 => n9532, A2 => n11225, B1 => n9724, B2 => 
                           n11130, ZN => n15964);
   U3685 : NAND4_X1 port map( A1 => n15967, A2 => n15966, A3 => n15965, A4 => 
                           n15964, ZN => n15968);
   U3686 : AOI22_X1 port map( A1 => n16087, A2 => n15969, B1 => n16085, B2 => 
                           n15968, ZN => n15970);
   U3687 : OAI21_X1 port map( B1 => n16090, B2 => n15971, A => n15970, ZN => 
                           OUT1(5));
   U3688 : AOI22_X1 port map( A1 => n9499, A2 => n10052, B1 => n9275, B2 => 
                           n11152, ZN => n15975);
   U3689 : AOI22_X1 port map( A1 => n9467, A2 => n10042, B1 => n9403, B2 => 
                           n11141, ZN => n15974);
   U3690 : AOI22_X1 port map( A1 => n9051, A2 => n11149, B1 => n9019, B2 => 
                           n10045, ZN => n15973);
   U3691 : AOI22_X1 port map( A1 => n9211, A2 => n10039, B1 => n9339, B2 => 
                           n10050, ZN => n15972);
   U3692 : NAND4_X1 port map( A1 => n15975, A2 => n15974, A3 => n15973, A4 => 
                           n15972, ZN => n15981);
   U3693 : AOI22_X1 port map( A1 => n9115, A2 => n11137, B1 => n9083, B2 => 
                           n11142, ZN => n15979);
   U3694 : AOI22_X1 port map( A1 => n9435, A2 => n11151, B1 => n9307, B2 => 
                           n10044, ZN => n15978);
   U3695 : AOI22_X1 port map( A1 => n9243, A2 => n11132, B1 => n9371, B2 => 
                           n10053, ZN => n15977);
   U3696 : AOI22_X1 port map( A1 => n9179, A2 => n10051, B1 => n9147, B2 => 
                           n11140, ZN => n15976);
   U3697 : NAND4_X1 port map( A1 => n15979, A2 => n15978, A3 => n15977, A4 => 
                           n15976, ZN => n15980);
   U3698 : NOR2_X1 port map( A1 => n15981, A2 => n15980, ZN => n15993);
   U3699 : AOI22_X1 port map( A1 => n9947, A2 => n11230, B1 => n9787, B2 => 
                           n11134, ZN => n15985);
   U3700 : AOI22_X1 port map( A1 => n9979, A2 => n11130, B1 => n9915, B2 => 
                           n11135, ZN => n15984);
   U3701 : AOI22_X1 port map( A1 => n10011, A2 => n16072, B1 => n9819, B2 => 
                           n11127, ZN => n15983);
   U3702 : AOI22_X1 port map( A1 => n9883, A2 => n11148, B1 => n9851, B2 => 
                           n11131, ZN => n15982);
   U3703 : NAND4_X1 port map( A1 => n15985, A2 => n15984, A3 => n15983, A4 => 
                           n15982, ZN => n15991);
   U3704 : AOI22_X1 port map( A1 => n9755, A2 => n16072, B1 => n9627, B2 => 
                           n11144, ZN => n15989);
   U3705 : AOI22_X1 port map( A1 => n9595, A2 => n16078, B1 => n9659, B2 => 
                           n11135, ZN => n15988);
   U3706 : AOI22_X1 port map( A1 => n9723, A2 => n16053, B1 => n9531, B2 => 
                           n16077, ZN => n15987);
   U3707 : AOI22_X1 port map( A1 => n9563, A2 => n11147, B1 => n9691, B2 => 
                           n11129, ZN => n15986);
   U3708 : NAND4_X1 port map( A1 => n15989, A2 => n15988, A3 => n15987, A4 => 
                           n15986, ZN => n15990);
   U3709 : AOI22_X1 port map( A1 => n16087, A2 => n15991, B1 => n16085, B2 => 
                           n15990, ZN => n15992);
   U3710 : OAI21_X1 port map( B1 => n16090, B2 => n15993, A => n15992, ZN => 
                           OUT1(4));
   U3711 : AOI22_X1 port map( A1 => n9082, A2 => n10040, B1 => n9146, B2 => 
                           n11140, ZN => n15997);
   U3712 : AOI22_X1 port map( A1 => n9114, A2 => n11137, B1 => n9178, B2 => 
                           n10051, ZN => n15996);
   U3713 : AOI22_X1 port map( A1 => n9050, A2 => n10043, B1 => n9210, B2 => 
                           n11143, ZN => n15995);
   U3714 : AOI22_X1 port map( A1 => n9018, A2 => n11150, B1 => n9370, B2 => 
                           n10053, ZN => n15994);
   U3715 : NAND4_X1 port map( A1 => n15997, A2 => n15996, A3 => n15995, A4 => 
                           n15994, ZN => n16003);
   U3716 : AOI22_X1 port map( A1 => n9498, A2 => n11136, B1 => n9466, B2 => 
                           n11133, ZN => n16001);
   U3717 : AOI22_X1 port map( A1 => n9402, A2 => n11141, B1 => n9434, B2 => 
                           n11151, ZN => n16000);
   U3718 : AOI22_X1 port map( A1 => n9274, A2 => n10049, B1 => n9338, B2 => 
                           n11139, ZN => n15999);
   U3719 : AOI22_X1 port map( A1 => n9242, A2 => n11132, B1 => n9306, B2 => 
                           n10044, ZN => n15998);
   U3720 : NAND4_X1 port map( A1 => n16001, A2 => n16000, A3 => n15999, A4 => 
                           n15998, ZN => n16002);
   U3721 : NOR2_X1 port map( A1 => n16003, A2 => n16002, ZN => n16015);
   U3722 : AOI22_X1 port map( A1 => n9946, A2 => n16048, B1 => n9786, B2 => 
                           n11225, ZN => n16007);
   U3723 : AOI22_X1 port map( A1 => n9850, A2 => n16078, B1 => n10010, B2 => 
                           n16072, ZN => n16006);
   U3724 : AOI22_X1 port map( A1 => n9818, A2 => n11147, B1 => n9914, B2 => 
                           n16079, ZN => n16005);
   U3725 : AOI22_X1 port map( A1 => n9882, A2 => n11128, B1 => n9978, B2 => 
                           n11130, ZN => n16004);
   U3726 : NAND4_X1 port map( A1 => n16007, A2 => n16006, A3 => n16005, A4 => 
                           n16004, ZN => n16013);
   U3727 : AOI22_X1 port map( A1 => n9594, A2 => n11229, B1 => n9530, B2 => 
                           n11225, ZN => n16011);
   U3728 : AOI22_X1 port map( A1 => n9626, A2 => n11144, B1 => n9690, B2 => 
                           n11129, ZN => n16010);
   U3729 : AOI22_X1 port map( A1 => n9658, A2 => n11232, B1 => n9754, B2 => 
                           n16072, ZN => n16009);
   U3730 : AOI22_X1 port map( A1 => n9722, A2 => n11130, B1 => n9562, B2 => 
                           n11147, ZN => n16008);
   U3731 : NAND4_X1 port map( A1 => n16011, A2 => n16010, A3 => n16009, A4 => 
                           n16008, ZN => n16012);
   U3732 : AOI22_X1 port map( A1 => n16087, A2 => n16013, B1 => n16085, B2 => 
                           n16012, ZN => n16014);
   U3733 : OAI21_X1 port map( B1 => n16090, B2 => n16015, A => n16014, ZN => 
                           OUT1(3));
   U3734 : AOI22_X1 port map( A1 => n9465, A2 => n11133, B1 => n9017, B2 => 
                           n10045, ZN => n16019);
   U3735 : AOI22_X1 port map( A1 => n9369, A2 => n11154, B1 => n9113, B2 => 
                           n11137, ZN => n16018);
   U3736 : AOI22_X1 port map( A1 => n9049, A2 => n11149, B1 => n9401, B2 => 
                           n11141, ZN => n16017);
   U3737 : AOI22_X1 port map( A1 => n9209, A2 => n10039, B1 => n9433, B2 => 
                           n11151, ZN => n16016);
   U3738 : NAND4_X1 port map( A1 => n16019, A2 => n16018, A3 => n16017, A4 => 
                           n16016, ZN => n16025);
   U3739 : AOI22_X1 port map( A1 => n9305, A2 => n11138, B1 => n9241, B2 => 
                           n10054, ZN => n16023);
   U3740 : AOI22_X1 port map( A1 => n9145, A2 => n10041, B1 => n9081, B2 => 
                           n11142, ZN => n16022);
   U3741 : AOI22_X1 port map( A1 => n9497, A2 => n10052, B1 => n9177, B2 => 
                           n10051, ZN => n16021);
   U3742 : AOI22_X1 port map( A1 => n9273, A2 => n10049, B1 => n9337, B2 => 
                           n10050, ZN => n16020);
   U3743 : NAND4_X1 port map( A1 => n16023, A2 => n16022, A3 => n16021, A4 => 
                           n16020, ZN => n16024);
   U3744 : NOR2_X1 port map( A1 => n16025, A2 => n16024, ZN => n16037);
   U3745 : AOI22_X1 port map( A1 => n9977, A2 => n11130, B1 => n9945, B2 => 
                           n11230, ZN => n16029);
   U3746 : AOI22_X1 port map( A1 => n9817, A2 => n11147, B1 => n9913, B2 => 
                           n11232, ZN => n16028);
   U3747 : AOI22_X1 port map( A1 => n10009, A2 => n11146, B1 => n9785, B2 => 
                           n11134, ZN => n16027);
   U3748 : AOI22_X1 port map( A1 => n9881, A2 => n11128, B1 => n9849, B2 => 
                           n11229, ZN => n16026);
   U3749 : NAND4_X1 port map( A1 => n16029, A2 => n16028, A3 => n16027, A4 => 
                           n16026, ZN => n16035);
   U3750 : AOI22_X1 port map( A1 => n9657, A2 => n11135, B1 => n9625, B2 => 
                           n11148, ZN => n16033);
   U3751 : AOI22_X1 port map( A1 => n9529, A2 => n11134, B1 => n9689, B2 => 
                           n11129, ZN => n16032);
   U3752 : AOI22_X1 port map( A1 => n9561, A2 => n11147, B1 => n9721, B2 => 
                           n11228, ZN => n16031);
   U3753 : AOI22_X1 port map( A1 => n9753, A2 => n16072, B1 => n9593, B2 => 
                           n16078, ZN => n16030);
   U3754 : NAND4_X1 port map( A1 => n16033, A2 => n16032, A3 => n16031, A4 => 
                           n16030, ZN => n16034);
   U3755 : AOI22_X1 port map( A1 => n16087, A2 => n16035, B1 => n16085, B2 => 
                           n16034, ZN => n16036);
   U3756 : OAI21_X1 port map( B1 => n16090, B2 => n16037, A => n16036, ZN => 
                           OUT1(2));
   U3757 : AOI22_X1 port map( A1 => n9336, A2 => n10050, B1 => n9080, B2 => 
                           n10040, ZN => n16041);
   U3758 : AOI22_X1 port map( A1 => n9432, A2 => n10047, B1 => n9400, B2 => 
                           n10048, ZN => n16040);
   U3759 : AOI22_X1 port map( A1 => n9272, A2 => n11152, B1 => n9176, B2 => 
                           n11153, ZN => n16039);
   U3760 : AOI22_X1 port map( A1 => n9112, A2 => n10046, B1 => n9496, B2 => 
                           n11136, ZN => n16038);
   U3761 : NAND4_X1 port map( A1 => n16041, A2 => n16040, A3 => n16039, A4 => 
                           n16038, ZN => n16047);
   U3762 : AOI22_X1 port map( A1 => n9464, A2 => n11133, B1 => n9048, B2 => 
                           n10043, ZN => n16045);
   U3763 : AOI22_X1 port map( A1 => n9208, A2 => n11143, B1 => n9016, B2 => 
                           n11150, ZN => n16044);
   U3764 : AOI22_X1 port map( A1 => n9368, A2 => n11154, B1 => n9144, B2 => 
                           n11140, ZN => n16043);
   U3765 : AOI22_X1 port map( A1 => n9240, A2 => n11132, B1 => n9304, B2 => 
                           n11138, ZN => n16042);
   U3766 : NAND4_X1 port map( A1 => n16045, A2 => n16044, A3 => n16043, A4 => 
                           n16042, ZN => n16046);
   U3767 : NOR2_X1 port map( A1 => n16047, A2 => n16046, ZN => n16061);
   U3768 : AOI22_X1 port map( A1 => n9912, A2 => n16079, B1 => n10008, B2 => 
                           n11231, ZN => n16052);
   U3769 : AOI22_X1 port map( A1 => n9848, A2 => n16078, B1 => n9976, B2 => 
                           n11228, ZN => n16051);
   U3770 : AOI22_X1 port map( A1 => n9816, A2 => n11147, B1 => n9944, B2 => 
                           n16048, ZN => n16050);
   U3771 : AOI22_X1 port map( A1 => n9784, A2 => n11225, B1 => n9880, B2 => 
                           n11148, ZN => n16049);
   U3772 : NAND4_X1 port map( A1 => n16052, A2 => n16051, A3 => n16050, A4 => 
                           n16049, ZN => n16059);
   U3773 : AOI22_X1 port map( A1 => n9688, A2 => n11129, B1 => n9592, B2 => 
                           n16078, ZN => n16057);
   U3774 : AOI22_X1 port map( A1 => n9624, A2 => n11128, B1 => n9656, B2 => 
                           n11135, ZN => n16056);
   U3775 : AOI22_X1 port map( A1 => n9528, A2 => n11225, B1 => n9720, B2 => 
                           n16053, ZN => n16055);
   U3776 : AOI22_X1 port map( A1 => n9560, A2 => n11145, B1 => n9752, B2 => 
                           n11146, ZN => n16054);
   U3777 : NAND4_X1 port map( A1 => n16057, A2 => n16056, A3 => n16055, A4 => 
                           n16054, ZN => n16058);
   U3778 : AOI22_X1 port map( A1 => n16087, A2 => n16059, B1 => n16085, B2 => 
                           n16058, ZN => n16060);
   U3779 : OAI21_X1 port map( B1 => n16090, B2 => n16061, A => n16060, ZN => 
                           OUT1(1));
   U3780 : AOI22_X1 port map( A1 => n9303, A2 => n11138, B1 => n9111, B2 => 
                           n11137, ZN => n16065);
   U3781 : AOI22_X1 port map( A1 => n9175, A2 => n10051, B1 => n9239, B2 => 
                           n10054, ZN => n16064);
   U3782 : AOI22_X1 port map( A1 => n9335, A2 => n11139, B1 => n9207, B2 => 
                           n11143, ZN => n16063);
   U3783 : AOI22_X1 port map( A1 => n9495, A2 => n10052, B1 => n9399, B2 => 
                           n10048, ZN => n16062);
   U3784 : NAND4_X1 port map( A1 => n16065, A2 => n16064, A3 => n16063, A4 => 
                           n16062, ZN => n16071);
   U3785 : AOI22_X1 port map( A1 => n9143, A2 => n10041, B1 => n9367, B2 => 
                           n11154, ZN => n16069);
   U3786 : AOI22_X1 port map( A1 => n9271, A2 => n10049, B1 => n9463, B2 => 
                           n11133, ZN => n16068);
   U3787 : AOI22_X1 port map( A1 => n9015, A2 => n11150, B1 => n9079, B2 => 
                           n11142, ZN => n16067);
   U3788 : AOI22_X1 port map( A1 => n9431, A2 => n11151, B1 => n9047, B2 => 
                           n10043, ZN => n16066);
   U3789 : NAND4_X1 port map( A1 => n16069, A2 => n16068, A3 => n16067, A4 => 
                           n16066, ZN => n16070);
   U3790 : NOR2_X1 port map( A1 => n16071, A2 => n16070, ZN => n16089);
   U3791 : AOI22_X1 port map( A1 => n9879, A2 => n11148, B1 => n9783, B2 => 
                           n11134, ZN => n16076);
   U3792 : AOI22_X1 port map( A1 => n10007, A2 => n16072, B1 => n9911, B2 => 
                           n11135, ZN => n16075);
   U3793 : AOI22_X1 port map( A1 => n9975, A2 => n11228, B1 => n9847, B2 => 
                           n16078, ZN => n16074);
   U3794 : AOI22_X1 port map( A1 => n9815, A2 => n11127, B1 => n9943, B2 => 
                           n11230, ZN => n16073);
   U3795 : NAND4_X1 port map( A1 => n16076, A2 => n16075, A3 => n16074, A4 => 
                           n16073, ZN => n16086);
   U3796 : AOI22_X1 port map( A1 => n9687, A2 => n11230, B1 => n9751, B2 => 
                           n11231, ZN => n16083);
   U3797 : AOI22_X1 port map( A1 => n9527, A2 => n16077, B1 => n9559, B2 => 
                           n11147, ZN => n16082);
   U3798 : AOI22_X1 port map( A1 => n9719, A2 => n11130, B1 => n9591, B2 => 
                           n16078, ZN => n16081);
   U3799 : AOI22_X1 port map( A1 => n9623, A2 => n11148, B1 => n9655, B2 => 
                           n16079, ZN => n16080);
   U3800 : NAND4_X1 port map( A1 => n16083, A2 => n16082, A3 => n16081, A4 => 
                           n16080, ZN => n16084);
   U3801 : AOI22_X1 port map( A1 => n16087, A2 => n16086, B1 => n16085, B2 => 
                           n16084, ZN => n16088);
   U3802 : OAI21_X1 port map( B1 => n16090, B2 => n16089, A => n16088, ZN => 
                           OUT1(0));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1808, n793, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, curr_instruction_to_cu_i_20_port, 
      curr_instruction_to_cu_i_19_port, curr_instruction_to_cu_i_18_port, 
      curr_instruction_to_cu_i_17_port, curr_instruction_to_cu_i_16_port, 
      curr_instruction_to_cu_i_15_port, curr_instruction_to_cu_i_14_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_4_port, curr_instruction_to_cu_i_3_port, 
      curr_instruction_to_cu_i_0_port, enable_rf_i, read_rf_p2_i, alu_cin_i, 
      write_rf_i, cu_i_n153, cu_i_n152, cu_i_n151, cu_i_n135, cu_i_n4, cu_i_n3,
      cu_i_n2, cu_i_n145, cu_i_cw2_4_port, cu_i_cw2_5_port, cu_i_cw2_6_port, 
      cu_i_cw2_7_port, cu_i_cw2_8_port, cu_i_cw1_5_port, cu_i_N279, cu_i_N278, 
      cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, cu_i_N273, cu_i_N267, 
      cu_i_N266, cu_i_N265, cu_i_N264, cu_i_cmd_alu_op_type_0_port, 
      cu_i_cmd_alu_op_type_1_port, cu_i_cmd_alu_op_type_2_port, 
      cu_i_cmd_alu_op_type_3_port, cu_i_cmd_word_3_port, cu_i_cmd_word_4_port, 
      cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, cu_i_cmd_word_8_port, 
      datapath_i_alu_output_val_i_0_port, datapath_i_alu_output_val_i_1_port, 
      datapath_i_alu_output_val_i_2_port, datapath_i_alu_output_val_i_3_port, 
      datapath_i_alu_output_val_i_4_port, datapath_i_alu_output_val_i_5_port, 
      datapath_i_alu_output_val_i_6_port, datapath_i_alu_output_val_i_7_port, 
      datapath_i_alu_output_val_i_8_port, datapath_i_alu_output_val_i_9_port, 
      datapath_i_alu_output_val_i_10_port, datapath_i_alu_output_val_i_11_port,
      datapath_i_alu_output_val_i_12_port, datapath_i_alu_output_val_i_13_port,
      datapath_i_alu_output_val_i_14_port, datapath_i_alu_output_val_i_15_port,
      datapath_i_alu_output_val_i_16_port, datapath_i_alu_output_val_i_17_port,
      datapath_i_alu_output_val_i_18_port, datapath_i_alu_output_val_i_19_port,
      datapath_i_alu_output_val_i_20_port, datapath_i_alu_output_val_i_21_port,
      datapath_i_alu_output_val_i_22_port, datapath_i_alu_output_val_i_23_port,
      datapath_i_alu_output_val_i_24_port, datapath_i_alu_output_val_i_25_port,
      datapath_i_alu_output_val_i_26_port, datapath_i_alu_output_val_i_27_port,
      datapath_i_alu_output_val_i_28_port, datapath_i_alu_output_val_i_29_port,
      datapath_i_alu_output_val_i_30_port, datapath_i_alu_output_val_i_31_port,
      datapath_i_val_immediate_i_0_port, datapath_i_val_immediate_i_1_port, 
      datapath_i_val_immediate_i_2_port, datapath_i_val_immediate_i_3_port, 
      datapath_i_val_immediate_i_4_port, datapath_i_val_immediate_i_5_port, 
      datapath_i_val_immediate_i_6_port, datapath_i_val_immediate_i_7_port, 
      datapath_i_val_immediate_i_8_port, datapath_i_val_immediate_i_9_port, 
      datapath_i_val_immediate_i_10_port, datapath_i_val_immediate_i_11_port, 
      datapath_i_val_immediate_i_12_port, datapath_i_val_immediate_i_13_port, 
      datapath_i_val_immediate_i_14_port, datapath_i_val_immediate_i_15_port, 
      datapath_i_val_immediate_i_16_port, datapath_i_val_immediate_i_17_port, 
      datapath_i_val_immediate_i_18_port, datapath_i_val_immediate_i_19_port, 
      datapath_i_val_immediate_i_20_port, datapath_i_val_immediate_i_21_port, 
      datapath_i_val_immediate_i_22_port, datapath_i_val_immediate_i_23_port, 
      datapath_i_val_immediate_i_24_port, datapath_i_val_immediate_i_25_port, 
      datapath_i_val_immediate_i_26_port, datapath_i_val_immediate_i_27_port, 
      datapath_i_val_immediate_i_28_port, datapath_i_val_immediate_i_29_port, 
      datapath_i_val_immediate_i_30_port, datapath_i_val_immediate_i_31_port, 
      datapath_i_val_b_i_0_port, datapath_i_val_b_i_1_port, 
      datapath_i_val_b_i_2_port, datapath_i_val_b_i_3_port, 
      datapath_i_val_b_i_4_port, datapath_i_val_b_i_5_port, 
      datapath_i_val_b_i_6_port, datapath_i_val_b_i_7_port, 
      datapath_i_val_b_i_8_port, datapath_i_val_b_i_9_port, 
      datapath_i_val_b_i_10_port, datapath_i_val_b_i_11_port, 
      datapath_i_val_b_i_12_port, datapath_i_val_b_i_13_port, 
      datapath_i_val_b_i_14_port, datapath_i_val_b_i_15_port, 
      datapath_i_val_b_i_16_port, datapath_i_val_b_i_17_port, 
      datapath_i_val_b_i_18_port, datapath_i_val_b_i_19_port, 
      datapath_i_val_b_i_20_port, datapath_i_val_b_i_21_port, 
      datapath_i_val_b_i_22_port, datapath_i_val_b_i_23_port, 
      datapath_i_val_b_i_24_port, datapath_i_val_b_i_25_port, 
      datapath_i_val_b_i_26_port, datapath_i_val_b_i_27_port, 
      datapath_i_val_b_i_28_port, datapath_i_val_b_i_29_port, 
      datapath_i_val_b_i_30_port, datapath_i_val_b_i_31_port, 
      datapath_i_val_a_i_0_port, datapath_i_val_a_i_1_port, 
      datapath_i_val_a_i_2_port, datapath_i_val_a_i_3_port, 
      datapath_i_val_a_i_4_port, datapath_i_val_a_i_5_port, 
      datapath_i_val_a_i_6_port, datapath_i_val_a_i_7_port, 
      datapath_i_val_a_i_8_port, datapath_i_val_a_i_9_port, 
      datapath_i_val_a_i_10_port, datapath_i_val_a_i_11_port, 
      datapath_i_val_a_i_12_port, datapath_i_val_a_i_13_port, 
      datapath_i_val_a_i_14_port, datapath_i_val_a_i_15_port, 
      datapath_i_val_a_i_16_port, datapath_i_val_a_i_17_port, 
      datapath_i_val_a_i_18_port, datapath_i_val_a_i_19_port, 
      datapath_i_val_a_i_20_port, datapath_i_val_a_i_21_port, 
      datapath_i_val_a_i_22_port, datapath_i_val_a_i_23_port, 
      datapath_i_val_a_i_24_port, datapath_i_val_a_i_25_port, 
      datapath_i_val_a_i_26_port, datapath_i_val_a_i_27_port, 
      datapath_i_val_a_i_28_port, datapath_i_val_a_i_29_port, 
      datapath_i_val_a_i_30_port, datapath_i_val_a_i_31_port, 
      datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_N40, 
      datapath_i_fetch_stage_dp_N39, datapath_i_decode_stage_dp_n44, 
      datapath_i_decode_stage_dp_n43, datapath_i_decode_stage_dp_n42, 
      datapath_i_decode_stage_dp_n41, datapath_i_decode_stage_dp_n40, 
      datapath_i_decode_stage_dp_n39, datapath_i_decode_stage_dp_n38, 
      datapath_i_decode_stage_dp_n37, datapath_i_decode_stage_dp_n36, 
      datapath_i_decode_stage_dp_n35, datapath_i_decode_stage_dp_n34, 
      datapath_i_decode_stage_dp_n33, datapath_i_decode_stage_dp_n32, 
      datapath_i_decode_stage_dp_n31, datapath_i_decode_stage_dp_n30, 
      datapath_i_decode_stage_dp_n29, datapath_i_decode_stage_dp_n28, 
      datapath_i_decode_stage_dp_n27, datapath_i_decode_stage_dp_n26, 
      datapath_i_decode_stage_dp_n25, datapath_i_decode_stage_dp_n24, 
      datapath_i_decode_stage_dp_n23, datapath_i_decode_stage_dp_n22, 
      datapath_i_decode_stage_dp_n21, datapath_i_decode_stage_dp_n20, 
      datapath_i_decode_stage_dp_n19, datapath_i_decode_stage_dp_n18, 
      datapath_i_decode_stage_dp_n17, datapath_i_decode_stage_dp_n16, 
      datapath_i_decode_stage_dp_n15, datapath_i_decode_stage_dp_n14, 
      datapath_i_decode_stage_dp_n13, datapath_i_decode_stage_dp_clk_immediate,
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, datapath_i_memory_stage_dp_n2, 
      n301, n302, n361, n375, n377, n380, n385, n390, n395, n400, n405, n415, 
      n420, n423, n426, n431, n436, n441, n464, n468, n474, n475, n477, n485, 
      n492, n493, n513, n514, n519, n523, n524, n526, n529, n535, n541, n547, 
      n553, n559, n565, n571, n577, n583, n589, n595, n601, n606, n676, n692, 
      n699, n700, n703, n705, n717, n719, n1301, n1302, n1303, n1304, n1305, 
      n1306, n1307, n1308, n1309, n1310, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1328, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1385, IRAM_ADDRESS_1_port, n1388, 
      IRAM_ADDRESS_0_port, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1916, n1429, IRAM_ADDRESS_29_port, n1431, IRAM_ADDRESS_27_port, 
      n1433, IRAM_ADDRESS_25_port, n1435, IRAM_ADDRESS_23_port, n1437, 
      IRAM_ADDRESS_21_port, n1439, IRAM_ADDRESS_19_port, n1441, 
      IRAM_ADDRESS_17_port, n1443, IRAM_ADDRESS_15_port, n1445, 
      IRAM_ADDRESS_13_port, n1447, IRAM_ADDRESS_11_port, n1449, 
      IRAM_ADDRESS_9_port, n1451, n1452, n1453, n1454, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_7_port, n1457, n1458, n1459, n1460, n1475, n1476, n1477, 
      n1478, n1485, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
      n1502, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, 
      IRAM_ENABLE_port, n1801, n1802, n1803, n1804, n1807, n1842, n1844, n1846,
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n2042, n2043, 
      n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, 
      n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, 
      n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, 
      n2074, n2075, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_3_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_28_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_22_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_16_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_10_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_4_port, n2275, 
      n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, 
      n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
      n2296, n2297, n2298, n2299, n2300, n2301, n2302, IRAM_ADDRESS_31_port, 
      n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, 
      n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
      n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
      n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, 
      n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, 
      n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, 
      n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
      n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, 
      n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, 
      n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, 
      n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, 
      n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, 
      n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, 
      n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, 
      n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, 
      n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
      n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, 
      n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, 
      n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
      n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
      n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, 
      n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
      n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, 
      n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, 
      n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, 
      n2575, n2576, n2577, n2578, n_3929, n_3930, n_3931, n_3932, n_3933, 
      n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, 
      n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, 
      n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, 
      n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, 
      n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, 
      n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, 
      n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, 
      n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, 
      n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014, 
      n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, 
      n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, 
      n_4033, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, 
      n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050, 
      n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, 
      n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, 
      n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, 
      n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, 
      n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, 
      n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, 
      n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, 
      n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122, 
      n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, 
      n_4132, n_4133, n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, 
      n_4141, n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, 
      n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158, 
      n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, 
      n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, 
      n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185, 
      n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193, n_4194, 
      n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, 
      n_4204, n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212, 
      n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, 
      n_4222, n_4223, n_4224, n_4225, n_4226, n_4227, n_4228, n_4229, n_4230, 
      n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, 
      n_4240, n_4241, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, 
      n_4249, n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, 
      n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, 
      n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, 
      n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, 
      n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, 
      n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301, n_4302, 
      n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, 
      n_4312, n_4313, n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, 
      n_4321, n_4322, n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, 
      n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, 
      n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346, n_4347, 
      n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, 
      n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, 
      n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, 
      n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383, 
      n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, 
      n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, 
      n_4402, n_4403, n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, 
      n_4411 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_n4);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_n2);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_n151);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_n152);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n1760, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n1760, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n1760, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n1760, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n1760, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n1760, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n1760, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n1760, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n1760, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n1760, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n1760, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n1760, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n1348, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n1348, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n1348, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n1348, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n1348, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n1760, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n1760, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n1760, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n1760, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n1760, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n1760, Z 
                           => DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n1760, Z 
                           => DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n1760, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n1760, Z 
                           => DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n1760, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n1760, Z 
                           => DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n1760, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n1760, Z 
                           => DRAM_ADDRESS_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n2578, D => n1390, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n301, D => n1391, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n301, D => n1392, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n301, D => n1393, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n2578, D => n1394, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n2578, D => n1395, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n2578, D => n1396, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n2578, D => n1397, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n2578, D => n1398, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n301, D => n1399, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n2578, D => n1400, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n2578, D => n1401, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n2578, D => n1402, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n2578, D => n1403, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n2578, D => n1404, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n2578, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n2578, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n2578, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n2578, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n301, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n2578, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n2578, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n2297, D => n1390, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n2575, D => n1391, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n2575, D => n1392, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n2297, D => n1393, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n2575, D => n1394, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n2297, D => n1395, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n2297, D => n1396, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n2575, D => n1397, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n2297, D => n1398, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n2575, D => n1399, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n2297, D => n1400, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n2575, D => n1401, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n2297, D => n1402, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n2575, D => n1403, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n2297, D => n1404, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n2297, D => n1405, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n2575, D => n1406, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n2297, D => n1407, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n2297, D => n1408, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n2297, D => n1409, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n2297, D => n1410, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n2297, D => n1411, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n2297, D => n1412, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n2297, D => n1413, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n2297, D => n1414, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n2297, D => n1415, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_26_inst : 
                           DLH_X1 port map( G => n2297, D => n1415, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_27_inst : 
                           DLH_X1 port map( G => n2297, D => n1415, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_28_inst : 
                           DLH_X1 port map( G => n2297, D => n1415, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_29_inst : 
                           DLH_X1 port map( G => n2297, D => n1415, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_30_inst : 
                           DLH_X1 port map( G => n2297, D => n1415, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n2297, D => n1415, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   clk_r_REG3253_S2 : DFFS_X1 port map( D => n361, CK => CLK, SN => RST, Q => 
                           n_3929, QN => DRAM_ENABLE);
   clk_r_REG1555_S9 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, CK => 
                           CLK, RN => RST, Q => n_3930, QN => n1854);
   clk_r_REG1463_S10 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, CK => 
                           CLK, RN => RST, Q => n_3931, QN => n1855);
   clk_r_REG115_S51 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, CK => 
                           CLK, RN => RST, Q => n_3932, QN => n1852);
   clk_r_REG104_S48 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, CK => 
                           CLK, RN => RST, Q => n_3933, QN => n1851);
   clk_r_REG90_S45 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, CK => 
                           CLK, RN => RST, Q => n_3934, QN => n1853);
   clk_r_REG78_S42 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, CK => 
                           CLK, RN => RST, Q => n_3935, QN => n1861);
   clk_r_REG163_S41 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, CK => 
                           CLK, RN => RST, Q => n_3936, QN => n1858);
   clk_r_REG66_S38 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, CK => 
                           CLK, RN => RST, Q => n_3937, QN => n1857);
   clk_r_REG55_S35 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, CK => 
                           CLK, RN => RST, Q => n_3938, QN => n1849);
   clk_r_REG40_S30 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, CK => 
                           CLK, RN => RST, Q => n_3939, QN => n1856);
   clk_r_REG293_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, CK => 
                           CLK, RN => RST, Q => n_3940, QN => n1850);
   clk_r_REG177_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, CK => 
                           CLK, RN => RST, Q => n_3941, QN => n1859);
   clk_r_REG406_S23 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, CK => 
                           CLK, RN => RST, Q => n_3942, QN => n1860);
   clk_r_REG460_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, CK => 
                           CLK, RN => RST, Q => n_3943, QN => n1848);
   clk_r_REG372_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, CK => 
                           CLK, RN => RST, Q => n_3944, QN => n1862);
   clk_r_REG902_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, CK => 
                           CLK, RN => RST, Q => n_3945, QN => n1847);
   clk_r_REG3181_S2 : DFFS_X1 port map( D => n793, CK => CLK, SN => RST, Q => 
                           IRAM_ENABLE_port, QN => n_3946);
   clk_r_REG2096_S4 : DFFS_X1 port map( D => n513, CK => CLK, SN => RST, Q => 
                           n1783, QN => n2550);
   clk_r_REG3486_S7 : DFFS_X1 port map( D => n2292, CK => CLK, SN => RST, Q => 
                           n1782, QN => n_3947);
   clk_r_REG3326_S1 : DFFR_X1 port map( D => n2578, CK => CLK, RN => RST, Q => 
                           n1781, QN => n_3948);
   clk_r_REG3476_S7 : DFFR_X1 port map( D => n2294, CK => CLK, RN => RST, Q => 
                           n1780, QN => n_3949);
   clk_r_REG3324_S3 : DFFR_X1 port map( D => n2254, CK => CLK, RN => RST, Q => 
                           n1779, QN => n_3950);
   clk_r_REG3261_S4 : DFFR_X1 port map( D => n2253, CK => CLK, RN => RST, Q => 
                           n1778, QN => n_3951);
   clk_r_REG3309_S1 : DFFR_X1 port map( D => n2575, CK => CLK, RN => RST, Q => 
                           n1777, QN => n_3952);
   clk_r_REG3296_S1 : DFFR_X1 port map( D => n2575, CK => CLK, RN => RST, Q => 
                           n1776, QN => n_3953);
   clk_r_REG3258_S2 : DFFR_X1 port map( D => n2252, CK => CLK, RN => RST, Q => 
                           DRAM_READNOTWRITE, QN => n_3954);
   clk_r_REG3274_S1 : DFFR_X1 port map( D => n2575, CK => CLK, RN => RST, Q => 
                           n1774, QN => n_3955);
   clk_r_REG3287_S2 : DFFR_X1 port map( D => n1774, CK => CLK, RN => RST, Q => 
                           n1773, QN => n_3956);
   clk_r_REG3284_S1 : DFFR_X1 port map( D => n2250, CK => CLK, RN => RST, Q => 
                           n1772, QN => n_3957);
   clk_r_REG3285_S2 : DFFR_X1 port map( D => n1772, CK => CLK, RN => RST, Q => 
                           n1771, QN => n_3958);
   clk_r_REG3286_S3 : DFFR_X1 port map( D => n1771, CK => CLK, RN => RST, Q => 
                           n1770, QN => n_3959);
   clk_r_REG3281_S1 : DFFR_X1 port map( D => n2249, CK => CLK, RN => RST, Q => 
                           n1769, QN => n_3960);
   clk_r_REG3282_S2 : DFFR_X1 port map( D => n1769, CK => CLK, RN => RST, Q => 
                           n1768, QN => n_3961);
   clk_r_REG3283_S3 : DFFR_X1 port map( D => n1768, CK => CLK, RN => RST, Q => 
                           n1767, QN => n_3962);
   clk_r_REG3278_S1 : DFFR_X1 port map( D => n2248, CK => CLK, RN => RST, Q => 
                           n1766, QN => n_3963);
   clk_r_REG3279_S2 : DFFR_X1 port map( D => n1766, CK => CLK, RN => RST, Q => 
                           n1765, QN => n_3964);
   clk_r_REG3280_S3 : DFFR_X1 port map( D => n1765, CK => CLK, RN => RST, Q => 
                           n1764, QN => n_3965);
   clk_r_REG3275_S1 : DFFR_X1 port map( D => n2247, CK => CLK, RN => RST, Q => 
                           n1763, QN => n_3966);
   clk_r_REG3276_S2 : DFFR_X1 port map( D => n1763, CK => CLK, RN => RST, Q => 
                           n1762, QN => n_3967);
   clk_r_REG3277_S3 : DFFR_X1 port map( D => n1762, CK => CLK, RN => RST, Q => 
                           n1761, QN => n_3968);
   clk_r_REG3254_S2 : DFFS_X1 port map( D => n361, CK => CLK, SN => RST, Q => 
                           n1760, QN => n_3969);
   clk_r_REG132_S4 : DFFR_X1 port map( D => n1310, CK => CLK, RN => RST, Q => 
                           n1759, QN => n_3970);
   clk_r_REG134_S4 : DFFS_X1 port map( D => n423, CK => CLK, SN => RST, Q => 
                           n1758, QN => n_3971);
   clk_r_REG2094_S5 : DFFR_X1 port map( D => n2280, CK => CLK, RN => RST, Q => 
                           n1757, QN => n_3972);
   clk_r_REG2093_S5 : DFFS_X1 port map( D => n2280, CK => CLK, SN => RST, Q => 
                           n1756, QN => n_3973);
   clk_r_REG740_S5 : DFFR_X1 port map( D => n2279, CK => CLK, RN => RST, Q => 
                           n1755, QN => n_3974);
   clk_r_REG2098_S4 : DFFS_X1 port map( D => n375, CK => CLK, SN => RST, Q => 
                           n1754, QN => n_3975);
   clk_r_REG2099_S5 : DFFS_X1 port map( D => n1754, CK => CLK, SN => RST, Q => 
                           n1753, QN => n_3976);
   clk_r_REG3019_S21 : DFFR_X1 port map( D => n2278, CK => CLK, RN => RST, Q =>
                           n1752, QN => n_3977);
   clk_r_REG3018_S21 : DFFS_X1 port map( D => n2278, CK => CLK, SN => RST, Q =>
                           n1751, QN => n_3978);
   clk_r_REG1458_S17 : DFFR_X1 port map( D => n2277, CK => CLK, RN => RST, Q =>
                           n1750, QN => n_3979);
   clk_r_REG1457_S17 : DFFS_X1 port map( D => n2277, CK => CLK, SN => RST, Q =>
                           n1749, QN => n_3980);
   clk_r_REG1712_S5 : DFFR_X1 port map( D => n2284, CK => CLK, RN => RST, Q => 
                           n1748, QN => n_3981);
   clk_r_REG1711_S5 : DFFS_X1 port map( D => n2284, CK => CLK, SN => RST, Q => 
                           n1747, QN => n_3982);
   clk_r_REG2100_S4 : DFFS_X1 port map( D => n375, CK => CLK, SN => RST, Q => 
                           n1746, QN => n_3983);
   clk_r_REG2101_S5 : DFFS_X1 port map( D => n1746, CK => CLK, SN => RST, Q => 
                           n1745, QN => n_3984);
   clk_r_REG2088_S5 : DFFR_X1 port map( D => n2283, CK => CLK, RN => RST, Q => 
                           n1744, QN => n_3985);
   clk_r_REG2087_S5 : DFFS_X1 port map( D => n2283, CK => CLK, SN => RST, Q => 
                           n1743, QN => n_3986);
   clk_r_REG2939_S33 : DFFR_X1 port map( D => n2285, CK => CLK, RN => RST, Q =>
                           n1742, QN => n_3987);
   clk_r_REG2938_S33 : DFFS_X1 port map( D => n2285, CK => CLK, SN => RST, Q =>
                           n1741, QN => n_3988);
   clk_r_REG2792_S36 : DFFR_X1 port map( D => n2286, CK => CLK, RN => RST, Q =>
                           n1740, QN => n_3989);
   clk_r_REG2791_S36 : DFFS_X1 port map( D => n2286, CK => CLK, SN => RST, Q =>
                           n1739, QN => n_3990);
   clk_r_REG1944_S39 : DFFR_X1 port map( D => n2287, CK => CLK, RN => RST, Q =>
                           n1738, QN => n_3991);
   clk_r_REG1943_S39 : DFFS_X1 port map( D => n2287, CK => CLK, SN => RST, Q =>
                           n1737, QN => n_3992);
   clk_r_REG2714_S40 : DFFR_X1 port map( D => n2282, CK => CLK, RN => RST, Q =>
                           n1736, QN => n_3993);
   clk_r_REG2713_S40 : DFFS_X1 port map( D => n2282, CK => CLK, SN => RST, Q =>
                           n1735, QN => n_3994);
   clk_r_REG2558_S43 : DFFR_X1 port map( D => n2281, CK => CLK, RN => RST, Q =>
                           n1734, QN => n_3995);
   clk_r_REG2557_S43 : DFFS_X1 port map( D => n2281, CK => CLK, SN => RST, Q =>
                           n1733, QN => n_3996);
   clk_r_REG2400_S46 : DFFR_X1 port map( D => n2276, CK => CLK, RN => RST, Q =>
                           n1732, QN => n_3997);
   clk_r_REG2399_S46 : DFFS_X1 port map( D => n2276, CK => CLK, SN => RST, Q =>
                           n1731, QN => n_3998);
   clk_r_REG2246_S49 : DFFR_X1 port map( D => n2275, CK => CLK, RN => RST, Q =>
                           n1730, QN => n_3999);
   clk_r_REG2245_S49 : DFFS_X1 port map( D => n2275, CK => CLK, SN => RST, Q =>
                           n1729, QN => n_4000);
   clk_r_REG3328_S1 : DFFS_X1 port map( D => n676, CK => CLK, SN => RST, Q => 
                           n1728, QN => n_4001);
   clk_r_REG3331_S2 : DFFR_X1 port map( D => n2288, CK => CLK, RN => RST, Q => 
                           n1726, QN => n2573);
   clk_r_REG3512_S4 : DFFR_X1 port map( D => n2246, CK => CLK, RN => RST, Q => 
                           n1725, QN => n_4002);
   clk_r_REG2169_S53 : DFFS_X1 port map( D => n1844, CK => CLK, SN => RST, Q =>
                           n1724, QN => n_4003);
   clk_r_REG3483_S7 : DFFS_X1 port map( D => n2298, CK => CLK, SN => RST, Q => 
                           n1723, QN => n_4004);
   clk_r_REG3489_S7 : DFFS_X1 port map( D => n2295, CK => CLK, SN => RST, Q => 
                           n1722, QN => n_4005);
   clk_r_REG3502_S7 : DFFS_X1 port map( D => n2291, CK => CLK, SN => RST, Q => 
                           n1721, QN => n_4006);
   clk_r_REG3507_S7 : DFFS_X1 port map( D => n2290, CK => CLK, SN => RST, Q => 
                           n1720, QN => n_4007);
   clk_r_REG3509_S7 : DFFS_X1 port map( D => n2289, CK => CLK, SN => RST, Q => 
                           n1719, QN => n_4008);
   clk_r_REG109_S49 : DFFS_X1 port map( D => n2275, CK => CLK, SN => RST, Q => 
                           n1718, QN => n_4009);
   clk_r_REG98_S46 : DFFS_X1 port map( D => n2276, CK => CLK, SN => RST, Q => 
                           n1717, QN => n_4010);
   clk_r_REG83_S43 : DFFS_X1 port map( D => n2281, CK => CLK, SN => RST, Q => 
                           n1716, QN => n_4011);
   clk_r_REG73_S40 : DFFS_X1 port map( D => n2282, CK => CLK, SN => RST, Q => 
                           n1715, QN => n_4012);
   clk_r_REG158_S39 : DFFS_X1 port map( D => n2287, CK => CLK, SN => RST, Q => 
                           n1714, QN => n_4013);
   clk_r_REG59_S36 : DFFS_X1 port map( D => n2286, CK => CLK, SN => RST, Q => 
                           n1713, QN => n_4014);
   clk_r_REG48_S33 : DFFS_X1 port map( D => n2285, CK => CLK, SN => RST, Q => 
                           n1712, QN => n_4015);
   clk_r_REG147_S5 : DFFS_X1 port map( D => n2283, CK => CLK, SN => RST, Q => 
                           n1711, QN => n_4016);
   clk_r_REG238_S5 : DFFS_X1 port map( D => n2284, CK => CLK, SN => RST, Q => 
                           n1710, QN => n_4017);
   clk_r_REG331_S17 : DFFS_X1 port map( D => n2277, CK => CLK, SN => RST, Q => 
                           n1709, QN => n_4018);
   clk_r_REG29_S21 : DFFS_X1 port map( D => n2278, CK => CLK, SN => RST, Q => 
                           n1708, QN => n_4019);
   clk_r_REG136_S5 : DFFS_X1 port map( D => n2280, CK => CLK, SN => RST, Q => 
                           n1707, QN => n_4020);
   clk_r_REG470_S5 : DFFS_X1 port map( D => n2279, CK => CLK, SN => RST, Q => 
                           n1706, QN => n_4021);
   clk_r_REG2244_S52 : DFFS_X1 port map( D => n1887, CK => CLK, SN => RST, Q =>
                           n1705, QN => n_4022);
   clk_r_REG2320_S50 : DFFS_X1 port map( D => n1881, CK => CLK, SN => RST, Q =>
                           n1704, QN => n2568);
   clk_r_REG2398_S49 : DFFS_X1 port map( D => n1893, CK => CLK, SN => RST, Q =>
                           n1703, QN => n_4023);
   clk_r_REG2477_S47 : DFFS_X1 port map( D => n1882, CK => CLK, SN => RST, Q =>
                           n1702, QN => n2567);
   clk_r_REG2556_S46 : DFFS_X1 port map( D => n1886, CK => CLK, SN => RST, Q =>
                           n1701, QN => n_4024);
   clk_r_REG2635_S44 : DFFS_X1 port map( D => n1883, CK => CLK, SN => RST, Q =>
                           n1700, QN => n2556);
   clk_r_REG2712_S43 : DFFS_X1 port map( D => n1884, CK => CLK, SN => RST, Q =>
                           n1699, QN => n_4025);
   clk_r_REG1795_S43 : DFFS_X1 port map( D => n1879, CK => CLK, SN => RST, Q =>
                           n1698, QN => n2563);
   clk_r_REG1941_S42 : DFFS_X1 port map( D => n1880, CK => CLK, SN => RST, Q =>
                           n1697, QN => n_4026);
   clk_r_REG2716_S40 : DFFS_X1 port map( D => n1877, CK => CLK, SN => RST, Q =>
                           n1696, QN => n2558);
   clk_r_REG2790_S39 : DFFS_X1 port map( D => n1892, CK => CLK, SN => RST, Q =>
                           n1695, QN => n_4027);
   clk_r_REG2865_S37 : DFFS_X1 port map( D => n1878, CK => CLK, SN => RST, Q =>
                           n1694, QN => n2559);
   clk_r_REG2937_S36 : DFFS_X1 port map( D => n1885, CK => CLK, SN => RST, Q =>
                           n1693, QN => n_4028);
   clk_r_REG2016_S36 : DFFS_X1 port map( D => n1875, CK => CLK, SN => RST, Q =>
                           n1692, QN => n2560);
   clk_r_REG2942_S33 : DFFS_X1 port map( D => n1876, CK => CLK, SN => RST, Q =>
                           n1691, QN => n_4029);
   clk_r_REG1557_S9 : DFFS_X1 port map( D => n1872, CK => CLK, SN => RST, Q => 
                           n1690, QN => n2562);
   clk_r_REG1710_S8 : DFFS_X1 port map( D => n1871, CK => CLK, SN => RST, Q => 
                           n1689, QN => n_4030);
   clk_r_REG1379_S8 : DFFS_X1 port map( D => n1873, CK => CLK, SN => RST, Q => 
                           n1688, QN => n2561);
   clk_r_REG1719_S8 : DFFS_X1 port map( D => n1896, CK => CLK, SN => RST, Q => 
                           n1687, QN => n_4031);
   clk_r_REG998_S25 : DFFS_X1 port map( D => n1874, CK => CLK, SN => RST, Q => 
                           n1686, QN => n2566);
   clk_r_REG3017_S24 : DFFS_X1 port map( D => n1889, CK => CLK, SN => RST, Q =>
                           n1685, QN => n_4032);
   clk_r_REG744_S7 : DFFS_X1 port map( D => n1870, CK => CLK, SN => RST, Q => 
                           n1684, QN => n2565);
   clk_r_REG2092_S8 : DFFS_X1 port map( D => n1890, CK => CLK, SN => RST, Q => 
                           n1683, QN => n_4033);
   clk_r_REG901_S11 : DFFS_X1 port map( D => n1897, CK => CLK, SN => RST, Q => 
                           n1682, QN => n2564);
   clk_r_REG1220_S8 : DFFS_X1 port map( D => n1894, CK => CLK, SN => RST, Q => 
                           n1681, QN => n_4034);
   clk_r_REG519_S8 : DFFS_X1 port map( D => n1895, CK => CLK, SN => RST, Q => 
                           n1680, QN => n2557);
   clk_r_REG1462_S11 : DFFS_X1 port map( D => n1869, CK => CLK, SN => RST, Q =>
                           n1679, QN => n_4035);
   clk_r_REG1464_S11 : DFFS_X1 port map( D => n1867, CK => CLK, SN => RST, Q =>
                           n1678, QN => n_4036);
   clk_r_REG1484_S11 : DFFS_X1 port map( D => n1868, CK => CLK, SN => RST, Q =>
                           n1677, QN => n_4037);
   clk_r_REG3036_S15 : DFFS_X1 port map( D => n1891, CK => CLK, SN => RST, Q =>
                           n1676, QN => n_4038);
   clk_r_REG3111_S13 : DFFS_X1 port map( D => n1888, CK => CLK, SN => RST, Q =>
                           n1675, QN => n_4039);
   clk_r_REG3335_S6 : DFFR_X1 port map( D => n719, CK => CLK, RN => RST, Q => 
                           n_4040, QN => n1674);
   clk_r_REG129_S3 : DFFR_X1 port map( D => n1673, CK => CLK, RN => RST, Q => 
                           n1672, QN => n_4041);
   clk_r_REG2180_S2 : DFF_X1 port map( D => datapath_i_val_a_i_30_port, CK => 
                           CLK, Q => n1671, QN => n_4042);
   clk_r_REG2181_S3 : DFFR_X1 port map( D => n1671, CK => CLK, RN => RST, Q => 
                           n1670, QN => n_4043);
   clk_r_REG2256_S2 : DFF_X1 port map( D => datapath_i_val_a_i_29_port, CK => 
                           CLK, Q => n1669, QN => n_4044);
   clk_r_REG2257_S3 : DFFR_X1 port map( D => n1669, CK => CLK, RN => RST, Q => 
                           n1668, QN => n_4045);
   clk_r_REG2332_S2 : DFF_X1 port map( D => datapath_i_val_a_i_28_port, CK => 
                           CLK, Q => n1667, QN => n_4046);
   clk_r_REG2333_S3 : DFFR_X1 port map( D => n1667, CK => CLK, RN => RST, Q => 
                           n1666, QN => n_4047);
   clk_r_REG2413_S2 : DFF_X1 port map( D => datapath_i_val_a_i_27_port, CK => 
                           CLK, Q => n1665, QN => n_4048);
   clk_r_REG2414_S3 : DFFR_X1 port map( D => n1665, CK => CLK, RN => RST, Q => 
                           n1664, QN => n_4049);
   clk_r_REG2491_S2 : DFF_X1 port map( D => datapath_i_val_a_i_26_port, CK => 
                           CLK, Q => n1663, QN => n_4050);
   clk_r_REG2492_S3 : DFFR_X1 port map( D => n1663, CK => CLK, RN => RST, Q => 
                           n1662, QN => n_4051);
   clk_r_REG2571_S2 : DFF_X1 port map( D => datapath_i_val_a_i_25_port, CK => 
                           CLK, Q => n1661, QN => n_4052);
   clk_r_REG2572_S3 : DFFR_X1 port map( D => n1661, CK => CLK, RN => RST, Q => 
                           n1660, QN => n_4053);
   clk_r_REG2647_S2 : DFF_X1 port map( D => datapath_i_val_a_i_24_port, CK => 
                           CLK, Q => n1659, QN => n_4054);
   clk_r_REG2648_S3 : DFFR_X1 port map( D => n1659, CK => CLK, RN => RST, Q => 
                           n1658, QN => n_4055);
   clk_r_REG1803_S2 : DFF_X1 port map( D => datapath_i_val_a_i_23_port, CK => 
                           CLK, Q => n1657, QN => n_4056);
   clk_r_REG1804_S3 : DFFR_X1 port map( D => n1657, CK => CLK, RN => RST, Q => 
                           n1656, QN => n_4057);
   clk_r_REG1877_S2 : DFF_X1 port map( D => datapath_i_val_a_i_22_port, CK => 
                           CLK, Q => n1655, QN => n_4058);
   clk_r_REG1878_S3 : DFFR_X1 port map( D => n1655, CK => CLK, RN => RST, Q => 
                           n1654, QN => n_4059);
   clk_r_REG1952_S2 : DFF_X1 port map( D => datapath_i_val_a_i_21_port, CK => 
                           CLK, Q => n1653, QN => n_4060);
   clk_r_REG1953_S3 : DFFR_X1 port map( D => n1653, CK => CLK, RN => RST, Q => 
                           n1652, QN => n_4061);
   clk_r_REG2726_S2 : DFF_X1 port map( D => datapath_i_val_a_i_20_port, CK => 
                           CLK, Q => n1651, QN => n_4062);
   clk_r_REG2727_S3 : DFFR_X1 port map( D => n1651, CK => CLK, RN => RST, Q => 
                           n1650, QN => n_4063);
   clk_r_REG2801_S2 : DFF_X1 port map( D => datapath_i_val_a_i_19_port, CK => 
                           CLK, Q => n1649, QN => n_4064);
   clk_r_REG2802_S3 : DFFR_X1 port map( D => n1649, CK => CLK, RN => RST, Q => 
                           n1648, QN => n_4065);
   clk_r_REG2873_S2 : DFF_X1 port map( D => datapath_i_val_a_i_18_port, CK => 
                           CLK, Q => n1647, QN => n_4066);
   clk_r_REG2874_S3 : DFFR_X1 port map( D => n1647, CK => CLK, RN => RST, Q => 
                           n1646, QN => n_4067);
   clk_r_REG2023_S2 : DFF_X1 port map( D => datapath_i_val_a_i_17_port, CK => 
                           CLK, Q => n1645, QN => n_4068);
   clk_r_REG2024_S3 : DFFR_X1 port map( D => n1645, CK => CLK, RN => RST, Q => 
                           n1644, QN => n_4069);
   clk_r_REG2950_S2 : DFF_X1 port map( D => datapath_i_val_a_i_16_port, CK => 
                           CLK, Q => n1643, QN => n_4070);
   clk_r_REG2951_S3 : DFFR_X1 port map( D => n1643, CK => CLK, RN => RST, Q => 
                           n1642, QN => n_4071);
   clk_r_REG1569_S2 : DFF_X1 port map( D => datapath_i_val_a_i_15_port, CK => 
                           CLK, Q => n1641, QN => n_4072);
   clk_r_REG1570_S3 : DFFR_X1 port map( D => n1641, CK => CLK, RN => RST, Q => 
                           n1640, QN => n_4073);
   clk_r_REG1646_S2 : DFF_X1 port map( D => datapath_i_val_a_i_14_port, CK => 
                           CLK, Q => n1639, QN => n_4074);
   clk_r_REG1647_S3 : DFFR_X1 port map( D => n1639, CK => CLK, RN => RST, Q => 
                           n1638, QN => n_4075);
   clk_r_REG1393_S2 : DFF_X1 port map( D => datapath_i_val_a_i_13_port, CK => 
                           CLK, Q => n1637, QN => n_4076);
   clk_r_REG1394_S3 : DFFR_X1 port map( D => n1637, CK => CLK, RN => RST, Q => 
                           n1636, QN => n_4077);
   clk_r_REG1730_S2 : DFF_X1 port map( D => datapath_i_val_a_i_12_port, CK => 
                           CLK, Q => n1635, QN => n_4078);
   clk_r_REG1731_S3 : DFFR_X1 port map( D => n1635, CK => CLK, RN => RST, Q => 
                           n1634, QN => n_4079);
   clk_r_REG1009_S2 : DFF_X1 port map( D => datapath_i_val_a_i_11_port, CK => 
                           CLK, Q => n1633, QN => n_4080);
   clk_r_REG1010_S3 : DFFR_X1 port map( D => n1633, CK => CLK, RN => RST, Q => 
                           n1632, QN => n_4081);
   clk_r_REG1084_S2 : DFF_X1 port map( D => datapath_i_val_a_i_10_port, CK => 
                           CLK, Q => n1631, QN => n_4082);
   clk_r_REG1085_S3 : DFFR_X1 port map( D => n1631, CK => CLK, RN => RST, Q => 
                           n1630, QN => n_4083);
   clk_r_REG758_S2 : DFF_X1 port map( D => datapath_i_val_a_i_9_port, CK => CLK
                           , Q => n1629, QN => n_4084);
   clk_r_REG759_S3 : DFFR_X1 port map( D => n1629, CK => CLK, RN => RST, Q => 
                           n1628, QN => n_4085);
   clk_r_REG835_S2 : DFF_X1 port map( D => datapath_i_val_a_i_8_port, CK => CLK
                           , Q => n1627, QN => n_4086);
   clk_r_REG836_S3 : DFFR_X1 port map( D => n1627, CK => CLK, RN => RST, Q => 
                           n1626, QN => n_4087);
   clk_r_REG1148_S2 : DFF_X1 port map( D => datapath_i_val_a_i_7_port, CK => 
                           CLK, Q => n1625, QN => n_4088);
   clk_r_REG1149_S3 : DFFR_X1 port map( D => n1625, CK => CLK, RN => RST, Q => 
                           n1624, QN => n_4089);
   clk_r_REG1228_S2 : DFF_X1 port map( D => datapath_i_val_a_i_6_port, CK => 
                           CLK, Q => n1623, QN => n_4090);
   clk_r_REG1229_S3 : DFFR_X1 port map( D => n1623, CK => CLK, RN => RST, Q => 
                           n1622, QN => n_4091);
   clk_r_REG675_S2 : DFF_X1 port map( D => datapath_i_val_a_i_5_port, CK => CLK
                           , Q => n1621, QN => n_4092);
   clk_r_REG676_S3 : DFFR_X1 port map( D => n1621, CK => CLK, RN => RST, Q => 
                           n1620, QN => n_4093);
   clk_r_REG934_S2 : DFF_X1 port map( D => datapath_i_val_a_i_4_port, CK => CLK
                           , Q => n1619, QN => n_4094);
   clk_r_REG935_S3 : DFFR_X1 port map( D => n1619, CK => CLK, RN => RST, Q => 
                           n1618, QN => n_4095);
   clk_r_REG1303_S2 : DFF_X1 port map( D => datapath_i_val_a_i_3_port, CK => 
                           CLK, Q => n1617, QN => n_4096);
   clk_r_REG1304_S3 : DFFR_X1 port map( D => n1617, CK => CLK, RN => RST, Q => 
                           n1616, QN => n_4097);
   clk_r_REG1492_S2 : DFF_X1 port map( D => datapath_i_val_a_i_2_port, CK => 
                           CLK, Q => n1615, QN => n_4098);
   clk_r_REG3043_S2 : DFF_X1 port map( D => datapath_i_val_a_i_1_port, CK => 
                           CLK, Q => n1614, QN => n_4099);
   clk_r_REG3115_S2 : DFF_X1 port map( D => datapath_i_val_a_i_0_port, CK => 
                           CLK, Q => n1613, QN => n_4100);
   clk_r_REG123_S1 : DFF_X1 port map( D => datapath_i_val_b_i_31_port, CK => 
                           CLK, Q => n1612, QN => n_4101);
   clk_r_REG124_S2 : DFFR_X1 port map( D => n1612, CK => CLK, RN => RST, Q => 
                           n1611, QN => n_4102);
   clk_r_REG125_S3 : DFFR_X1 port map( D => n1611, CK => CLK, RN => RST, Q => 
                           n1610, QN => n_4103);
   clk_r_REG2173_S1 : DFF_X1 port map( D => datapath_i_val_b_i_30_port, CK => 
                           CLK, Q => n1609, QN => n_4104);
   clk_r_REG2174_S2 : DFFR_X1 port map( D => n1609, CK => CLK, RN => RST, Q => 
                           n1608, QN => n_4105);
   clk_r_REG2175_S3 : DFFR_X1 port map( D => n1608, CK => CLK, RN => RST, Q => 
                           n1607, QN => n_4106);
   clk_r_REG2250_S1 : DFF_X1 port map( D => datapath_i_val_b_i_29_port, CK => 
                           CLK, Q => n1606, QN => n_4107);
   clk_r_REG2251_S2 : DFFR_X1 port map( D => n1606, CK => CLK, RN => RST, Q => 
                           n1605, QN => n_4108);
   clk_r_REG2252_S3 : DFFR_X1 port map( D => n1605, CK => CLK, RN => RST, Q => 
                           n1604, QN => n_4109);
   clk_r_REG2324_S1 : DFF_X1 port map( D => datapath_i_val_b_i_28_port, CK => 
                           CLK, Q => n1603, QN => n_4110);
   clk_r_REG2325_S2 : DFFR_X1 port map( D => n1603, CK => CLK, RN => RST, Q => 
                           n1602, QN => n_4111);
   clk_r_REG2326_S3 : DFFR_X1 port map( D => n1602, CK => CLK, RN => RST, Q => 
                           n1601, QN => n_4112);
   clk_r_REG2404_S1 : DFF_X1 port map( D => datapath_i_val_b_i_27_port, CK => 
                           CLK, Q => n1600, QN => n_4113);
   clk_r_REG2405_S2 : DFFR_X1 port map( D => n1600, CK => CLK, RN => RST, Q => 
                           n1599, QN => n_4114);
   clk_r_REG2406_S3 : DFFR_X1 port map( D => n1599, CK => CLK, RN => RST, Q => 
                           n1598, QN => n_4115);
   clk_r_REG2481_S1 : DFF_X1 port map( D => datapath_i_val_b_i_26_port, CK => 
                           CLK, Q => n1597, QN => n_4116);
   clk_r_REG2482_S2 : DFFR_X1 port map( D => n1597, CK => CLK, RN => RST, Q => 
                           n1596, QN => n_4117);
   clk_r_REG2483_S3 : DFFR_X1 port map( D => n1596, CK => CLK, RN => RST, Q => 
                           n1595, QN => n_4118);
   clk_r_REG2562_S1 : DFF_X1 port map( D => datapath_i_val_b_i_25_port, CK => 
                           CLK, Q => n1594, QN => n_4119);
   clk_r_REG2563_S2 : DFFR_X1 port map( D => n1594, CK => CLK, RN => RST, Q => 
                           n1593, QN => n_4120);
   clk_r_REG2564_S3 : DFFR_X1 port map( D => n1593, CK => CLK, RN => RST, Q => 
                           n1592, QN => n_4121);
   clk_r_REG2639_S1 : DFF_X1 port map( D => datapath_i_val_b_i_24_port, CK => 
                           CLK, Q => n1591, QN => n_4122);
   clk_r_REG2640_S2 : DFFR_X1 port map( D => n1591, CK => CLK, RN => RST, Q => 
                           n1590, QN => n_4123);
   clk_r_REG2641_S3 : DFFR_X1 port map( D => n1590, CK => CLK, RN => RST, Q => 
                           n1589, QN => n_4124);
   clk_r_REG1799_S1 : DFF_X1 port map( D => datapath_i_val_b_i_23_port, CK => 
                           CLK, Q => n1588, QN => n_4125);
   clk_r_REG1800_S2 : DFFR_X1 port map( D => n1588, CK => CLK, RN => RST, Q => 
                           n1587, QN => n_4126);
   clk_r_REG1801_S3 : DFFR_X1 port map( D => n1587, CK => CLK, RN => RST, Q => 
                           n1586, QN => n_4127);
   clk_r_REG1871_S1 : DFF_X1 port map( D => datapath_i_val_b_i_22_port, CK => 
                           CLK, Q => n1585, QN => n_4128);
   clk_r_REG1872_S2 : DFFR_X1 port map( D => n1585, CK => CLK, RN => RST, Q => 
                           n1584, QN => n_4129);
   clk_r_REG1873_S3 : DFFR_X1 port map( D => n1584, CK => CLK, RN => RST, Q => 
                           n1583, QN => n_4130);
   clk_r_REG1948_S1 : DFF_X1 port map( D => datapath_i_val_b_i_21_port, CK => 
                           CLK, Q => n1582, QN => n_4131);
   clk_r_REG1949_S2 : DFFR_X1 port map( D => n1582, CK => CLK, RN => RST, Q => 
                           n1581, QN => n_4132);
   clk_r_REG1950_S3 : DFFR_X1 port map( D => n1581, CK => CLK, RN => RST, Q => 
                           n1580, QN => n_4133);
   clk_r_REG2720_S1 : DFF_X1 port map( D => datapath_i_val_b_i_20_port, CK => 
                           CLK, Q => n1579, QN => n_4134);
   clk_r_REG2721_S2 : DFFR_X1 port map( D => n1579, CK => CLK, RN => RST, Q => 
                           n1578, QN => n_4135);
   clk_r_REG2722_S3 : DFFR_X1 port map( D => n1578, CK => CLK, RN => RST, Q => 
                           n1577, QN => n_4136);
   clk_r_REG2796_S1 : DFF_X1 port map( D => datapath_i_val_b_i_19_port, CK => 
                           CLK, Q => n1576, QN => n_4137);
   clk_r_REG2797_S2 : DFFR_X1 port map( D => n1576, CK => CLK, RN => RST, Q => 
                           n1575, QN => n_4138);
   clk_r_REG2798_S3 : DFFR_X1 port map( D => n1575, CK => CLK, RN => RST, Q => 
                           n1574, QN => n_4139);
   clk_r_REG2869_S1 : DFF_X1 port map( D => datapath_i_val_b_i_18_port, CK => 
                           CLK, Q => n1573, QN => n_4140);
   clk_r_REG2870_S2 : DFFR_X1 port map( D => n1573, CK => CLK, RN => RST, Q => 
                           n1572, QN => n_4141);
   clk_r_REG2871_S3 : DFFR_X1 port map( D => n1572, CK => CLK, RN => RST, Q => 
                           n1571, QN => n_4142);
   clk_r_REG2020_S1 : DFF_X1 port map( D => datapath_i_val_b_i_17_port, CK => 
                           CLK, Q => n1570, QN => n_4143);
   clk_r_REG2021_S2 : DFFR_X1 port map( D => n1570, CK => CLK, RN => RST, Q => 
                           n1569, QN => n_4144);
   clk_r_REG2022_S3 : DFFR_X1 port map( D => n1569, CK => CLK, RN => RST, Q => 
                           n1568, QN => n_4145);
   clk_r_REG2946_S1 : DFF_X1 port map( D => datapath_i_val_b_i_16_port, CK => 
                           CLK, Q => n1567, QN => n_4146);
   clk_r_REG2947_S2 : DFFR_X1 port map( D => n1567, CK => CLK, RN => RST, Q => 
                           n1566, QN => n_4147);
   clk_r_REG2948_S3 : DFFR_X1 port map( D => n1566, CK => CLK, RN => RST, Q => 
                           n1565, QN => n_4148);
   clk_r_REG1561_S1 : DFF_X1 port map( D => datapath_i_val_b_i_15_port, CK => 
                           CLK, Q => n1564, QN => n_4149);
   clk_r_REG1562_S2 : DFFR_X1 port map( D => n1564, CK => CLK, RN => RST, Q => 
                           n1563, QN => n_4150);
   clk_r_REG1563_S3 : DFFR_X1 port map( D => n1563, CK => CLK, RN => RST, Q => 
                           n1562, QN => n_4151);
   clk_r_REG1637_S1 : DFF_X1 port map( D => datapath_i_val_b_i_14_port, CK => 
                           CLK, Q => n1561, QN => n_4152);
   clk_r_REG1638_S2 : DFFR_X1 port map( D => n1561, CK => CLK, RN => RST, Q => 
                           n1560, QN => n_4153);
   clk_r_REG1639_S3 : DFFR_X1 port map( D => n1560, CK => CLK, RN => RST, Q => 
                           n1559, QN => n_4154);
   clk_r_REG1383_S1 : DFF_X1 port map( D => datapath_i_val_b_i_13_port, CK => 
                           CLK, Q => n1558, QN => n_4155);
   clk_r_REG1384_S2 : DFFR_X1 port map( D => n1558, CK => CLK, RN => RST, Q => 
                           n1557, QN => n_4156);
   clk_r_REG1385_S3 : DFFR_X1 port map( D => n1557, CK => CLK, RN => RST, Q => 
                           n1556, QN => n_4157);
   clk_r_REG1723_S1 : DFF_X1 port map( D => datapath_i_val_b_i_12_port, CK => 
                           CLK, Q => n1555, QN => n_4158);
   clk_r_REG1724_S2 : DFFR_X1 port map( D => n1555, CK => CLK, RN => RST, Q => 
                           n1554, QN => n_4159);
   clk_r_REG1725_S3 : DFFR_X1 port map( D => n1554, CK => CLK, RN => RST, Q => 
                           n1553, QN => n_4160);
   clk_r_REG1002_S1 : DFF_X1 port map( D => datapath_i_val_b_i_11_port, CK => 
                           CLK, Q => n1552, QN => n_4161);
   clk_r_REG1003_S2 : DFFR_X1 port map( D => n1552, CK => CLK, RN => RST, Q => 
                           n1551, QN => n_4162);
   clk_r_REG1004_S3 : DFFR_X1 port map( D => n1551, CK => CLK, RN => RST, Q => 
                           n1550, QN => n_4163);
   clk_r_REG1077_S1 : DFF_X1 port map( D => datapath_i_val_b_i_10_port, CK => 
                           CLK, Q => n1549, QN => n_4164);
   clk_r_REG1078_S2 : DFFR_X1 port map( D => n1549, CK => CLK, RN => RST, Q => 
                           n1548, QN => n_4165);
   clk_r_REG1079_S3 : DFFR_X1 port map( D => n1548, CK => CLK, RN => RST, Q => 
                           n1547, QN => n_4166);
   clk_r_REG748_S1 : DFF_X1 port map( D => datapath_i_val_b_i_9_port, CK => CLK
                           , Q => n1546, QN => n_4167);
   clk_r_REG749_S2 : DFFR_X1 port map( D => n1546, CK => CLK, RN => RST, Q => 
                           n1545, QN => n_4168);
   clk_r_REG750_S3 : DFFR_X1 port map( D => n1545, CK => CLK, RN => RST, Q => 
                           n1544, QN => n_4169);
   clk_r_REG826_S1 : DFF_X1 port map( D => datapath_i_val_b_i_8_port, CK => CLK
                           , Q => n1543, QN => n_4170);
   clk_r_REG827_S2 : DFFR_X1 port map( D => n1543, CK => CLK, RN => RST, Q => 
                           n1542, QN => n_4171);
   clk_r_REG828_S3 : DFFR_X1 port map( D => n1542, CK => CLK, RN => RST, Q => 
                           n1541, QN => n_4172);
   clk_r_REG387_S1 : DFF_X1 port map( D => datapath_i_val_b_i_7_port, CK => CLK
                           , Q => n1540, QN => n_4173);
   clk_r_REG388_S2 : DFFR_X1 port map( D => n1540, CK => CLK, RN => RST, Q => 
                           n1539, QN => n_4174);
   clk_r_REG389_S3 : DFFR_X1 port map( D => n1539, CK => CLK, RN => RST, Q => 
                           n1538, QN => n_4175);
   clk_r_REG1224_S1 : DFF_X1 port map( D => datapath_i_val_b_i_6_port, CK => 
                           CLK, Q => n1537, QN => n_4176);
   clk_r_REG1225_S2 : DFFR_X1 port map( D => n1537, CK => CLK, RN => RST, Q => 
                           n1536, QN => n_4177);
   clk_r_REG1226_S3 : DFFR_X1 port map( D => n1536, CK => CLK, RN => RST, Q => 
                           n1535, QN => n_4178);
   clk_r_REG523_S1 : DFF_X1 port map( D => datapath_i_val_b_i_5_port, CK => CLK
                           , Q => n1534, QN => n_4179);
   clk_r_REG524_S2 : DFFR_X1 port map( D => n1534, CK => CLK, RN => RST, Q => 
                           n1533, QN => n_4180);
   clk_r_REG525_S3 : DFFR_X1 port map( D => n1533, CK => CLK, RN => RST, Q => 
                           n1532, QN => n_4181);
   clk_r_REG907_S1 : DFF_X1 port map( D => datapath_i_val_b_i_4_port, CK => CLK
                           , Q => n1531, QN => n_4182);
   clk_r_REG908_S2 : DFFR_X1 port map( D => n1531, CK => CLK, RN => RST, Q => 
                           n1530, QN => n_4183);
   clk_r_REG909_S3 : DFFR_X1 port map( D => n1530, CK => CLK, RN => RST, Q => 
                           n1529, QN => n_4184);
   clk_r_REG360_S1 : DFF_X1 port map( D => datapath_i_val_b_i_3_port, CK => CLK
                           , Q => n1528, QN => n_4185);
   clk_r_REG361_S2 : DFFR_X1 port map( D => n1528, CK => CLK, RN => RST, Q => 
                           n1527, QN => n_4186);
   clk_r_REG362_S3 : DFFR_X1 port map( D => n1527, CK => CLK, RN => RST, Q => 
                           n1526, QN => n_4187);
   clk_r_REG1488_S1 : DFF_X1 port map( D => datapath_i_val_b_i_2_port, CK => 
                           CLK, Q => n1525, QN => n_4188);
   clk_r_REG1489_S2 : DFFR_X1 port map( D => n1525, CK => CLK, RN => RST, Q => 
                           n1524, QN => n_4189);
   clk_r_REG1490_S3 : DFFR_X1 port map( D => n1524, CK => CLK, RN => RST, Q => 
                           n1523, QN => n_4190);
   clk_r_REG3040_S1 : DFF_X1 port map( D => datapath_i_val_b_i_1_port, CK => 
                           CLK, Q => n1522, QN => n_4191);
   clk_r_REG3041_S2 : DFFR_X1 port map( D => n1522, CK => CLK, RN => RST, Q => 
                           n1521, QN => n_4192);
   clk_r_REG3042_S3 : DFFR_X1 port map( D => n1521, CK => CLK, RN => RST, Q => 
                           n1520, QN => n_4193);
   clk_r_REG0_S1 : DFF_X1 port map( D => datapath_i_val_b_i_0_port, CK => CLK, 
                           Q => n1519, QN => n_4194);
   clk_r_REG1_S2 : DFFR_X1 port map( D => n1519, CK => CLK, RN => RST, Q => 
                           n1518, QN => n_4195);
   clk_r_REG2_S3 : DFFR_X1 port map( D => n1518, CK => CLK, RN => RST, Q => 
                           n1517, QN => n_4196);
   clk_r_REG3472_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port, CK =>
                           CLK, RN => RST, Q => n1516, QN => n_4197);
   clk_r_REG3477_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port, CK =>
                           CLK, RN => RST, Q => n1515, QN => n_4198);
   clk_r_REG3471_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port, CK =>
                           CLK, RN => RST, Q => n1514, QN => n_4199);
   clk_r_REG3515_S4 : DFFR_X1 port map( D => cu_i_n4, CK => CLK, RN => RST, Q 
                           => n1513, QN => n_4200);
   clk_r_REG3332_S4 : DFFR_X1 port map( D => cu_i_n2, CK => CLK, RN => RST, Q 
                           => n1512, QN => n2551);
   clk_r_REG3513_S4 : DFFR_X1 port map( D => cu_i_n151, CK => CLK, RN => RST, Q
                           => n1511, QN => n2571);
   clk_r_REG3514_S4 : DFFR_X1 port map( D => cu_i_n152, CK => CLK, RN => RST, Q
                           => n1510, QN => n_4201);
   clk_r_REG3473_S9 : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port, CK =>
                           CLK, RN => RST, Q => n1508, QN => n_4202);
   clk_r_REG133_S4 : DFFS_X1 port map( D => n423, CK => CLK, SN => RST, Q => 
                           n1506, QN => n_4203);
   clk_r_REG2095_S4 : DFFS_X1 port map( D => n513, CK => CLK, SN => RST, Q => 
                           n1505, QN => n2549);
   clk_r_REG3329_S2 : DFFS_X1 port map( D => n2293, CK => CLK, SN => RST, Q => 
                           n_4204, QN => n1504);
   clk_r_REG3487_S7 : DFFS_X1 port map( D => n474, CK => CLK, SN => RST, Q => 
                           n_4205, QN => n1842);
   clk_r_REG3485_S7 : DFFS_X1 port map( D => n2292, CK => CLK, SN => RST, Q => 
                           n_4206, QN => n1502);
   clk_r_REG3480_S7 : DFFS_X1 port map( D => n2299, CK => CLK, SN => RST, Q => 
                           n_4207, QN => n1501);
   clk_r_REG3469_S7 : DFFR_X1 port map( D => n475, CK => CLK, RN => RST, Q => 
                           n1500, QN => n_4208);
   clk_r_REG3257_S2 : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => CLK, 
                           RN => RST, Q => n1499, QN => n_4209);
   clk_r_REG3259_S2 : DFFR_X1 port map( D => cu_i_cw1_5_port, CK => CLK, RN => 
                           RST, Q => n1498, QN => n_4210);
   clk_r_REG3255_S2 : DFFS_X1 port map( D => datapath_i_memory_stage_dp_n2, CK 
                           => CLK, SN => RST, Q => n1497, QN => n_4211);
   clk_r_REG3268_S1 : DFFR_X1 port map( D => cu_i_n135, CK => CLK, RN => RST, Q
                           => n1496, QN => n_4212);
   clk_r_REG3475_S7 : DFFS_X1 port map( D => n477, CK => CLK, SN => RST, Q => 
                           n1495, QN => n_4213);
   clk_r_REG427_S9 : DFFR_X1 port map( D => n526, CK => CLK, RN => RST, Q => 
                           n1494, QN => n_4214);
   clk_r_REG1556_S9 : DFFS_X1 port map( D => n514, CK => CLK, SN => RST, Q => 
                           n2555, QN => n1846);
   clk_r_REG428_S10 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_7_port, CK => CLK, RN
                           => RST, Q => n_4215, QN => n1897);
   clk_r_REG472_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_5_port, CK => CLK, RN
                           => RST, Q => n_4216, QN => n1895);
   clk_r_REG461_S6 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_9_port, CK => CLK, RN
                           => RST, Q => n_4217, QN => n1870);
   clk_r_REG407_S24 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_11_port, CK => CLK, 
                           RN => RST, Q => n_4218, QN => n1874);
   clk_r_REG333_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_13_port, CK => CLK, 
                           RN => RST, Q => n_4219, QN => n1873);
   clk_r_REG294_S8 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_15_port, CK => CLK, 
                           RN => RST, Q => n_4220, QN => n1872);
   clk_r_REG149_S35 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_17_port, CK => CLK, 
                           RN => RST, Q => n_4221, QN => n1875);
   clk_r_REG3330_S2 : DFFR_X1 port map( D => n2288, CK => CLK, RN => RST, Q => 
                           n_4222, QN => n1485);
   clk_r_REG56_S36 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_19_port, CK => CLK, 
                           RN => RST, Q => n_4223, QN => n1878);
   clk_r_REG67_S39 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_21_port, CK => CLK, 
                           RN => RST, Q => n_4224, QN => n1877);
   clk_r_REG164_S42 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_23_port, CK => CLK, 
                           RN => RST, Q => n_4225, QN => n1879);
   clk_r_REG79_S43 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_25_port, CK => CLK, 
                           RN => RST, Q => n_4226, QN => n1883);
   clk_r_REG91_S46 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_27_port, CK => CLK, 
                           RN => RST, Q => n_4227, QN => n1882);
   clk_r_REG105_S49 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_29_port, CK => CLK, 
                           RN => RST, Q => n_4228, QN => n1881);
   clk_r_REG3270_S1 : DFFR_X1 port map( D => n703, CK => CLK, RN => RST, Q => 
                           n1478, QN => n_4229);
   clk_r_REG3510_S7 : DFFR_X1 port map( D => n493, CK => CLK, RN => RST, Q => 
                           n1477, QN => n_4230);
   clk_r_REG3504_S7 : DFFS_X1 port map( D => n492, CK => CLK, SN => RST, Q => 
                           n1476, QN => n_4231);
   clk_r_REG3516_S2 : DFFR_X1 port map( D => cu_i_n3, CK => CLK, RN => RST, Q 
                           => n1475, QN => n_4232);
   clk_r_REG322_S10 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_4_port, CK => CLK, RN
                           => RST, Q => n_4233, QN => n1869);
   clk_r_REG374_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_6_port, CK => CLK, RN
                           => RST, Q => n_4234, QN => n1894);
   clk_r_REG138_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_8_port, CK => CLK, RN
                           => RST, Q => n_4235, QN => n1890);
   clk_r_REG31_S23 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_10_port, CK => CLK, 
                           RN => RST, Q => n_4236, QN => n1889);
   clk_r_REG179_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_12_port, CK => CLK, 
                           RN => RST, Q => n_4237, QN => n1896);
   clk_r_REG240_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_14_port, CK => CLK, 
                           RN => RST, Q => n_4238, QN => n1871);
   clk_r_REG42_S32 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_16_port, CK => CLK, 
                           RN => RST, Q => n_4239, QN => n1876);
   clk_r_REG50_S35 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_18_port, CK => CLK, 
                           RN => RST, Q => n_4240, QN => n1885);
   clk_r_REG61_S38 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_20_port, CK => CLK, 
                           RN => RST, Q => n_4241, QN => n1892);
   clk_r_REG160_S41 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_22_port, CK => CLK, 
                           RN => RST, Q => n_4242, QN => n1880);
   clk_r_REG75_S42 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_24_port, CK => CLK, 
                           RN => RST, Q => n_4243, QN => n1884);
   clk_r_REG85_S45 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_26_port, CK => CLK, 
                           RN => RST, Q => n_4244, QN => n1886);
   clk_r_REG100_S48 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_28_port, CK => CLK, 
                           RN => RST, Q => n_4245, QN => n1893);
   clk_r_REG111_S51 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_30_port, CK => CLK, 
                           RN => RST, Q => n_4246, QN => n1887);
   clk_r_REG119_S53 : DFFS_X1 port map( D => n606, CK => CLK, SN => RST, Q => 
                           n1460, QN => n_4247);
   clk_r_REG3251_S2 : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => CLK, 
                           RN => RST, Q => n1459, QN => n_4248);
   clk_r_REG3333_S4 : DFFS_X1 port map( D => cu_i_n145, CK => CLK, SN => RST, Q
                           => n1458, QN => n_4249);
   clk_r_REG320_S10 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_3_port, CK => 
                           CLK, RN => RST, Q => n1457, QN => n_4250);
   clk_r_REG135_S5 : DFFS_X1 port map( D => n2280, CK => CLK, SN => RST, Q => 
                           n_4251, QN => IRAM_ADDRESS_7_port);
   clk_r_REG469_S5 : DFFS_X1 port map( D => n2279, CK => CLK, SN => RST, Q => 
                           n_4252, QN => IRAM_ADDRESS_5_port);
   clk_r_REG425_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, CK => 
                           CLK, RN => RST, Q => n1454, QN => n_4253);
   clk_r_REG371_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, CK => 
                           CLK, RN => RST, Q => n1453, QN => n_4254);
   clk_r_REG3267_S1 : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK => CLK, 
                           RN => RST, Q => n1452, QN => n_4255);
   clk_r_REG426_S9 : DFFR_X1 port map( D => n519, CK => CLK, RN => RST, Q => 
                           n1451, QN => n_4256);
   clk_r_REG28_S21 : DFFS_X1 port map( D => n2278, CK => CLK, SN => RST, Q => 
                           n_4257, QN => IRAM_ADDRESS_9_port);
   clk_r_REG459_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, CK => 
                           CLK, RN => RST, Q => n1449, QN => n_4258);
   clk_r_REG330_S17 : DFFS_X1 port map( D => n2277, CK => CLK, SN => RST, Q => 
                           n_4259, QN => IRAM_ADDRESS_11_port);
   clk_r_REG405_S23 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, CK => 
                           CLK, RN => RST, Q => n1447, QN => n_4260);
   clk_r_REG237_S5 : DFFS_X1 port map( D => n2284, CK => CLK, SN => RST, Q => 
                           n_4261, QN => IRAM_ADDRESS_13_port);
   clk_r_REG176_S5 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, CK => 
                           CLK, RN => RST, Q => n1445, QN => n_4262);
   clk_r_REG146_S5 : DFFS_X1 port map( D => n2283, CK => CLK, SN => RST, Q => 
                           n_4263, QN => IRAM_ADDRESS_15_port);
   clk_r_REG292_S7 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, CK => 
                           CLK, RN => RST, Q => n1443, QN => n_4264);
   clk_r_REG47_S33 : DFFS_X1 port map( D => n2285, CK => CLK, SN => RST, Q => 
                           n_4265, QN => IRAM_ADDRESS_17_port);
   clk_r_REG39_S30 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, CK => 
                           CLK, RN => RST, Q => n1441, QN => n_4266);
   clk_r_REG58_S36 : DFFS_X1 port map( D => n2286, CK => CLK, SN => RST, Q => 
                           n_4267, QN => IRAM_ADDRESS_19_port);
   clk_r_REG54_S35 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, CK => 
                           CLK, RN => RST, Q => n1439, QN => n_4268);
   clk_r_REG157_S39 : DFFS_X1 port map( D => n2287, CK => CLK, SN => RST, Q => 
                           n_4269, QN => IRAM_ADDRESS_21_port);
   clk_r_REG65_S38 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, CK => 
                           CLK, RN => RST, Q => n1437, QN => n_4270);
   clk_r_REG72_S40 : DFFS_X1 port map( D => n2282, CK => CLK, SN => RST, Q => 
                           n_4271, QN => IRAM_ADDRESS_23_port);
   clk_r_REG162_S41 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, CK => 
                           CLK, RN => RST, Q => n1435, QN => n_4272);
   clk_r_REG82_S43 : DFFS_X1 port map( D => n2281, CK => CLK, SN => RST, Q => 
                           n_4273, QN => IRAM_ADDRESS_25_port);
   clk_r_REG77_S42 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, CK => 
                           CLK, RN => RST, Q => n1433, QN => n_4274);
   clk_r_REG97_S46 : DFFS_X1 port map( D => n2276, CK => CLK, SN => RST, Q => 
                           n_4275, QN => IRAM_ADDRESS_27_port);
   clk_r_REG89_S45 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, CK => 
                           CLK, RN => RST, Q => n1431, QN => n_4276);
   clk_r_REG108_S49 : DFFS_X1 port map( D => n2275, CK => CLK, SN => RST, Q => 
                           n_4277, QN => IRAM_ADDRESS_29_port);
   clk_r_REG103_S48 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, CK => 
                           CLK, RN => RST, Q => n1429, QN => n_4278);
   clk_r_REG118_S52 : DFFR_X1 port map( D => n1808, CK => CLK, RN => RST, Q => 
                           n1916, QN => n_4279);
   clk_r_REG114_S51 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, CK => 
                           CLK, RN => RST, Q => n1427, QN => n_4280);
   clk_r_REG3273_S2 : DFFR_X1 port map( D => cu_i_cw2_4_port, CK => CLK, RN => 
                           RST, Q => n1426, QN => n2569);
   clk_r_REG3262_S3 : DFFR_X1 port map( D => cu_i_cw2_7_port, CK => CLK, RN => 
                           RST, Q => n1425, QN => n_4281);
   clk_r_REG3263_S3 : DFFR_X1 port map( D => cu_i_cw2_8_port, CK => CLK, RN => 
                           RST, Q => n1424, QN => n_4282);
   clk_r_REG3323_S2 : DFFR_X1 port map( D => cu_i_cw2_6_port, CK => CLK, RN => 
                           RST, Q => n1423, QN => n_4283);
   clk_r_REG3260_S3 : DFFR_X1 port map( D => cu_i_cw2_5_port, CK => CLK, RN => 
                           RST, Q => n1422, QN => n_4284);
   clk_r_REG3178_S1 : DFFS_X1 port map( D => n2302, CK => CLK, SN => RST, Q => 
                           n_4285, QN => n1421);
   clk_r_REG3468_S7 : DFFS_X1 port map( D => n2301, CK => CLK, SN => RST, Q => 
                           n_4286, QN => n1420);
   clk_r_REG3481_S7 : DFFS_X1 port map( D => n2300, CK => CLK, SN => RST, Q => 
                           n_4287, QN => n1419);
   clk_r_REG3482_S7 : DFFS_X1 port map( D => n2298, CK => CLK, SN => RST, Q => 
                           n_4288, QN => n1418);
   clk_r_REG3484_S7 : DFFS_X1 port map( D => n2296, CK => CLK, SN => RST, Q => 
                           n_4289, QN => n1417);
   clk_r_REG3488_S7 : DFFS_X1 port map( D => n2295, CK => CLK, SN => RST, Q => 
                           n_4290, QN => n1416);
   clk_r_REG3490_S7 : DFFR_X1 port map( D => datapath_i_n9, CK => CLK, RN => 
                           RST, Q => n1415, QN => n_4291);
   clk_r_REG3492_S7 : DFFR_X1 port map( D => datapath_i_n10, CK => CLK, RN => 
                           RST, Q => n1414, QN => n_4292);
   clk_r_REG3337_S7 : DFFR_X1 port map( D => datapath_i_n11, CK => CLK, RN => 
                           RST, Q => n1413, QN => n_4293);
   clk_r_REG3388_S7 : DFFR_X1 port map( D => datapath_i_n12, CK => CLK, RN => 
                           RST, Q => n1412, QN => n_4294);
   clk_r_REG3389_S7 : DFFR_X1 port map( D => datapath_i_n13, CK => CLK, RN => 
                           RST, Q => n1411, QN => n_4295);
   clk_r_REG3390_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_20_port, 
                           CK => CLK, RN => RST, Q => n1410, QN => n_4296);
   clk_r_REG3424_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_19_port, 
                           CK => CLK, RN => RST, Q => n1409, QN => n_4297);
   clk_r_REG3427_S7 : DFFS_X1 port map( D => n2258, CK => CLK, SN => RST, Q => 
                           n_4298, QN => n1408);
   clk_r_REG3450_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_17_port, 
                           CK => CLK, RN => RST, Q => n1407, QN => n_4299);
   clk_r_REG3451_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_16_port, 
                           CK => CLK, RN => RST, Q => n1406, QN => n_4300);
   clk_r_REG3453_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_14_port, 
                           CK => CLK, RN => RST, Q => n1404, QN => n_4301);
   clk_r_REG3454_S7 : DFFS_X1 port map( D => n2257, CK => CLK, SN => RST, Q => 
                           n_4302, QN => n1403);
   clk_r_REG3455_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_12_port, 
                           CK => CLK, RN => RST, Q => n1402, QN => n_4303);
   clk_r_REG3495_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_11_port, 
                           CK => CLK, RN => RST, Q => n1401, QN => n_4304);
   clk_r_REG3496_S7 : DFFR_X1 port map( D => datapath_i_n14, CK => CLK, RN => 
                           RST, Q => n1400, QN => n_4305);
   clk_r_REG3497_S7 : DFFR_X1 port map( D => datapath_i_n15, CK => CLK, RN => 
                           RST, Q => n1399, QN => n_4306);
   clk_r_REG3498_S7 : DFFR_X1 port map( D => datapath_i_n16, CK => CLK, RN => 
                           RST, Q => n1398, QN => n_4307);
   clk_r_REG3499_S7 : DFFR_X1 port map( D => datapath_i_n17, CK => CLK, RN => 
                           RST, Q => n1397, QN => n_4308);
   clk_r_REG3500_S7 : DFFR_X1 port map( D => datapath_i_n18, CK => CLK, RN => 
                           RST, Q => n1396, QN => n_4309);
   clk_r_REG3501_S7 : DFFS_X1 port map( D => n2291, CK => CLK, SN => RST, Q => 
                           n_4310, QN => n1395);
   clk_r_REG3503_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_4_port, 
                           CK => CLK, RN => RST, Q => n1394, QN => n_4311);
   clk_r_REG3505_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_3_port, 
                           CK => CLK, RN => RST, Q => n1393, QN => n_4312);
   clk_r_REG3506_S7 : DFFS_X1 port map( D => n2290, CK => CLK, SN => RST, Q => 
                           n_4313, QN => n1392);
   clk_r_REG3508_S7 : DFFS_X1 port map( D => n2289, CK => CLK, SN => RST, Q => 
                           n2572, QN => n1391);
   clk_r_REG3511_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_0_port, 
                           CK => CLK, RN => RST, Q => n1390, QN => n2570);
   clk_r_REG10_S11 : DFFR_X1 port map( D => datapath_i_fetch_stage_dp_N39, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_0_port, QN => 
                           n_4314);
   clk_r_REG11_S11 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_0_port, CK => CLK, RN
                           => RST, Q => n1388, QN => n_4315);
   clk_r_REG3110_S12 : DFFR_X1 port map( D => n1388, CK => CLK, RN => RST, Q =>
                           n_4316, QN => n1888);
   clk_r_REG17_S13 : DFFR_X1 port map( D => datapath_i_fetch_stage_dp_N40, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_1_port, QN => 
                           n_4317);
   clk_r_REG18_S13 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_1_port, CK => CLK, RN
                           => RST, Q => n1385, QN => n_4318);
   clk_r_REG3035_S14 : DFFR_X1 port map( D => n1385, CK => CLK, RN => RST, Q =>
                           n_4319, QN => n1891);
   clk_r_REG3288_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1383, QN => n_4320);
   clk_r_REG3289_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1382, QN => n_4321);
   clk_r_REG3290_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1381, QN => n_4322);
   clk_r_REG3291_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1380, QN => n_4323);
   clk_r_REG3292_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1379, QN => n_4324);
   clk_r_REG3293_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1378, QN => n_4325);
   clk_r_REG3294_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1377, QN => n_4326);
   clk_r_REG3295_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1376, QN => n_4327);
   clk_r_REG3297_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1375, QN => n_4328);
   clk_r_REG3298_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1374, QN => n_4329);
   clk_r_REG3299_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1373, QN => n_4330);
   clk_r_REG3300_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1372, QN => n_4331);
   clk_r_REG3301_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1371, QN => n_4332);
   clk_r_REG3302_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1370, QN => n_4333);
   clk_r_REG3303_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1369, QN => n_4334);
   clk_r_REG3304_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1368, QN => n_4335);
   clk_r_REG3305_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1367, QN => n_4336);
   clk_r_REG3306_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1366, QN => n_4337);
   clk_r_REG3307_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_25_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1365, QN => n_4338);
   clk_r_REG3308_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_26_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1364, QN => n_4339);
   clk_r_REG3310_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1363, QN => n_4340);
   clk_r_REG3311_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_27_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1362, QN => n_4341);
   clk_r_REG3312_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_28_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1361, QN => n_4342);
   clk_r_REG3313_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_29_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1360, QN => n_4343);
   clk_r_REG3314_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_30_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1359, QN => n_4344);
   clk_r_REG3315_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => n1358, QN => n_4345);
   clk_r_REG3316_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1357, QN => n_4346);
   clk_r_REG3317_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1356, QN => n_4347);
   clk_r_REG3318_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1355, QN => n_4348);
   clk_r_REG3319_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1354, QN => n_4349);
   clk_r_REG3320_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1353, QN => n_4350);
   clk_r_REG3321_S2 : DFFR_X1 port map( D => datapath_i_val_immediate_i_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => n1352, QN => n_4351);
   clk_r_REG3474_S7 : DFFR_X1 port map( D => n2294, CK => CLK, RN => RST, Q => 
                           n_4352, QN => n1351);
   clk_r_REG3479_S7 : DFFR_X1 port map( D => n468, CK => CLK, RN => RST, Q => 
                           n1350, QN => n_4353);
   clk_r_REG3470_S7 : DFFS_X1 port map( D => n485, CK => CLK, SN => RST, Q => 
                           n1349, QN => n_4354);
   clk_r_REG3252_S2 : DFFR_X1 port map( D => n2251, CK => CLK, RN => RST, Q => 
                           n_4355, QN => n1348);
   clk_r_REG3325_S2 : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK => CLK, 
                           RN => RST, Q => n1347, QN => n_4356);
   clk_r_REG739_S6 : DFFR_X1 port map( D => n377, CK => CLK, RN => RST, Q => 
                           n1346, QN => n_4357);
   clk_r_REG471_S6 : DFFR_X1 port map( D => n380, CK => CLK, RN => RST, Q => 
                           n1345, QN => n_4358);
   clk_r_REG822_S22 : DFFR_X1 port map( D => n385, CK => CLK, RN => RST, Q => 
                           n1344, QN => n_4359);
   clk_r_REG1073_S18 : DFFR_X1 port map( D => n390, CK => CLK, RN => RST, Q => 
                           n1343, QN => n_4360);
   clk_r_REG332_S6 : DFFR_X1 port map( D => n395, CK => CLK, RN => RST, Q => 
                           n1342, QN => n_4361);
   clk_r_REG1633_S6 : DFFR_X1 port map( D => n400, CK => CLK, RN => RST, Q => 
                           n1341, QN => n_4362);
   clk_r_REG148_S34 : DFFR_X1 port map( D => n405, CK => CLK, RN => RST, Q => 
                           n1340, QN => n_4363);
   clk_r_REG2103_S37 : DFFR_X1 port map( D => n415, CK => CLK, RN => RST, Q => 
                           n1339, QN => n_4364);
   clk_r_REG1942_S40 : DFFR_X1 port map( D => n420, CK => CLK, RN => RST, Q => 
                           n1338, QN => n_4365);
   clk_r_REG1867_S41 : DFFR_X1 port map( D => n426, CK => CLK, RN => RST, Q => 
                           n1337, QN => n_4366);
   clk_r_REG2104_S44 : DFFR_X1 port map( D => n431, CK => CLK, RN => RST, Q => 
                           n1336, QN => n_4367);
   clk_r_REG2105_S47 : DFFR_X1 port map( D => n436, CK => CLK, RN => RST, Q => 
                           n1335, QN => n_4368);
   clk_r_REG2106_S50 : DFFR_X1 port map( D => n441, CK => CLK, RN => RST, Q => 
                           n1334, QN => n_4369);
   clk_r_REG3327_S1 : DFFS_X1 port map( D => n676, CK => CLK, SN => RST, Q => 
                           n1333, QN => n_4370);
   clk_r_REG3248_S2 : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK => CLK, 
                           RN => RST, Q => n1332, QN => n_4371);
   clk_r_REG3180_S1 : DFFS_X1 port map( D => cu_i_n153, CK => CLK, SN => RST, Q
                           => n1331, QN => n2553);
   clk_r_REG1465_S9 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_2_port, CK => CLK, RN
                           => RST, Q => n1330, QN => n_4372);
   clk_r_REG1483_S10 : DFFR_X1 port map( D => n1330, CK => CLK, RN => RST, Q =>
                           n_4373, QN => n1868);
   clk_r_REG318_S9 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_3_port, CK => CLK, RN
                           => RST, Q => n1328, QN => n_4374);
   clk_r_REG319_S10 : DFFR_X1 port map( D => n1328, CK => CLK, RN => RST, Q => 
                           n_4375, QN => n1867);
   clk_r_REG321_S9 : DFFS_X1 port map( D => n524, CK => CLK, SN => RST, Q => 
                           n1326, QN => n_4376);
   clk_r_REG903_S6 : DFFS_X1 port map( D => n523, CK => CLK, SN => RST, Q => 
                           n1325, QN => n_4377);
   clk_r_REG373_S6 : DFFS_X1 port map( D => n529, CK => CLK, SN => RST, Q => 
                           n1324, QN => n_4378);
   clk_r_REG137_S6 : DFFS_X1 port map( D => n535, CK => CLK, SN => RST, Q => 
                           n1323, QN => n_4379);
   clk_r_REG30_S22 : DFFS_X1 port map( D => n541, CK => CLK, SN => RST, Q => 
                           n1322, QN => n_4380);
   clk_r_REG178_S6 : DFFS_X1 port map( D => n547, CK => CLK, SN => RST, Q => 
                           n1321, QN => n_4381);
   clk_r_REG239_S6 : DFFS_X1 port map( D => n553, CK => CLK, SN => RST, Q => 
                           n1320, QN => n_4382);
   clk_r_REG41_S31 : DFFS_X1 port map( D => n559, CK => CLK, SN => RST, Q => 
                           n1319, QN => n_4383);
   clk_r_REG49_S34 : DFFS_X1 port map( D => n565, CK => CLK, SN => RST, Q => 
                           n1318, QN => n_4384);
   clk_r_REG60_S37 : DFFS_X1 port map( D => n571, CK => CLK, SN => RST, Q => 
                           n1317, QN => n_4385);
   clk_r_REG159_S40 : DFFS_X1 port map( D => n577, CK => CLK, SN => RST, Q => 
                           n1316, QN => n_4386);
   clk_r_REG74_S41 : DFFS_X1 port map( D => n583, CK => CLK, SN => RST, Q => 
                           n1315, QN => n_4387);
   clk_r_REG84_S44 : DFFS_X1 port map( D => n589, CK => CLK, SN => RST, Q => 
                           n1314, QN => n_4388);
   clk_r_REG99_S47 : DFFS_X1 port map( D => n595, CK => CLK, SN => RST, Q => 
                           n1313, QN => n_4389);
   clk_r_REG110_S50 : DFFS_X1 port map( D => n601, CK => CLK, SN => RST, Q => 
                           n1312, QN => n_4390);
   clk_r_REG116_S52 : DFFR_X1 port map( D => 
                           datapath_i_new_pc_value_decode_31_port, CK => CLK, 
                           RN => RST, Q => n_4391, QN => n1844);
   clk_r_REG130_S3 : DFFR_X1 port map( D => n717, CK => CLK, RN => RST, Q => 
                           n1310, QN => n1866);
   clk_r_REG12_S11 : DFFS_X1 port map( D => n692, CK => CLK, SN => RST, Q => 
                           n1308, QN => n_4392);
   clk_r_REG19_S13 : DFFS_X1 port map( D => n699, CK => CLK, SN => RST, Q => 
                           n1307, QN => n_4393);
   clk_r_REG1466_S9 : DFFS_X1 port map( D => n700, CK => CLK, SN => RST, Q => 
                           n1306, QN => n_4394);
   clk_r_REG3478_S7 : DFFS_X1 port map( D => n464, CK => CLK, SN => RST, Q => 
                           n1305, QN => n_4395);
   clk_r_REG3264_S1 : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           CK => CLK, RN => RST, Q => n1304, QN => n_4396);
   clk_r_REG3265_S2 : DFFR_X1 port map( D => n1304, CK => CLK, RN => RST, Q => 
                           n1303, QN => n_4397);
   clk_r_REG3266_S3 : DFFR_X1 port map( D => n1303, CK => CLK, RN => RST, Q => 
                           n1302, QN => n_4398);
   clk_r_REG3322_S1 : DFFR_X1 port map( D => n302, CK => CLK, RN => RST, Q => 
                           n1301, QN => n_4399);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => n1770, ADD_WR(3) => n1767, ADD_WR(2) =>
                           n1302, ADD_WR(1) => n1761, ADD_WR(0) => n1764, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n43, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n44, OUT1(31) => 
                           datapath_i_val_a_i_31_port, OUT1(30) => 
                           datapath_i_val_a_i_30_port, OUT1(29) => 
                           datapath_i_val_a_i_29_port, OUT1(28) => 
                           datapath_i_val_a_i_28_port, OUT1(27) => 
                           datapath_i_val_a_i_27_port, OUT1(26) => 
                           datapath_i_val_a_i_26_port, OUT1(25) => 
                           datapath_i_val_a_i_25_port, OUT1(24) => 
                           datapath_i_val_a_i_24_port, OUT1(23) => 
                           datapath_i_val_a_i_23_port, OUT1(22) => 
                           datapath_i_val_a_i_22_port, OUT1(21) => 
                           datapath_i_val_a_i_21_port, OUT1(20) => 
                           datapath_i_val_a_i_20_port, OUT1(19) => 
                           datapath_i_val_a_i_19_port, OUT1(18) => 
                           datapath_i_val_a_i_18_port, OUT1(17) => 
                           datapath_i_val_a_i_17_port, OUT1(16) => 
                           datapath_i_val_a_i_16_port, OUT1(15) => 
                           datapath_i_val_a_i_15_port, OUT1(14) => 
                           datapath_i_val_a_i_14_port, OUT1(13) => 
                           datapath_i_val_a_i_13_port, OUT1(12) => 
                           datapath_i_val_a_i_12_port, OUT1(11) => 
                           datapath_i_val_a_i_11_port, OUT1(10) => 
                           datapath_i_val_a_i_10_port, OUT1(9) => 
                           datapath_i_val_a_i_9_port, OUT1(8) => 
                           datapath_i_val_a_i_8_port, OUT1(7) => 
                           datapath_i_val_a_i_7_port, OUT1(6) => 
                           datapath_i_val_a_i_6_port, OUT1(5) => 
                           datapath_i_val_a_i_5_port, OUT1(4) => 
                           datapath_i_val_a_i_4_port, OUT1(3) => 
                           datapath_i_val_a_i_3_port, OUT1(2) => 
                           datapath_i_val_a_i_2_port, OUT1(1) => 
                           datapath_i_val_a_i_1_port, OUT1(0) => 
                           datapath_i_val_a_i_0_port, OUT2(31) => 
                           datapath_i_val_b_i_31_port, OUT2(30) => 
                           datapath_i_val_b_i_30_port, OUT2(29) => 
                           datapath_i_val_b_i_29_port, OUT2(28) => 
                           datapath_i_val_b_i_28_port, OUT2(27) => 
                           datapath_i_val_b_i_27_port, OUT2(26) => 
                           datapath_i_val_b_i_26_port, OUT2(25) => 
                           datapath_i_val_b_i_25_port, OUT2(24) => 
                           datapath_i_val_b_i_24_port, OUT2(23) => 
                           datapath_i_val_b_i_23_port, OUT2(22) => 
                           datapath_i_val_b_i_22_port, OUT2(21) => 
                           datapath_i_val_b_i_21_port, OUT2(20) => 
                           datapath_i_val_b_i_20_port, OUT2(19) => 
                           datapath_i_val_b_i_19_port, OUT2(18) => 
                           datapath_i_val_b_i_18_port, OUT2(17) => 
                           datapath_i_val_b_i_17_port, OUT2(16) => 
                           datapath_i_val_b_i_16_port, OUT2(15) => 
                           datapath_i_val_b_i_15_port, OUT2(14) => 
                           datapath_i_val_b_i_14_port, OUT2(13) => 
                           datapath_i_val_b_i_13_port, OUT2(12) => 
                           datapath_i_val_b_i_12_port, OUT2(11) => 
                           datapath_i_val_b_i_11_port, OUT2(10) => 
                           datapath_i_val_b_i_10_port, OUT2(9) => 
                           datapath_i_val_b_i_9_port, OUT2(8) => 
                           datapath_i_val_b_i_8_port, OUT2(7) => 
                           datapath_i_val_b_i_7_port, OUT2(6) => 
                           datapath_i_val_b_i_6_port, OUT2(5) => 
                           datapath_i_val_b_i_5_port, OUT2(4) => 
                           datapath_i_val_b_i_4_port, OUT2(3) => 
                           datapath_i_val_b_i_3_port, OUT2(2) => 
                           datapath_i_val_b_i_2_port, OUT2(1) => 
                           datapath_i_val_b_i_1_port, OUT2(0) => 
                           datapath_i_val_b_i_0_port, RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_4400, mul_exeception => 
                           n_4401, FUNC(0) => n2245, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_4402, 
                           OUTALU(31) => datapath_i_alu_output_val_i_31_port, 
                           OUTALU(30) => datapath_i_alu_output_val_i_30_port, 
                           OUTALU(29) => datapath_i_alu_output_val_i_29_port, 
                           OUTALU(28) => datapath_i_alu_output_val_i_28_port, 
                           OUTALU(27) => datapath_i_alu_output_val_i_27_port, 
                           OUTALU(26) => datapath_i_alu_output_val_i_26_port, 
                           OUTALU(25) => datapath_i_alu_output_val_i_25_port, 
                           OUTALU(24) => datapath_i_alu_output_val_i_24_port, 
                           OUTALU(23) => datapath_i_alu_output_val_i_23_port, 
                           OUTALU(22) => datapath_i_alu_output_val_i_22_port, 
                           OUTALU(21) => datapath_i_alu_output_val_i_21_port, 
                           OUTALU(20) => datapath_i_alu_output_val_i_20_port, 
                           OUTALU(19) => datapath_i_alu_output_val_i_19_port, 
                           OUTALU(18) => datapath_i_alu_output_val_i_18_port, 
                           OUTALU(17) => datapath_i_alu_output_val_i_17_port, 
                           OUTALU(16) => datapath_i_alu_output_val_i_16_port, 
                           OUTALU(15) => datapath_i_alu_output_val_i_15_port, 
                           OUTALU(14) => datapath_i_alu_output_val_i_14_port, 
                           OUTALU(13) => datapath_i_alu_output_val_i_13_port, 
                           OUTALU(12) => datapath_i_alu_output_val_i_12_port, 
                           OUTALU(11) => datapath_i_alu_output_val_i_11_port, 
                           OUTALU(10) => datapath_i_alu_output_val_i_10_port, 
                           OUTALU(9) => datapath_i_alu_output_val_i_9_port, 
                           OUTALU(8) => datapath_i_alu_output_val_i_8_port, 
                           OUTALU(7) => datapath_i_alu_output_val_i_7_port, 
                           OUTALU(6) => datapath_i_alu_output_val_i_6_port, 
                           OUTALU(5) => datapath_i_alu_output_val_i_5_port, 
                           OUTALU(4) => datapath_i_alu_output_val_i_4_port, 
                           OUTALU(3) => datapath_i_alu_output_val_i_3_port, 
                           OUTALU(2) => datapath_i_alu_output_val_i_2_port, 
                           OUTALU(1) => datapath_i_alu_output_val_i_1_port, 
                           OUTALU(0) => datapath_i_alu_output_val_i_0_port, 
                           rst_BAR => RST);
   U934 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_31_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(31), ZN => n2042
                           );
   U936 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_30_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(30), ZN => n2043
                           );
   U938 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_29_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(29), ZN => n2044
                           );
   U940 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_28_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(28), ZN => n2045
                           );
   U942 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_27_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(27), ZN => n2046
                           );
   U944 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_26_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(26), ZN => n2047
                           );
   U946 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_25_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(25), ZN => n2048
                           );
   U948 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_24_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(24), ZN => n2049
                           );
   U950 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_23_port, A2 => 
                           n2576, B1 => n2577, B2 => DRAM_DATA(23), ZN => n2050
                           );
   U952 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_22_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(22), ZN => n2051
                           );
   U954 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_21_port, A2 => 
                           n2576, B1 => n2073, B2 => DRAM_DATA(21), ZN => n2052
                           );
   U956 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_20_port, A2 => 
                           n2576, B1 => n2073, B2 => DRAM_DATA(20), ZN => n2053
                           );
   U958 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_19_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(19), ZN => n2054
                           );
   U960 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_18_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(18), ZN => n2055
                           );
   U962 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_17_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(17), ZN => n2056
                           );
   U964 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_16_port, A2 => 
                           n2576, B1 => n2073, B2 => DRAM_DATA(16), ZN => n2057
                           );
   U966 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_15_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(15), ZN => n2058
                           );
   U968 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_14_port, A2 => 
                           n2576, B1 => n2073, B2 => DRAM_DATA(14), ZN => n2059
                           );
   U970 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_13_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(13), ZN => n2060
                           );
   U972 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(12), B1 => n2074, B2 
                           => datapath_i_alu_output_val_i_12_port, ZN => n2061)
                           ;
   U974 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(11), B1 => n2074, B2 
                           => datapath_i_alu_output_val_i_11_port, ZN => n2062)
                           ;
   U976 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(10), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_10_port, ZN => n2063)
                           ;
   U978 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(9), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_9_port, ZN => n2064);
   U980 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(8), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_8_port, ZN => n2065);
   U982 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(7), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_7_port, ZN => n2066);
   U984 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(6), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_6_port, ZN => n2067);
   U986 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(5), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_5_port, ZN => n2068);
   U988 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(4), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_4_port, ZN => n2069);
   U990 : AOI22_X1 port map( A1 => n2073, A2 => DRAM_DATA(3), B1 => n2576, B2 
                           => datapath_i_alu_output_val_i_3_port, ZN => n2070);
   U992 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_2_port, A2 => 
                           n2576, B1 => n2073, B2 => DRAM_DATA(2), ZN => n2071)
                           ;
   U994 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_1_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(1), ZN => n2072)
                           ;
   U996 : AOI22_X1 port map( A1 => datapath_i_alu_output_val_i_0_port, A2 => 
                           n2074, B1 => n2073, B2 => DRAM_DATA(0), ZN => n2075)
                           ;
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   clk_r_REG3256_S2 : DFFS_X1 port map( D => datapath_i_memory_stage_dp_n2, CK 
                           => CLK, SN => RST, Q => n1807, QN => n_4403);
   clk_r_REG2102_S5 : DFFR_X1 port map( D => n1804, CK => CLK, RN => RST, Q => 
                           n1803, QN => n_4404);
   clk_r_REG128_S2 : DFF_X1 port map( D => datapath_i_val_a_i_31_port, CK => 
                           CLK, Q => n1673, QN => n_4405);
   clk_r_REG3336_S6 : DFFR_X1 port map( D => n719, CK => CLK, RN => RST, Q => 
                           n1801, QN => n2554);
   clk_r_REG3269_S1 : DFFS_X1 port map( D => n2256, CK => CLK, SN => RST, Q => 
                           n1802, QN => n_4406);
   clk_r_REG3272_S1 : DFFS_X1 port map( D => n705, CK => CLK, SN => RST, Q => 
                           n1507, QN => n_4407);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => n1458, Q => n719
                           );
   clk_r_REG3452_S7 : DFFR_X1 port map( D => curr_instruction_to_cu_i_15_port, 
                           CK => CLK, RN => RST, Q => n1405, QN => n_4408);
   clk_r_REG2097_S4 : DFFS_X1 port map( D => n375, CK => CLK, SN => RST, Q => 
                           n_4409, QN => n1804);
   clk_r_REG131_S4 : DFFS_X1 port map( D => n1866, CK => CLK, SN => RST, Q => 
                           n_4410, QN => n1309);
   clk_r_REG3271_S1 : DFFR_X1 port map( D => n703, CK => CLK, RN => RST, Q => 
                           n1727, QN => n_4411);
   clk_r_REG3334_S6 : DFFS_X1 port map( D => n2255, CK => CLK, SN => RST, Q => 
                           n2552, QN => n1509);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X2 port map( A => 
                           n1541, EN => n2574, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X2 port map( A => 
                           n1547, EN => n1807, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X2 port map( A => 
                           n1526, EN => n1497, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X2 port map( A => 
                           n1553, EN => n1807, Z => DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X2 port map( A => 
                           n1550, EN => n2574, Z => DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X2 port map( A => 
                           n1544, EN => n2574, Z => DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X2 port map( A => 
                           n1538, EN => n1497, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X2 port map( A => 
                           n1535, EN => n1497, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X2 port map( A => 
                           n1532, EN => n1497, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X2 port map( A => 
                           n1529, EN => n1497, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X2 port map( A => 
                           n1607, EN => n2574, Z => DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X2 port map( A => 
                           n1601, EN => n2574, Z => DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X2 port map( A => 
                           n1595, EN => n2574, Z => DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X2 port map( A => 
                           n1589, EN => n2574, Z => DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X2 port map( A => 
                           n1583, EN => n2574, Z => DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X2 port map( A => 
                           n1562, EN => n2574, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X2 port map( A => 
                           n1556, EN => n2574, Z => DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X2 port map( A => 
                           n1610, EN => n1807, Z => DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X2 port map( A => 
                           n1604, EN => n1807, Z => DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X2 port map( A => 
                           n1598, EN => n1807, Z => DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X2 port map( A => 
                           n1592, EN => n1807, Z => DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X2 port map( A => 
                           n1586, EN => n1807, Z => DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X2 port map( A => 
                           n1580, EN => n1807, Z => DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X2 port map( A => 
                           n1559, EN => n1807, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X2 port map( A => 
                           n1517, EN => n2574, Z => DRAM_DATA(0));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X2 port map( A => 
                           n1577, EN => n1497, Z => DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X2 port map( A => 
                           n1574, EN => n1497, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X2 port map( A => 
                           n1571, EN => n1497, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X2 port map( A => 
                           n1568, EN => n1497, Z => DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X2 port map( A => 
                           n1565, EN => n1497, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X2 port map( A => 
                           n1523, EN => n1497, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X2 port map( A => 
                           n1520, EN => n1497, Z => DRAM_DATA(1));
   U1255 : OAI21_X2 port map( B1 => n2544, B2 => n1685, A => n2365, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U1256 : OAI21_X2 port map( B1 => n1507, B2 => n1689, A => n2371, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U1257 : INV_X2 port map( A => n2336, ZN => n2513);
   U1258 : BUF_X1 port map( A => n1916, Z => IRAM_ADDRESS_31_port);
   U1259 : AOI22_X1 port map( A1 => n1801, A2 => cu_i_cmd_alu_op_type_3_port, 
                           B1 => n1674, B2 => n1514, ZN => n2514);
   U1260 : AOI22_X1 port map( A1 => n1801, A2 => cu_i_cmd_alu_op_type_1_port, 
                           B1 => n1674, B2 => n1516, ZN => n2518);
   U1261 : NOR2_X1 port map( A1 => n2515, A2 => n2338, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U1262 : NOR2_X1 port map( A1 => n2516, A2 => n2340, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U1263 : NOR2_X1 port map( A1 => n1475, A2 => n2553, ZN => n2461);
   U1264 : MUX2_X1 port map( A => n1355, B => n1527, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U1265 : MUX2_X1 port map( A => n1363, B => n1518, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U1266 : INV_X1 port map( A => n719, ZN => n2255);
   U1267 : OAI22_X1 port map( A1 => n2255, A2 => n1778, B1 => n1422, B2 => n719
                           , ZN => n2305);
   U1268 : INV_X1 port map( A => n2305, ZN => n2253);
   U1269 : AOI22_X1 port map( A1 => n1801, A2 => n1408, B1 => IRAM_DATA(18), B2
                           => n2554, ZN => n2258);
   U1270 : INV_X1 port map( A => n2258, ZN => curr_instruction_to_cu_i_18_port)
                           ;
   U1271 : AOI22_X1 port map( A1 => n1509, A2 => n1419, B1 => IRAM_DATA(29), B2
                           => n2552, ZN => n2300);
   U1272 : AOI22_X1 port map( A1 => n1509, A2 => n1416, B1 => IRAM_DATA(26), B2
                           => n2552, ZN => n2295);
   U1273 : AOI22_X1 port map( A1 => n1509, A2 => n1421, B1 => IRAM_DATA(31), B2
                           => n2552, ZN => n2302);
   U1274 : AOI22_X1 port map( A1 => n1509, A2 => n1420, B1 => IRAM_DATA(30), B2
                           => n2552, ZN => n2301);
   U1275 : AOI22_X1 port map( A1 => n1509, A2 => n1418, B1 => IRAM_DATA(28), B2
                           => n2552, ZN => n2298);
   U1276 : AOI22_X1 port map( A1 => n1509, A2 => n1417, B1 => IRAM_DATA(27), B2
                           => n2552, ZN => n2296);
   U1277 : INV_X1 port map( A => n2300, ZN => n2310);
   U1278 : INV_X1 port map( A => n2296, ZN => n2315);
   U1279 : NAND3_X1 port map( A1 => n2301, A2 => n2298, A3 => n2315, ZN => 
                           n2465);
   U1280 : NOR3_X1 port map( A1 => n2295, A2 => n2302, A3 => n2465, ZN => n2329
                           );
   U1281 : NAND2_X1 port map( A1 => n2461, A2 => n2329, ZN => n2509);
   U1282 : NOR2_X1 port map( A1 => n2310, A2 => n2509, ZN => 
                           cu_i_cmd_word_3_port);
   U1283 : OAI22_X1 port map( A1 => n2255, A2 => cu_i_cmd_word_3_port, B1 => 
                           n1425, B2 => n719, ZN => n2407);
   U1284 : INV_X1 port map( A => n2407, ZN => n2252);
   U1285 : INV_X1 port map( A => n2509, ZN => cu_i_cmd_word_4_port);
   U1286 : OAI22_X1 port map( A1 => n2255, A2 => cu_i_cmd_word_4_port, B1 => 
                           n1424, B2 => n719, ZN => n361);
   U1287 : INV_X1 port map( A => n361, ZN => n2251);
   U1288 : INV_X1 port map( A => n2295, ZN => n2307);
   U1289 : NOR2_X1 port map( A1 => n2307, A2 => n2315, ZN => n2292);
   U1290 : INV_X1 port map( A => n2292, ZN => n2327);
   U1291 : INV_X1 port map( A => n2301, ZN => n2313);
   U1292 : INV_X1 port map( A => n2302, ZN => n2308);
   U1293 : NOR3_X1 port map( A1 => n2298, A2 => n2313, A3 => n2308, ZN => n2326
                           );
   U1294 : NAND3_X1 port map( A1 => n2300, A2 => n2461, A3 => n2326, ZN => 
                           n2306);
   U1295 : NAND2_X1 port map( A1 => n2300, A2 => n2302, ZN => n2311);
   U1296 : NOR2_X1 port map( A1 => n2311, A2 => n2465, ZN => n2330);
   U1297 : NAND2_X1 port map( A1 => n2461, A2 => n2330, ZN => n2510);
   U1298 : OAI21_X1 port map( B1 => n2327, B2 => n2306, A => n2510, ZN => 
                           cu_i_cmd_word_6_port);
   U1299 : NAND2_X1 port map( A1 => n2296, A2 => n2307, ZN => n474);
   U1300 : NOR2_X1 port map( A1 => n474, A2 => n2306, ZN => 
                           cu_i_cmd_word_7_port);
   U1301 : OR2_X1 port map( A1 => cu_i_cmd_word_6_port, A2 => 
                           cu_i_cmd_word_7_port, ZN => cu_i_n135);
   U1302 : AOI22_X1 port map( A1 => n719, A2 => cu_i_n135, B1 => n1496, B2 => 
                           n2255, ZN => n2256);
   U1303 : NOR4_X1 port map( A1 => n2298, A2 => n2301, A3 => n2307, A4 => n2311
                           , ZN => n468);
   U1304 : NOR2_X1 port map( A1 => n2308, A2 => n2300, ZN => n2460);
   U1305 : AND2_X1 port map( A1 => n2313, A2 => n2460, ZN => n475);
   U1306 : INV_X1 port map( A => n2298, ZN => n2312);
   U1307 : OAI211_X1 port map( C1 => n2307, C2 => n2312, A => n2296, B => n475,
                           ZN => n485);
   U1308 : NAND2_X1 port map( A1 => n2326, A2 => n2310, ZN => n2299);
   U1309 : AOI211_X1 port map( C1 => n2296, C2 => n2298, A => n2313, B => n2308
                           , ZN => n2309);
   U1310 : NAND3_X1 port map( A1 => n2295, A2 => n2310, A3 => n2309, ZN => n464
                           );
   U1311 : NOR4_X1 port map( A1 => n2313, A2 => n2312, A3 => n2311, A4 => n2327
                           , ZN => n2413);
   U1312 : NAND2_X1 port map( A1 => n2461, A2 => n2413, ZN => n2293);
   U1313 : AOI22_X1 port map( A1 => n1509, A2 => n1392, B1 => IRAM_DATA(2), B2 
                           => n2552, ZN => n2290);
   U1314 : AOI22_X1 port map( A1 => n1509, A2 => n1391, B1 => IRAM_DATA(1), B2 
                           => n2552, ZN => n2289);
   U1315 : MUX2_X1 port map( A => IRAM_DATA(4), B => n1394, S => n1509, Z => 
                           curr_instruction_to_cu_i_4_port);
   U1316 : MUX2_X1 port map( A => IRAM_DATA(0), B => n1390, S => n1509, Z => 
                           curr_instruction_to_cu_i_0_port);
   U1317 : AOI22_X1 port map( A1 => n1509, A2 => n1395, B1 => IRAM_DATA(5), B2 
                           => n2552, ZN => n2291);
   U1318 : MUX2_X1 port map( A => IRAM_DATA(3), B => n1393, S => n1509, Z => 
                           curr_instruction_to_cu_i_3_port);
   U1319 : INV_X1 port map( A => n2461, ZN => n2474);
   U1320 : INV_X1 port map( A => n485, ZN => n2317);
   U1321 : NAND3_X1 port map( A1 => n2301, A2 => n2292, A3 => n2460, ZN => 
                           n2314);
   U1322 : OAI211_X1 port map( C1 => n2315, C2 => n2299, A => n2314, B => n464,
                           ZN => n2316);
   U1323 : NOR3_X1 port map( A1 => n468, A2 => n2317, A3 => n2316, ZN => n2468)
                           ;
   U1324 : INV_X1 port map( A => n2291, ZN => n2462);
   U1325 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => 
                           curr_instruction_to_cu_i_0_port, A3 => n2462, A4 => 
                           curr_instruction_to_cu_i_3_port, ZN => n2318);
   U1326 : NOR3_X1 port map( A1 => n2290, A2 => n2289, A3 => n2318, ZN => n2412
                           );
   U1327 : OAI222_X1 port map( A1 => n2474, A2 => n2468, B1 => n2510, B2 => 
                           n2295, C1 => n2293, C2 => n2412, ZN => n302);
   U1328 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n302, ZN => 
                           cu_i_cw1_5_port);
   U1329 : INV_X1 port map( A => n2413, ZN => n2294);
   U1330 : NOR2_X1 port map( A1 => cu_i_n2, A2 => cu_i_n4, ZN => n2320);
   U1331 : NAND3_X1 port map( A1 => cu_i_n152, A2 => cu_i_n151, A3 => n2320, ZN
                           => cu_i_n145);
   U1332 : INV_X1 port map( A => cu_i_n151, ZN => n2319);
   U1333 : NOR2_X1 port map( A1 => n2320, A2 => n2319, ZN => n2246);
   U1334 : MUX2_X1 port map( A => IRAM_DATA(19), B => n1409, S => n1801, Z => 
                           curr_instruction_to_cu_i_19_port);
   U1335 : MUX2_X1 port map( A => IRAM_DATA(14), B => n1404, S => n1801, Z => 
                           curr_instruction_to_cu_i_14_port);
   U1336 : INV_X1 port map( A => n2510, ZN => n2297);
   U1337 : CLKBUF_X1 port map( A => n2297, Z => n2575);
   U1338 : INV_X1 port map( A => n2246, ZN => n2321);
   U1339 : NAND2_X1 port map( A1 => cu_i_n145, A2 => n2321, ZN => n2414);
   U1340 : AOI21_X1 port map( B1 => n2412, B2 => n2414, A => n2293, ZN => n2512
                           );
   U1341 : INV_X1 port map( A => n2512, ZN => n2511);
   U1342 : AOI221_X1 port map( B1 => n2511, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n2512, C2 =>
                           curr_instruction_to_cu_i_14_port, A => n2575, ZN => 
                           n2322);
   U1343 : INV_X1 port map( A => n2322, ZN => n2249);
   U1344 : MUX2_X1 port map( A => IRAM_DATA(17), B => n1407, S => n1801, Z => 
                           curr_instruction_to_cu_i_17_port);
   U1345 : MUX2_X1 port map( A => IRAM_DATA(12), B => n1402, S => n1801, Z => 
                           curr_instruction_to_cu_i_12_port);
   U1346 : AOI221_X1 port map( B1 => n2511, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n2512, C2 =>
                           curr_instruction_to_cu_i_12_port, A => n2575, ZN => 
                           n2323);
   U1347 : INV_X1 port map( A => n2323, ZN => n2247);
   U1348 : MUX2_X1 port map( A => IRAM_DATA(20), B => n1410, S => n1801, Z => 
                           curr_instruction_to_cu_i_20_port);
   U1349 : MUX2_X1 port map( A => IRAM_DATA(15), B => n1405, S => n1801, Z => 
                           curr_instruction_to_cu_i_15_port);
   U1350 : AOI221_X1 port map( B1 => n2511, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n2512, C2 =>
                           curr_instruction_to_cu_i_15_port, A => n2575, ZN => 
                           n2324);
   U1351 : INV_X1 port map( A => n2324, ZN => n2250);
   U1352 : MUX2_X1 port map( A => IRAM_DATA(16), B => n1406, S => n1801, Z => 
                           curr_instruction_to_cu_i_16_port);
   U1353 : MUX2_X1 port map( A => IRAM_DATA(11), B => n1401, S => n1509, Z => 
                           curr_instruction_to_cu_i_11_port);
   U1354 : AOI221_X1 port map( B1 => n2511, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n2512, C2 =>
                           curr_instruction_to_cu_i_11_port, A => n2575, ZN => 
                           n2325);
   U1355 : INV_X1 port map( A => n2325, ZN => n2248);
   U1356 : INV_X1 port map( A => n2326, ZN => n2328);
   U1357 : OAI21_X1 port map( B1 => n2328, B2 => n2327, A => n2468, ZN => n2331
                           );
   U1358 : NOR3_X1 port map( A1 => n2330, A2 => n2329, A3 => n2331, ZN => n2472
                           );
   U1359 : INV_X1 port map( A => cu_i_cmd_word_7_port, ZN => n2332);
   U1360 : OAI21_X1 port map( B1 => n2472, B2 => n2474, A => n2332, ZN => n301)
                           ;
   U1361 : CLKBUF_X1 port map( A => n301, Z => n2578);
   U1362 : AOI211_X1 port map( C1 => n2461, C2 => n2331, A => 
                           cu_i_cmd_word_4_port, B => n2512, ZN => n2333);
   U1363 : NAND2_X1 port map( A1 => n2333, A2 => n2332, ZN => enable_rf_i);
   U1364 : INV_X1 port map( A => n2293, ZN => n2415);
   U1365 : AND2_X1 port map( A1 => n2415, A2 => n2412, ZN => n2288);
   U1366 : AND2_X1 port map( A1 => n2246, A2 => n2288, ZN => n2334);
   U1367 : OR2_X1 port map( A1 => n1778, A2 => n2334, ZN => write_rf_i);
   U1368 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U1369 : NOR2_X1 port map( A1 => n2334, A2 => n1779, ZN => n2337);
   U1370 : AND4_X1 port map( A1 => n1767, A2 => n1302, A3 => n1761, A4 => n1764
                           , ZN => n2335);
   U1371 : AND2_X1 port map( A1 => n1770, A2 => n2335, ZN => n2336);
   U1372 : AND3_X1 port map( A1 => n2337, A2 => DRAM_READY, A3 => n2513, ZN => 
                           n2073);
   U1373 : CLKBUF_X1 port map( A => n2073, Z => n2577);
   U1374 : NOR2_X1 port map( A1 => n2337, A2 => n2336, ZN => n2074);
   U1375 : CLKBUF_X1 port map( A => n2074, Z => n2576);
   U1376 : AOI22_X1 port map( A1 => n1801, A2 => cu_i_cmd_alu_op_type_0_port, 
                           B1 => n1674, B2 => n1508, ZN => n2515);
   U1377 : AOI22_X1 port map( A1 => n1801, A2 => cu_i_cmd_alu_op_type_2_port, 
                           B1 => n1674, B2 => n1515, ZN => n2516);
   U1378 : AOI21_X1 port map( B1 => n2516, B2 => n2518, A => n2514, ZN => n2338
                           );
   U1379 : INV_X1 port map( A => n2514, ZN => n2340);
   U1380 : OAI211_X1 port map( C1 => n2515, C2 => n2518, A => n2340, B => n2516
                           , ZN => n2339);
   U1381 : INV_X1 port map( A => n2339, ZN => n2245);
   U1382 : MUX2_X1 port map( A => n1354, B => n1530, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U1383 : MUX2_X1 port map( A => n1353, B => n1533, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U1384 : NAND2_X1 port map( A1 => n1453, A2 => n1494, ZN => n2399);
   U1385 : NOR2_X1 port map( A1 => n1756, A2 => n2399, ZN => n2359);
   U1386 : NAND2_X1 port map( A1 => n2359, A2 => n1449, ZN => n2358);
   U1387 : NOR2_X1 port map( A1 => n1751, A2 => n2358, ZN => n2363);
   U1388 : NAND2_X1 port map( A1 => n2363, A2 => n1447, ZN => n2362);
   U1389 : NOR2_X1 port map( A1 => n1749, A2 => n2362, ZN => n2395);
   U1390 : NAND2_X1 port map( A1 => n2395, A2 => n1445, ZN => n2394);
   U1391 : NOR2_X1 port map( A1 => n1747, A2 => n2394, ZN => n2369);
   U1392 : NAND2_X1 port map( A1 => n2369, A2 => n1443, ZN => n2368);
   U1393 : NOR2_X1 port map( A1 => n1743, A2 => n2368, ZN => n2391);
   U1394 : NAND2_X1 port map( A1 => n2391, A2 => n1441, ZN => n2390);
   U1395 : NOR2_X1 port map( A1 => n1741, A2 => n2390, ZN => n2403);
   U1396 : NAND2_X1 port map( A1 => n2403, A2 => n1439, ZN => n2402);
   U1397 : NOR2_X1 port map( A1 => n1739, A2 => n2402, ZN => n2375);
   U1398 : NAND2_X1 port map( A1 => n2375, A2 => n1437, ZN => n2374);
   U1399 : NOR2_X1 port map( A1 => n1737, A2 => n2374, ZN => n2426);
   U1400 : NAND2_X1 port map( A1 => n2426, A2 => n1435, ZN => n2425);
   U1401 : NOR2_X1 port map( A1 => n1735, A2 => n2425, ZN => n2383);
   U1402 : NAND2_X1 port map( A1 => n2383, A2 => n1433, ZN => n2382);
   U1403 : NOR2_X1 port map( A1 => n1733, A2 => n2382, ZN => n2379);
   U1404 : NAND2_X1 port map( A1 => n2379, A2 => n1431, ZN => n2378);
   U1405 : NOR2_X1 port map( A1 => n1731, A2 => n2378, ZN => n2355);
   U1406 : NAND2_X1 port map( A1 => n2355, A2 => n1429, ZN => n2354);
   U1407 : NOR2_X1 port map( A1 => n1729, A2 => n2354, ZN => n2435);
   U1408 : AOI211_X1 port map( C1 => n1730, C2 => n2354, A => n1745, B => n2435
                           , ZN => n2341);
   U1409 : OR2_X1 port map( A1 => n1334, A2 => n2341, ZN => 
                           datapath_i_new_pc_value_decode_29_port);
   U1410 : AOI211_X1 port map( C1 => n1750, C2 => n2362, A => n1753, B => n2395
                           , ZN => n2342);
   U1411 : OR2_X1 port map( A1 => n1343, A2 => n2342, ZN => 
                           datapath_i_new_pc_value_decode_11_port);
   U1412 : AOI211_X1 port map( C1 => n1748, C2 => n2394, A => n1745, B => n2369
                           , ZN => n2343);
   U1413 : OR2_X1 port map( A1 => n1342, A2 => n2343, ZN => 
                           datapath_i_new_pc_value_decode_13_port);
   U1414 : AOI211_X1 port map( C1 => n1738, C2 => n2374, A => n1745, B => n2426
                           , ZN => n2344);
   U1415 : OR2_X1 port map( A1 => n1338, A2 => n2344, ZN => 
                           datapath_i_new_pc_value_decode_21_port);
   U1416 : AOI211_X1 port map( C1 => n1740, C2 => n2402, A => n1745, B => n2375
                           , ZN => n2345);
   U1417 : OR2_X1 port map( A1 => n1339, A2 => n2345, ZN => 
                           datapath_i_new_pc_value_decode_19_port);
   U1418 : AOI211_X1 port map( C1 => n1742, C2 => n2390, A => n1745, B => n2403
                           , ZN => n2346);
   U1419 : OR2_X1 port map( A1 => n1340, A2 => n2346, ZN => 
                           datapath_i_new_pc_value_decode_17_port);
   U1420 : AOI211_X1 port map( C1 => n1736, C2 => n2425, A => n1745, B => n2383
                           , ZN => n2347);
   U1421 : OR2_X1 port map( A1 => n1337, A2 => n2347, ZN => 
                           datapath_i_new_pc_value_decode_23_port);
   U1422 : AOI211_X1 port map( C1 => n1752, C2 => n2358, A => n1753, B => n2363
                           , ZN => n2348);
   U1423 : OR2_X1 port map( A1 => n1344, A2 => n2348, ZN => 
                           datapath_i_new_pc_value_decode_9_port);
   U1424 : AOI211_X1 port map( C1 => n1451, C2 => n1755, A => n1494, B => n1753
                           , ZN => n2349);
   U1425 : OR2_X1 port map( A1 => n1345, A2 => n2349, ZN => 
                           datapath_i_new_pc_value_decode_5_port);
   U1426 : AOI211_X1 port map( C1 => n1757, C2 => n2399, A => n1753, B => n2359
                           , ZN => n2350);
   U1427 : OR2_X1 port map( A1 => n1346, A2 => n2350, ZN => 
                           datapath_i_new_pc_value_decode_7_port);
   U1428 : AOI211_X1 port map( C1 => n1744, C2 => n2368, A => n1753, B => n2391
                           , ZN => n2351);
   U1429 : OR2_X1 port map( A1 => n1341, A2 => n2351, ZN => 
                           datapath_i_new_pc_value_decode_15_port);
   U1430 : AOI211_X1 port map( C1 => n1734, C2 => n2382, A => n1745, B => n2379
                           , ZN => n2352);
   U1431 : OR2_X1 port map( A1 => n1336, A2 => n2352, ZN => 
                           datapath_i_new_pc_value_decode_25_port);
   U1432 : AOI211_X1 port map( C1 => n1732, C2 => n2378, A => n1745, B => n2355
                           , ZN => n2353);
   U1433 : OR2_X1 port map( A1 => n1335, A2 => n2353, ZN => 
                           datapath_i_new_pc_value_decode_27_port);
   U1434 : CLKBUF_X1 port map( A => n1807, Z => n2574);
   U1435 : OR2_X1 port map( A1 => n1781, A2 => n1504, ZN => cu_i_N278);
   U1436 : INV_X1 port map( A => n1854, ZN => IRAM_ADDRESS_2_port);
   U1437 : INV_X1 port map( A => n1855, ZN => IRAM_ADDRESS_3_port);
   U1438 : INV_X1 port map( A => n1847, ZN => IRAM_ADDRESS_4_port);
   U1439 : INV_X1 port map( A => n1862, ZN => IRAM_ADDRESS_6_port);
   U1440 : INV_X1 port map( A => n1848, ZN => IRAM_ADDRESS_8_port);
   U1441 : INV_X1 port map( A => n1860, ZN => IRAM_ADDRESS_10_port);
   U1442 : INV_X1 port map( A => n1859, ZN => IRAM_ADDRESS_12_port);
   U1443 : INV_X1 port map( A => n1850, ZN => IRAM_ADDRESS_14_port);
   U1444 : INV_X1 port map( A => n1856, ZN => IRAM_ADDRESS_16_port);
   U1445 : INV_X1 port map( A => n1849, ZN => IRAM_ADDRESS_18_port);
   U1446 : INV_X1 port map( A => n1857, ZN => IRAM_ADDRESS_20_port);
   U1447 : INV_X1 port map( A => n1858, ZN => IRAM_ADDRESS_22_port);
   U1448 : INV_X1 port map( A => n1861, ZN => IRAM_ADDRESS_24_port);
   U1449 : INV_X1 port map( A => n1853, ZN => IRAM_ADDRESS_26_port);
   U1450 : INV_X1 port map( A => n1851, ZN => IRAM_ADDRESS_28_port);
   U1451 : INV_X1 port map( A => n1852, ZN => IRAM_ADDRESS_30_port);
   U1452 : OAI211_X1 port map( C1 => n2355, C2 => n1429, A => n1803, B => n2354
                           , ZN => n2356);
   U1453 : NAND2_X1 port map( A1 => n1313, A2 => n2356, ZN => 
                           datapath_i_new_pc_value_decode_28_port);
   U1454 : CLKBUF_X1 port map( A => n1507, Z => n2544);
   U1455 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_28_port, B1 => n1802,
                           B2 => n1666, ZN => n2357);
   U1456 : OAI21_X1 port map( B1 => n2544, B2 => n1703, A => n2357, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U1457 : OAI211_X1 port map( C1 => n2359, C2 => n1449, A => n1803, B => n2358
                           , ZN => n2360);
   U1458 : NAND2_X1 port map( A1 => n1323, A2 => n2360, ZN => 
                           datapath_i_new_pc_value_decode_8_port);
   U1459 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_8_port, B1 => n1802, 
                           B2 => n1626, ZN => n2361);
   U1460 : OAI21_X1 port map( B1 => n1507, B2 => n1683, A => n2361, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U1461 : OAI211_X1 port map( C1 => n2363, C2 => n1447, A => n1803, B => n2362
                           , ZN => n2364);
   U1462 : NAND2_X1 port map( A1 => n1322, A2 => n2364, ZN => 
                           datapath_i_new_pc_value_decode_10_port);
   U1463 : CLKBUF_X1 port map( A => n1802, Z => n2541);
   U1464 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_10_port, B1 => n2541,
                           B2 => n1630, ZN => n2365);
   U1465 : OAI21_X1 port map( B1 => n2544, B2 => n1676, A => n1307, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U1466 : AOI22_X1 port map( A1 => n1802, A2 => n1620, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_5_port, ZN => n2366);
   U1467 : OAI21_X1 port map( B1 => n2544, B2 => n1680, A => n2366, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U1468 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_7_port, B1 => n1802, 
                           B2 => n1624, ZN => n2367);
   U1469 : OAI21_X1 port map( B1 => n2544, B2 => n1682, A => n2367, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U1470 : OAI211_X1 port map( C1 => n2369, C2 => n1443, A => n1803, B => n2368
                           , ZN => n2370);
   U1471 : NAND2_X1 port map( A1 => n1320, A2 => n2370, ZN => 
                           datapath_i_new_pc_value_decode_14_port);
   U1472 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_14_port, B1 => n2541,
                           B2 => n1638, ZN => n2371);
   U1473 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_15_port, B1 => n1802,
                           B2 => n1640, ZN => n2372);
   U1474 : OAI21_X1 port map( B1 => n2544, B2 => n1690, A => n2372, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U1475 : AOI22_X1 port map( A1 => n2541, A2 => n1648, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_19_port, ZN => n2373)
                           ;
   U1476 : OAI21_X1 port map( B1 => n2544, B2 => n1694, A => n2373, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U1477 : OAI211_X1 port map( C1 => n2375, C2 => n1437, A => n1803, B => n2374
                           , ZN => n2376);
   U1478 : NAND2_X1 port map( A1 => n1317, A2 => n2376, ZN => 
                           datapath_i_new_pc_value_decode_20_port);
   U1479 : AOI22_X1 port map( A1 => n1802, A2 => n1650, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_20_port, ZN => n2377)
                           ;
   U1480 : OAI21_X1 port map( B1 => n2544, B2 => n1695, A => n2377, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U1481 : OAI211_X1 port map( C1 => n2379, C2 => n1431, A => n1803, B => n2378
                           , ZN => n2380);
   U1482 : NAND2_X1 port map( A1 => n1314, A2 => n2380, ZN => 
                           datapath_i_new_pc_value_decode_26_port);
   U1483 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_26_port, B1 => n1802,
                           B2 => n1662, ZN => n2381);
   U1484 : OAI21_X1 port map( B1 => n2544, B2 => n1701, A => n2381, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U1485 : OAI211_X1 port map( C1 => n2383, C2 => n1433, A => n1803, B => n2382
                           , ZN => n2384);
   U1486 : NAND2_X1 port map( A1 => n1315, A2 => n2384, ZN => 
                           datapath_i_new_pc_value_decode_24_port);
   U1487 : AOI22_X1 port map( A1 => n2541, A2 => n1658, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_24_port, ZN => n2385)
                           ;
   U1488 : OAI21_X1 port map( B1 => n1507, B2 => n1699, A => n2385, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U1489 : MUX2_X1 port map( A => n1357, B => n1521, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U1490 : MUX2_X1 port map( A => n1356, B => n1524, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U1491 : OR2_X1 port map( A1 => n1485, A2 => n2571, ZN => n2387);
   U1492 : NAND2_X1 port map( A1 => n1513, A2 => n1510, ZN => n2459);
   U1493 : NOR2_X1 port map( A1 => n2551, A2 => n2459, ZN => n2458);
   U1494 : OAI221_X1 port map( B1 => n1511, B2 => n2458, C1 => n2571, C2 => 
                           n2459, A => n1726, ZN => n2386);
   U1495 : OAI21_X1 port map( B1 => n1512, B2 => n2387, A => n2386, ZN => 
                           cu_i_N277);
   U1496 : INV_X1 port map( A => n2256, ZN => n2388);
   U1497 : NAND2_X1 port map( A1 => n1773, A2 => n2388, ZN => n705);
   U1498 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_9_port, B1 => n1802, 
                           B2 => n1628, ZN => n2389);
   U1499 : OAI21_X1 port map( B1 => n1507, B2 => n1684, A => n2389, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U1500 : OAI211_X1 port map( C1 => n2391, C2 => n1441, A => n1803, B => n2390
                           , ZN => n2392);
   U1501 : NAND2_X1 port map( A1 => n1319, A2 => n2392, ZN => 
                           datapath_i_new_pc_value_decode_16_port);
   U1502 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_16_port, B1 => n2541,
                           B2 => n1642, ZN => n2393);
   U1503 : OAI21_X1 port map( B1 => n1507, B2 => n1691, A => n2393, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U1504 : OAI211_X1 port map( C1 => n2395, C2 => n1445, A => n1803, B => n2394
                           , ZN => n2396);
   U1505 : NAND2_X1 port map( A1 => n1321, A2 => n2396, ZN => 
                           datapath_i_new_pc_value_decode_12_port);
   U1506 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_12_port, B1 => n2541,
                           B2 => n1634, ZN => n2397);
   U1507 : OAI21_X1 port map( B1 => n1507, B2 => n1687, A => n2397, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U1508 : NAND2_X1 port map( A1 => n1325, A2 => n1326, ZN => 
                           datapath_i_new_pc_value_decode_4_port);
   U1509 : AOI22_X1 port map( A1 => n2541, A2 => n1618, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_4_port, ZN => n2398);
   U1510 : OAI21_X1 port map( B1 => n1507, B2 => n1679, A => n2398, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U1511 : OAI211_X1 port map( C1 => n1453, C2 => n1494, A => n1803, B => n2399
                           , ZN => n2400);
   U1512 : NAND2_X1 port map( A1 => n1324, A2 => n2400, ZN => 
                           datapath_i_new_pc_value_decode_6_port);
   U1513 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_6_port, B1 => n2541, 
                           B2 => n1622, ZN => n2401);
   U1514 : OAI21_X1 port map( B1 => n1507, B2 => n1681, A => n2401, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);
   U1515 : OAI211_X1 port map( C1 => n2403, C2 => n1439, A => n1803, B => n2402
                           , ZN => n2404);
   U1516 : NAND2_X1 port map( A1 => n1318, A2 => n2404, ZN => 
                           datapath_i_new_pc_value_decode_18_port);
   U1517 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_18_port, B1 => n1802,
                           B2 => n1646, ZN => n2405);
   U1518 : OAI21_X1 port map( B1 => n1507, B2 => n1693, A => n2405, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U1519 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_11_port, B1 => n1802,
                           B2 => n1632, ZN => n2406);
   U1520 : OAI21_X1 port map( B1 => n1507, B2 => n1686, A => n2406, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U1521 : NOR2_X1 port map( A1 => n1773, A2 => n1310, ZN => n423);
   U1522 : NAND2_X1 port map( A1 => n1773, A2 => n1866, ZN => n513);
   U1523 : NAND2_X1 port map( A1 => n2251, A2 => n2407, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U1524 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_6_port, B1 => n1759, 
                           B2 => datapath_i_alu_output_val_i_6_port, ZN => 
                           n2408);
   U1525 : OAI21_X1 port map( B1 => n1505, B2 => n1681, A => n2408, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U1526 : AOI222_X1 port map( A1 => n2557, A2 => n2549, B1 => n1759, B2 => 
                           datapath_i_alu_output_val_i_5_port, C1 => 
                           datapath_i_new_pc_value_decode_5_port, C2 => n1758, 
                           ZN => n2279);
   U1527 : AOI22_X1 port map( A1 => n1309, A2 => 
                           datapath_i_alu_output_val_i_2_port, B1 => n1506, B2 
                           => n1330, ZN => n2409);
   U1528 : OAI21_X1 port map( B1 => n1783, B2 => n1677, A => n2409, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U1529 : AOI22_X1 port map( A1 => n1309, A2 => 
                           datapath_i_alu_output_val_i_3_port, B1 => n1506, B2 
                           => n1328, ZN => n2410);
   U1530 : OAI21_X1 port map( B1 => n1783, B2 => n1678, A => n2410, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U1531 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_4_port, B1 => n1759, 
                           B2 => datapath_i_alu_output_val_i_4_port, ZN => 
                           n2411);
   U1532 : OAI21_X1 port map( B1 => n1783, B2 => n1679, A => n2411, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U1533 : NAND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_2_port,
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, ZN
                           => n2476);
   U1534 : INV_X1 port map( A => n2476, ZN => n2479);
   U1535 : NAND2_X1 port map( A1 => n2479, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, ZN => 
                           n519);
   U1536 : NOR2_X1 port map( A1 => n2279, A2 => n519, ZN => n526);
   U1537 : AOI221_X1 port map( B1 => n1426, B2 => n2255, C1 => cu_i_n135, C2 =>
                           n719, A => n1310, ZN => n375);
   U1538 : NAND2_X1 port map( A1 => n2413, A2 => n2412, ZN => n477);
   U1539 : AOI22_X1 port map( A1 => n2461, A2 => n477, B1 => n2415, B2 => n2414
                           , ZN => n2417);
   U1540 : NAND2_X1 port map( A1 => n1475, A2 => n2553, ZN => n2416);
   U1541 : AOI21_X1 port map( B1 => n2417, B2 => n2416, A => n719, ZN => n793);
   U1542 : NAND2_X1 port map( A1 => n793, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, ZN => 
                           n514);
   U1543 : NAND3_X1 port map( A1 => n1846, A2 => n1457, A3 => n1454, ZN => 
                           n2481);
   U1544 : NOR2_X1 port map( A1 => n1706, A2 => n2481, ZN => n2484);
   U1545 : NAND2_X1 port map( A1 => n1453, A2 => n2484, ZN => n2483);
   U1546 : NOR2_X1 port map( A1 => n1707, A2 => n2483, ZN => n2486);
   U1547 : AOI211_X1 port map( C1 => n1707, C2 => n2483, A => n2486, B => n1804
                           , ZN => n377);
   U1548 : AOI211_X1 port map( C1 => n1706, C2 => n2481, A => n2484, B => n1804
                           , ZN => n380);
   U1549 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_8_port, B1 => n1759, 
                           B2 => datapath_i_alu_output_val_i_8_port, ZN => 
                           n2418);
   U1550 : OAI21_X1 port map( B1 => n1505, B2 => n1683, A => n2418, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U1551 : NAND2_X1 port map( A1 => n1449, A2 => n2486, ZN => n2485);
   U1552 : NOR2_X1 port map( A1 => n1708, A2 => n2485, ZN => n2488);
   U1553 : AOI211_X1 port map( C1 => n1708, C2 => n2485, A => n2488, B => n1804
                           , ZN => n385);
   U1554 : AOI22_X1 port map( A1 => n1759, A2 => 
                           datapath_i_alu_output_val_i_10_port, B1 => n1506, B2
                           => datapath_i_new_pc_value_decode_10_port, ZN => 
                           n2419);
   U1555 : OAI21_X1 port map( B1 => n1505, B2 => n1685, A => n2419, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U1556 : NAND2_X1 port map( A1 => n1447, A2 => n2488, ZN => n2487);
   U1557 : NOR2_X1 port map( A1 => n1709, A2 => n2487, ZN => n2490);
   U1558 : AOI211_X1 port map( C1 => n1709, C2 => n2487, A => n2490, B => n1804
                           , ZN => n390);
   U1559 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_12_port, B1 => n1759,
                           B2 => datapath_i_alu_output_val_i_12_port, ZN => 
                           n2420);
   U1560 : OAI21_X1 port map( B1 => n1505, B2 => n1687, A => n2420, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U1561 : NAND2_X1 port map( A1 => n1445, A2 => n2490, ZN => n2489);
   U1562 : NOR2_X1 port map( A1 => n1710, A2 => n2489, ZN => n2492);
   U1563 : AOI211_X1 port map( C1 => n1710, C2 => n2489, A => n2492, B => n1804
                           , ZN => n395);
   U1564 : AOI22_X1 port map( A1 => n1309, A2 => 
                           datapath_i_alu_output_val_i_14_port, B1 => n1506, B2
                           => datapath_i_new_pc_value_decode_14_port, ZN => 
                           n2421);
   U1565 : OAI21_X1 port map( B1 => n1505, B2 => n1689, A => n2421, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U1566 : NAND2_X1 port map( A1 => n1443, A2 => n2492, ZN => n2491);
   U1567 : NOR2_X1 port map( A1 => n1711, A2 => n2491, ZN => n2494);
   U1568 : AOI211_X1 port map( C1 => n1711, C2 => n2491, A => n2494, B => n1804
                           , ZN => n400);
   U1569 : AOI22_X1 port map( A1 => n1309, A2 => 
                           datapath_i_alu_output_val_i_16_port, B1 => n1506, B2
                           => datapath_i_new_pc_value_decode_16_port, ZN => 
                           n2422);
   U1570 : OAI21_X1 port map( B1 => n1505, B2 => n1691, A => n2422, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U1571 : NAND2_X1 port map( A1 => n1441, A2 => n2494, ZN => n2493);
   U1572 : NOR2_X1 port map( A1 => n1712, A2 => n2493, ZN => n2496);
   U1573 : AOI211_X1 port map( C1 => n1712, C2 => n2493, A => n2496, B => n1804
                           , ZN => n405);
   U1574 : AOI22_X1 port map( A1 => n1309, A2 => 
                           datapath_i_alu_output_val_i_18_port, B1 => n1506, B2
                           => datapath_i_new_pc_value_decode_18_port, ZN => 
                           n2423);
   U1575 : OAI21_X1 port map( B1 => n1505, B2 => n1693, A => n2423, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U1576 : NAND2_X1 port map( A1 => n1439, A2 => n2496, ZN => n2495);
   U1577 : NOR2_X1 port map( A1 => n1713, A2 => n2495, ZN => n2498);
   U1578 : AOI211_X1 port map( C1 => n1713, C2 => n2495, A => n2498, B => n1804
                           , ZN => n415);
   U1579 : AOI22_X1 port map( A1 => n1309, A2 => 
                           datapath_i_alu_output_val_i_20_port, B1 => n1506, B2
                           => datapath_i_new_pc_value_decode_20_port, ZN => 
                           n2424);
   U1580 : OAI21_X1 port map( B1 => n1505, B2 => n1695, A => n2424, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U1581 : NAND2_X1 port map( A1 => n1437, A2 => n2498, ZN => n2497);
   U1582 : NOR2_X1 port map( A1 => n1714, A2 => n2497, ZN => n2500);
   U1583 : AOI211_X1 port map( C1 => n1714, C2 => n2497, A => n2500, B => n1804
                           , ZN => n420);
   U1584 : OAI211_X1 port map( C1 => n2426, C2 => n1435, A => n1803, B => n2425
                           , ZN => n2427);
   U1585 : NAND2_X1 port map( A1 => n1316, A2 => n2427, ZN => 
                           datapath_i_new_pc_value_decode_22_port);
   U1586 : AOI22_X1 port map( A1 => n1309, A2 => 
                           datapath_i_alu_output_val_i_22_port, B1 => n1506, B2
                           => datapath_i_new_pc_value_decode_22_port, ZN => 
                           n2428);
   U1587 : OAI21_X1 port map( B1 => n1505, B2 => n1697, A => n2428, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U1588 : NAND2_X1 port map( A1 => n1435, A2 => n2500, ZN => n2499);
   U1589 : NOR2_X1 port map( A1 => n1715, A2 => n2499, ZN => n2502);
   U1590 : AOI211_X1 port map( C1 => n1715, C2 => n2499, A => n2502, B => n1804
                           , ZN => n426);
   U1591 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_24_port, B1 => n1309,
                           B2 => datapath_i_alu_output_val_i_24_port, ZN => 
                           n2429);
   U1592 : OAI21_X1 port map( B1 => n1505, B2 => n1699, A => n2429, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U1593 : NAND2_X1 port map( A1 => n1433, A2 => n2502, ZN => n2501);
   U1594 : NOR2_X1 port map( A1 => n1716, A2 => n2501, ZN => n2504);
   U1595 : AOI211_X1 port map( C1 => n1716, C2 => n2501, A => n2504, B => n1804
                           , ZN => n431);
   U1596 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_26_port, B1 => n1309,
                           B2 => datapath_i_alu_output_val_i_26_port, ZN => 
                           n2430);
   U1597 : OAI21_X1 port map( B1 => n1783, B2 => n1701, A => n2430, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U1598 : NAND2_X1 port map( A1 => n1431, A2 => n2504, ZN => n2503);
   U1599 : NOR2_X1 port map( A1 => n1717, A2 => n2503, ZN => n2506);
   U1600 : AOI211_X1 port map( C1 => n1717, C2 => n2503, A => n2506, B => n1804
                           , ZN => n436);
   U1601 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_28_port, B1 => n1309,
                           B2 => datapath_i_alu_output_val_i_28_port, ZN => 
                           n2431);
   U1602 : OAI21_X1 port map( B1 => n1783, B2 => n1703, A => n2431, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U1603 : NAND2_X1 port map( A1 => n1429, A2 => n2506, ZN => n2505);
   U1604 : NOR2_X1 port map( A1 => n1718, A2 => n2505, ZN => n2507);
   U1605 : AOI211_X1 port map( C1 => n1718, C2 => n2505, A => n2507, B => n1804
                           , ZN => n441);
   U1606 : AOI22_X1 port map( A1 => n719, A2 => n2578, B1 => n1781, B2 => n2255
                           , ZN => n676);
   U1607 : NAND2_X1 port map( A1 => n2435, A2 => n1427, ZN => n2434);
   U1608 : XOR2_X1 port map( A => n1916, B => n2434, Z => n2432);
   U1609 : AOI22_X1 port map( A1 => n1803, A2 => n2432, B1 => n1745, B2 => 
                           n1460, ZN => datapath_i_new_pc_value_decode_31_port)
                           ;
   U1610 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_31_port, B1 => n1759,
                           B2 => datapath_i_alu_output_val_i_31_port, ZN => 
                           n2433);
   U1611 : OAI21_X1 port map( B1 => n1783, B2 => n1724, A => n2433, ZN => n1808
                           );
   U1612 : OAI211_X1 port map( C1 => n2435, C2 => n1427, A => n1803, B => n2434
                           , ZN => n2436);
   U1613 : NAND2_X1 port map( A1 => n1312, A2 => n2436, ZN => 
                           datapath_i_new_pc_value_decode_30_port);
   U1614 : AOI22_X1 port map( A1 => n1758, A2 => 
                           datapath_i_new_pc_value_decode_30_port, B1 => n1309,
                           B2 => datapath_i_alu_output_val_i_30_port, ZN => 
                           n2437);
   U1615 : OAI21_X1 port map( B1 => n1783, B2 => n1705, A => n2437, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   datapath_i_execute_stage_dp_n9 <= '0';
   U1617 : NOR4_X1 port map( A1 => n1394, A2 => n1393, A3 => n1721, A4 => n1780
                           , ZN => n2452);
   U1618 : NOR2_X1 port map( A1 => n1723, A2 => n1502, ZN => n2438);
   U1619 : AOI22_X1 port map( A1 => n2452, A2 => n1477, B1 => n1500, B2 => 
                           n2438, ZN => n2443);
   U1620 : NAND2_X1 port map( A1 => n1476, A2 => n1351, ZN => n2444);
   U1621 : NOR3_X1 port map( A1 => n1394, A2 => n1721, A3 => n1780, ZN => n2439
                           );
   U1622 : NAND3_X1 port map( A1 => n1393, A2 => n2439, A3 => n2572, ZN => 
                           n2456);
   U1623 : OAI21_X1 port map( B1 => n1719, B2 => n2444, A => n2456, ZN => n2440
                           );
   U1624 : NOR2_X1 port map( A1 => n1390, A2 => n1720, ZN => n2449);
   U1625 : OAI21_X1 port map( B1 => n2452, B2 => n2440, A => n2449, ZN => n2442
                           );
   U1626 : NAND2_X1 port map( A1 => n1417, A2 => n1350, ZN => n2441);
   U1627 : NAND4_X1 port map( A1 => n1305, A2 => n2443, A3 => n2442, A4 => 
                           n2441, ZN => cu_i_N264);
   U1628 : NOR2_X1 port map( A1 => n2444, A2 => n1395, ZN => n2445);
   U1629 : AOI21_X1 port map( B1 => n2445, B2 => n2449, A => n1350, ZN => n2454
                           );
   U1630 : NOR3_X1 port map( A1 => n1392, A2 => n2570, A3 => n2456, ZN => n2448
                           );
   U1631 : NAND3_X1 port map( A1 => n1723, A2 => n1842, A3 => n1500, ZN => 
                           n2446);
   U1632 : NAND2_X1 port map( A1 => n2446, A2 => n1495, ZN => n2447);
   U1633 : AOI211_X1 port map( C1 => n1501, C2 => n1782, A => n2448, B => n2447
                           , ZN => n2451);
   U1634 : NAND3_X1 port map( A1 => n2452, A2 => n2449, A3 => n1719, ZN => 
                           n2450);
   U1635 : NAND3_X1 port map( A1 => n2454, A2 => n2451, A3 => n2450, ZN => 
                           cu_i_N265);
   U1636 : OAI221_X1 port map( B1 => n1477, B2 => n1390, C1 => n1477, C2 => 
                           n1719, A => n2452, ZN => n2455);
   U1637 : OAI221_X1 port map( B1 => n1842, B2 => n1417, C1 => n1842, C2 => 
                           n1722, A => n1501, ZN => n2453);
   U1638 : OAI211_X1 port map( C1 => n1720, C2 => n2455, A => n2454, B => n2453
                           , ZN => cu_i_N266);
   U1639 : OAI221_X1 port map( B1 => n2456, B2 => n1720, C1 => n2456, C2 => 
                           n2570, A => n1349, ZN => cu_i_N267);
   U1640 : NAND2_X1 port map( A1 => n1801, A2 => n1485, ZN => cu_i_N274);
   U1641 : OAI21_X1 port map( B1 => n1513, B2 => n1510, A => n2459, ZN => n2457
                           );
   U1642 : NOR2_X1 port map( A1 => n1485, A2 => n2457, ZN => cu_i_N275);
   U1643 : NOR2_X1 port map( A1 => n1485, A2 => n1510, ZN => cu_i_N273);
   U1644 : AOI211_X1 port map( C1 => n2551, C2 => n2459, A => n2458, B => n2573
                           , ZN => cu_i_N276);
   U1645 : AOI211_X1 port map( C1 => n1801, C2 => n1458, A => n1485, B => n1725
                           , ZN => cu_i_N279);
   U1646 : NOR2_X1 port map( A1 => n2289, A2 => curr_instruction_to_cu_i_0_port
                           , ZN => n493);
   U1647 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => 
                           curr_instruction_to_cu_i_3_port, ZN => n492);
   U1648 : NAND3_X1 port map( A1 => n2295, A2 => n2461, A3 => n2460, ZN => 
                           n2464);
   U1649 : NAND4_X1 port map( A1 => n2290, A2 => n493, A3 => n492, A4 => n2462,
                           ZN => n2463);
   U1650 : OAI22_X1 port map( A1 => n2465, A2 => n2464, B1 => n2293, B2 => 
                           n2463, ZN => cu_i_cmd_word_8_port);
   U1651 : MUX2_X1 port map( A => n1332, B => cu_i_cmd_word_8_port, S => n719, 
                           Z => alu_cin_i);
   U1652 : NAND2_X1 port map( A1 => n1496, A2 => n2255, ZN => n2466);
   U1653 : OAI21_X1 port map( B1 => n2255, B2 => n2569, A => n2466, ZN => 
                           cu_i_cw2_4_port);
   U1654 : MUX2_X1 port map( A => n1499, B => n1425, S => n719, Z => 
                           cu_i_cw2_7_port);
   U1655 : MUX2_X1 port map( A => n1459, B => n1424, S => n719, Z => 
                           cu_i_cw2_8_port);
   U1656 : AOI22_X1 port map( A1 => n1801, A2 => n1403, B1 => IRAM_DATA(13), B2
                           => n2554, ZN => n2257);
   U1657 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_14_port, A2 => 
                           curr_instruction_to_cu_i_15_port, A3 => 
                           curr_instruction_to_cu_i_12_port, A4 => 
                           curr_instruction_to_cu_i_11_port, ZN => n2467);
   U1658 : AOI21_X1 port map( B1 => n2257, B2 => n2467, A => n2294, ZN => n2471
                           );
   U1659 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_19_port, A2 => 
                           curr_instruction_to_cu_i_20_port, A3 => 
                           curr_instruction_to_cu_i_17_port, A4 => 
                           curr_instruction_to_cu_i_16_port, ZN => n2469);
   U1660 : AOI21_X1 port map( B1 => n2258, B2 => n2469, A => n2468, ZN => n2470
                           );
   U1661 : AOI211_X1 port map( C1 => n2472, C2 => n2294, A => n2471, B => n2470
                           , ZN => n2475);
   U1662 : AOI211_X1 port map( C1 => n1475, C2 => n2553, A => 
                           cu_i_cmd_word_4_port, B => cu_i_n135, ZN => n2473);
   U1663 : OAI21_X1 port map( B1 => n2475, B2 => n2474, A => n2473, ZN => 
                           cu_i_n153);
   U1664 : AND2_X1 port map( A1 => n1475, A2 => n1331, ZN => cu_i_n3);
   U1665 : MUX2_X1 port map( A => n1301, B => n1423, S => n719, Z => 
                           cu_i_cw2_6_port);
   U1666 : MUX2_X1 port map( A => n1498, B => n1422, S => n719, Z => 
                           cu_i_cw2_5_port);
   U1667 : MUX2_X1 port map( A => IRAM_DATA(25), B => n1415, S => n1509, Z => 
                           datapath_i_n9);
   U1668 : MUX2_X1 port map( A => IRAM_DATA(24), B => n1414, S => n1509, Z => 
                           datapath_i_n10);
   U1669 : MUX2_X1 port map( A => IRAM_DATA(23), B => n1413, S => n1801, Z => 
                           datapath_i_n11);
   U1670 : MUX2_X1 port map( A => IRAM_DATA(22), B => n1412, S => n1801, Z => 
                           datapath_i_n12);
   U1671 : MUX2_X1 port map( A => IRAM_DATA(21), B => n1411, S => n1801, Z => 
                           datapath_i_n13);
   U1672 : MUX2_X1 port map( A => IRAM_DATA(10), B => n1400, S => n1509, Z => 
                           datapath_i_n14);
   U1673 : MUX2_X1 port map( A => IRAM_DATA(9), B => n1399, S => n1509, Z => 
                           datapath_i_n15);
   U1674 : MUX2_X1 port map( A => IRAM_DATA(8), B => n1398, S => n1509, Z => 
                           datapath_i_n16);
   U1675 : MUX2_X1 port map( A => IRAM_DATA(7), B => n1397, S => n1509, Z => 
                           datapath_i_n17);
   U1676 : MUX2_X1 port map( A => IRAM_DATA(6), B => n1396, S => n1509, Z => 
                           datapath_i_n18);
   U1677 : NAND2_X1 port map( A1 => n1846, A2 => n1457, ZN => n2480);
   U1678 : OAI211_X1 port map( C1 => n1846, C2 => IRAM_ADDRESS_3_port, A => 
                           n1746, B => n2480, ZN => n2478);
   U1679 : OAI211_X1 port map( C1 => datapath_i_new_pc_value_mem_stage_i_2_port
                           , C2 => datapath_i_new_pc_value_mem_stage_i_3_port, 
                           A => n1804, B => n2476, ZN => n2477);
   U1680 : NAND2_X1 port map( A1 => n2478, A2 => n2477, ZN => 
                           datapath_i_new_pc_value_decode_3_port);
   U1681 : OAI211_X1 port map( C1 => n2479, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n1804, B => n519, ZN => n524);
   U1682 : INV_X1 port map( A => n2480, ZN => n2482);
   U1683 : OAI211_X1 port map( C1 => n2482, C2 => IRAM_ADDRESS_4_port, A => 
                           n1746, B => n2481, ZN => n523);
   U1684 : OAI211_X1 port map( C1 => n2484, C2 => IRAM_ADDRESS_6_port, A => 
                           n1754, B => n2483, ZN => n529);
   U1685 : OAI211_X1 port map( C1 => n2486, C2 => IRAM_ADDRESS_8_port, A => 
                           n1754, B => n2485, ZN => n535);
   U1686 : OAI211_X1 port map( C1 => n2488, C2 => IRAM_ADDRESS_10_port, A => 
                           n1754, B => n2487, ZN => n541);
   U1687 : OAI211_X1 port map( C1 => n2490, C2 => IRAM_ADDRESS_12_port, A => 
                           n1754, B => n2489, ZN => n547);
   U1688 : OAI211_X1 port map( C1 => n2492, C2 => IRAM_ADDRESS_14_port, A => 
                           n1754, B => n2491, ZN => n553);
   U1689 : OAI211_X1 port map( C1 => n2494, C2 => IRAM_ADDRESS_16_port, A => 
                           n1754, B => n2493, ZN => n559);
   U1690 : OAI211_X1 port map( C1 => n2496, C2 => IRAM_ADDRESS_18_port, A => 
                           n1754, B => n2495, ZN => n565);
   U1691 : OAI211_X1 port map( C1 => n2498, C2 => IRAM_ADDRESS_20_port, A => 
                           n1754, B => n2497, ZN => n571);
   U1692 : OAI211_X1 port map( C1 => n2500, C2 => IRAM_ADDRESS_22_port, A => 
                           n1746, B => n2499, ZN => n577);
   U1693 : OAI211_X1 port map( C1 => n2502, C2 => IRAM_ADDRESS_24_port, A => 
                           n1754, B => n2501, ZN => n583);
   U1694 : OAI211_X1 port map( C1 => n2504, C2 => IRAM_ADDRESS_26_port, A => 
                           n1754, B => n2503, ZN => n589);
   U1695 : OAI211_X1 port map( C1 => n2506, C2 => IRAM_ADDRESS_28_port, A => 
                           n1746, B => n2505, ZN => n595);
   U1696 : NAND2_X1 port map( A1 => n1427, A2 => n2507, ZN => n2508);
   U1697 : OAI211_X1 port map( C1 => n2507, C2 => IRAM_ADDRESS_30_port, A => 
                           n1754, B => n2508, ZN => n601);
   U1698 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n2508, Z => n606);
   U1699 : AND2_X1 port map( A1 => n1781, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U1700 : OAI21_X1 port map( B1 => n2300, B2 => n2509, A => n2511, ZN => 
                           read_rf_p2_i);
   U1701 : OAI221_X1 port map( B1 => n2512, B2 => n2258, C1 => n2511, C2 => 
                           n2257, A => n2510, ZN => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port);
   U1702 : OAI21_X1 port map( B1 => n1888, B2 => n2513, A => n2075, ZN => 
                           datapath_i_decode_stage_dp_n44);
   U1703 : OAI21_X1 port map( B1 => n1891, B2 => n2513, A => n2072, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U1704 : OAI21_X1 port map( B1 => n1868, B2 => n2513, A => n2071, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U1705 : OAI21_X1 port map( B1 => n1867, B2 => n2513, A => n2070, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U1706 : OAI21_X1 port map( B1 => n1869, B2 => n2513, A => n2069, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U1707 : OAI21_X1 port map( B1 => n1895, B2 => n2513, A => n2068, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U1708 : OAI21_X1 port map( B1 => n1894, B2 => n2513, A => n2067, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U1709 : OAI21_X1 port map( B1 => n1897, B2 => n2513, A => n2066, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U1710 : OAI21_X1 port map( B1 => n1890, B2 => n2513, A => n2065, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U1711 : OAI21_X1 port map( B1 => n1870, B2 => n2513, A => n2064, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U1712 : OAI21_X1 port map( B1 => n1889, B2 => n2513, A => n2063, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U1713 : OAI21_X1 port map( B1 => n1874, B2 => n2513, A => n2062, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U1714 : OAI21_X1 port map( B1 => n1896, B2 => n2513, A => n2061, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U1715 : OAI21_X1 port map( B1 => n1873, B2 => n2513, A => n2060, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U1716 : OAI21_X1 port map( B1 => n1871, B2 => n2513, A => n2059, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U1717 : OAI21_X1 port map( B1 => n1872, B2 => n2513, A => n2058, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U1718 : OAI21_X1 port map( B1 => n1876, B2 => n2513, A => n2057, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U1719 : OAI21_X1 port map( B1 => n1875, B2 => n2513, A => n2056, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U1720 : OAI21_X1 port map( B1 => n1885, B2 => n2513, A => n2055, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U1721 : OAI21_X1 port map( B1 => n1878, B2 => n2513, A => n2054, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U1722 : OAI21_X1 port map( B1 => n1892, B2 => n2513, A => n2053, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U1723 : OAI21_X1 port map( B1 => n1877, B2 => n2513, A => n2052, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U1724 : OAI21_X1 port map( B1 => n1880, B2 => n2513, A => n2051, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U1725 : OAI21_X1 port map( B1 => n1879, B2 => n2513, A => n2050, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U1726 : OAI21_X1 port map( B1 => n1884, B2 => n2513, A => n2049, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U1727 : OAI21_X1 port map( B1 => n1883, B2 => n2513, A => n2048, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U1728 : OAI21_X1 port map( B1 => n1886, B2 => n2513, A => n2047, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U1729 : OAI21_X1 port map( B1 => n1882, B2 => n2513, A => n2046, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U1730 : OAI21_X1 port map( B1 => n1893, B2 => n2513, A => n2045, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U1731 : OAI21_X1 port map( B1 => n1881, B2 => n2513, A => n2044, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U1732 : OAI21_X1 port map( B1 => n1887, B2 => n2513, A => n2043, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U1733 : OAI21_X1 port map( B1 => n1844, B2 => n2513, A => n2042, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U1734 : AOI21_X1 port map( B1 => n2516, B2 => n2515, A => n2514, ZN => n2517
                           );
   U1735 : NOR2_X1 port map( A1 => n2518, A2 => n2517, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U1736 : AOI22_X1 port map( A1 => n719, A2 => cu_i_cmd_word_6_port, B1 => 
                           n1452, B2 => n2255, ZN => n2532);
   U1737 : NOR4_X1 port map( A1 => n1641, A2 => n1643, A3 => n1645, A4 => n1647
                           , ZN => n2522);
   U1738 : NOR4_X1 port map( A1 => n1649, A2 => n1651, A3 => n1653, A4 => n1655
                           , ZN => n2521);
   U1739 : NOR4_X1 port map( A1 => n1625, A2 => n1627, A3 => n1629, A4 => n1631
                           , ZN => n2520);
   U1740 : NOR4_X1 port map( A1 => n1633, A2 => n1635, A3 => n1637, A4 => n1639
                           , ZN => n2519);
   U1741 : NAND4_X1 port map( A1 => n2522, A2 => n2521, A3 => n2520, A4 => 
                           n2519, ZN => n2528);
   U1742 : NOR4_X1 port map( A1 => n1663, A2 => n1617, A3 => n1619, A4 => n1621
                           , ZN => n2526);
   U1743 : NOR4_X1 port map( A1 => n1613, A2 => n1614, A3 => n1615, A4 => n1661
                           , ZN => n2525);
   U1744 : NOR4_X1 port map( A1 => n1667, A2 => n1669, A3 => n1657, A4 => n1659
                           , ZN => n2524);
   U1745 : NOR4_X1 port map( A1 => n1623, A2 => n1671, A3 => n1673, A4 => n1665
                           , ZN => n2523);
   U1746 : NAND4_X1 port map( A1 => n2526, A2 => n2525, A3 => n2524, A4 => 
                           n2523, ZN => n2527);
   U1747 : NOR2_X1 port map( A1 => n2528, A2 => n2527, ZN => n2530);
   U1748 : AOI22_X1 port map( A1 => n719, A2 => cu_i_cmd_word_7_port, B1 => 
                           n1347, B2 => n2255, ZN => n2529);
   U1749 : NAND2_X1 port map( A1 => n2530, A2 => n2529, ZN => n2531);
   U1750 : OAI22_X1 port map( A1 => n2532, A2 => n2531, B1 => n2530, B2 => 
                           n2529, ZN => n717);
   U1751 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_7_port);
   U1752 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_8_port);
   U1753 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_9_port);
   U1754 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_10_port);
   U1755 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_11_port);
   U1756 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_12_port);
   U1757 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_13_port);
   U1758 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, S 
                           => n1774, Z => datapath_i_val_immediate_i_14_port);
   U1759 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_15_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_15_port);
   U1760 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_16_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_16_port);
   U1761 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_17_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_17_port);
   U1762 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_18_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_18_port);
   U1763 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_19_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_19_port);
   U1764 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_20_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_20_port);
   U1765 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_21_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_21_port);
   U1766 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_22_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_22_port);
   U1767 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_23_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_23_port);
   U1768 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_24_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_24_port);
   U1769 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_25_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_25_port);
   U1770 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_26_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_26_port, S 
                           => n1776, Z => datapath_i_val_immediate_i_26_port);
   U1771 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_0_port);
   U1772 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_27_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_27_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_27_port);
   U1773 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_28_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_28_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_28_port);
   U1774 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_29_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_29_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_29_port);
   U1775 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_30_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_30_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_30_port);
   U1776 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_31_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_31_port);
   U1777 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_1_port);
   U1778 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_2_port);
   U1779 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_3_port);
   U1780 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_4_port);
   U1781 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_5_port);
   U1782 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, S 
                           => n1777, Z => datapath_i_val_immediate_i_6_port);
   U1783 : MUX2_X1 port map( A => n1383, B => n1539, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U1784 : MUX2_X1 port map( A => n1382, B => n1542, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U1785 : MUX2_X1 port map( A => n1381, B => n1545, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U1786 : MUX2_X1 port map( A => n1380, B => n1548, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_10_port);
   U1787 : MUX2_X1 port map( A => n1379, B => n1551, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_11_port);
   U1788 : MUX2_X1 port map( A => n1378, B => n1554, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_12_port);
   U1789 : MUX2_X1 port map( A => n1377, B => n1557, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_13_port);
   U1790 : MUX2_X1 port map( A => n1376, B => n1560, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_14_port);
   U1791 : MUX2_X1 port map( A => n1375, B => n1563, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_15_port);
   U1792 : MUX2_X1 port map( A => n1374, B => n1566, S => n1333, Z => 
                           datapath_i_execute_stage_dp_opb_16_port);
   U1793 : MUX2_X1 port map( A => n1373, B => n1569, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_17_port);
   U1794 : MUX2_X1 port map( A => n1372, B => n1572, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_18_port);
   U1795 : MUX2_X1 port map( A => n1371, B => n1575, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_19_port);
   U1796 : MUX2_X1 port map( A => n1370, B => n1578, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_20_port);
   U1797 : MUX2_X1 port map( A => n1369, B => n1581, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_21_port);
   U1798 : MUX2_X1 port map( A => n1368, B => n1584, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_22_port);
   U1799 : MUX2_X1 port map( A => n1367, B => n1587, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_23_port);
   U1800 : MUX2_X1 port map( A => n1366, B => n1590, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_24_port);
   U1801 : MUX2_X1 port map( A => n1365, B => n1593, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U1802 : MUX2_X1 port map( A => n1364, B => n1596, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U1803 : MUX2_X1 port map( A => n1362, B => n1599, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U1804 : MUX2_X1 port map( A => n1361, B => n1602, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U1805 : MUX2_X1 port map( A => n1360, B => n1605, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U1806 : MUX2_X1 port map( A => n1359, B => n1608, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U1807 : MUX2_X1 port map( A => n1358, B => n1611, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U1808 : MUX2_X1 port map( A => n1352, B => n1536, S => n1728, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U1809 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_13_port, B1 => n1802,
                           B2 => n1636, ZN => n2533);
   U1810 : OAI21_X1 port map( B1 => n1507, B2 => n1688, A => n2533, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U1811 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_17_port, B1 => n2541,
                           B2 => n1644, ZN => n2534);
   U1812 : OAI21_X1 port map( B1 => n1507, B2 => n1692, A => n2534, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U1813 : AOI22_X1 port map( A1 => n1802, A2 => n1652, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_21_port, ZN => n2535)
                           ;
   U1814 : OAI21_X1 port map( B1 => n2544, B2 => n1696, A => n2535, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U1815 : AOI22_X1 port map( A1 => n1802, A2 => n1654, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_22_port, ZN => n2536)
                           ;
   U1816 : OAI21_X1 port map( B1 => n1507, B2 => n1697, A => n2536, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U1817 : AOI22_X1 port map( A1 => n2541, A2 => n1656, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_23_port, ZN => n2537)
                           ;
   U1818 : OAI21_X1 port map( B1 => n1507, B2 => n1698, A => n2537, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U1819 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_25_port, B1 => n2541,
                           B2 => n1660, ZN => n2538);
   U1820 : OAI21_X1 port map( B1 => n2544, B2 => n1700, A => n2538, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U1821 : NOR2_X1 port map( A1 => n1773, A2 => n2256, ZN => n703);
   U1822 : AOI22_X1 port map( A1 => n1758, A2 => n1388, B1 => n1759, B2 => 
                           datapath_i_alu_output_val_i_0_port, ZN => n2539);
   U1823 : OAI21_X1 port map( B1 => n1505, B2 => n1675, A => n2539, ZN => 
                           datapath_i_fetch_stage_dp_N39);
   U1824 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N39, B => 
                           IRAM_ADDRESS_0_port, S => n1746, Z => 
                           datapath_i_new_pc_value_decode_0_port);
   U1825 : AOI22_X1 port map( A1 => n2256, A2 => n1613, B1 => n703, B2 => 
                           datapath_i_new_pc_value_decode_0_port, ZN => n692);
   U1826 : OAI21_X1 port map( B1 => n1507, B2 => n1675, A => n1308, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U1827 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_27_port, B1 => n1802,
                           B2 => n1664, ZN => n2540);
   U1828 : OAI21_X1 port map( B1 => n1507, B2 => n1702, A => n2540, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U1829 : AOI22_X1 port map( A1 => n2541, A2 => n1668, B1 => n1478, B2 => 
                           datapath_i_new_pc_value_decode_29_port, ZN => n2542)
                           ;
   U1830 : OAI21_X1 port map( B1 => n2544, B2 => n1704, A => n2542, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U1831 : AOI22_X1 port map( A1 => n1727, A2 => 
                           datapath_i_new_pc_value_decode_30_port, B1 => n1802,
                           B2 => n1670, ZN => n2543);
   U1832 : OAI21_X1 port map( B1 => n2544, B2 => n1705, A => n2543, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U1833 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n1727, B1 => n1802, B2 => n1672, ZN => n2545);
   U1834 : OAI21_X1 port map( B1 => n1724, B2 => n1507, A => n2545, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U1835 : AOI22_X1 port map( A1 => n1758, A2 => n1385, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_1_port, ZN => n2546);
   U1836 : OAI21_X1 port map( B1 => n1505, B2 => n1676, A => n2546, ZN => 
                           datapath_i_fetch_stage_dp_N40);
   U1837 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N40, B => 
                           IRAM_ADDRESS_1_port, S => n1746, Z => 
                           datapath_i_new_pc_value_decode_1_port);
   U1838 : AOI22_X1 port map( A1 => n2256, A2 => n1614, B1 => n703, B2 => 
                           datapath_i_new_pc_value_decode_1_port, ZN => n699);
   U1839 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port
                           , A => n2555, ZN => n2547);
   U1840 : AOI22_X1 port map( A1 => n1804, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B1 => 
                           n1746, B2 => n2547, ZN => 
                           datapath_i_new_pc_value_decode_2_port);
   U1841 : AOI22_X1 port map( A1 => n2256, A2 => n1615, B1 => n703, B2 => 
                           datapath_i_new_pc_value_decode_2_port, ZN => n700);
   U1842 : OAI21_X1 port map( B1 => n1507, B2 => n1677, A => n1306, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U1843 : AOI22_X1 port map( A1 => n1802, A2 => n1616, B1 => n1478, B2 => 
                           n1328, ZN => n2548);
   U1844 : OAI21_X1 port map( B1 => n1507, B2 => n1678, A => n2548, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U1845 : AOI222_X1 port map( A1 => n2558, A2 => n2549, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_21_port, C1 => 
                           datapath_i_new_pc_value_decode_21_port, C2 => n1506,
                           ZN => n2287);
   U1846 : AOI222_X1 port map( A1 => n2559, A2 => n2549, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_19_port, C1 => 
                           datapath_i_new_pc_value_decode_19_port, C2 => n1506,
                           ZN => n2286);
   U1847 : AOI222_X1 port map( A1 => n2560, A2 => n2549, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_17_port, C1 => 
                           datapath_i_new_pc_value_decode_17_port, C2 => n1506,
                           ZN => n2285);
   U1848 : AOI222_X1 port map( A1 => n2561, A2 => n2549, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_13_port, C1 => 
                           datapath_i_new_pc_value_decode_13_port, C2 => n1758,
                           ZN => n2284);
   U1849 : AOI222_X1 port map( A1 => n2562, A2 => n2549, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_15_port, C1 => 
                           datapath_i_new_pc_value_decode_15_port, C2 => n1758,
                           ZN => n2283);
   U1850 : AOI222_X1 port map( A1 => n2563, A2 => n2549, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_23_port, C1 => 
                           datapath_i_new_pc_value_decode_23_port, C2 => n1758,
                           ZN => n2282);
   U1851 : AOI222_X1 port map( A1 => n2549, A2 => n2556, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_25_port, C1 => 
                           datapath_i_new_pc_value_decode_25_port, C2 => n1758,
                           ZN => n2281);
   U1852 : AOI222_X1 port map( A1 => n2564, A2 => n2549, B1 => n1759, B2 => 
                           datapath_i_alu_output_val_i_7_port, C1 => 
                           datapath_i_new_pc_value_decode_7_port, C2 => n1758, 
                           ZN => n2280);
   U1853 : AOI222_X1 port map( A1 => n2565, A2 => n2549, B1 => n1759, B2 => 
                           datapath_i_alu_output_val_i_9_port, C1 => 
                           datapath_i_new_pc_value_decode_9_port, C2 => n1758, 
                           ZN => n2278);
   U1854 : AOI222_X1 port map( A1 => n2566, A2 => n2549, B1 => n1759, B2 => 
                           datapath_i_alu_output_val_i_11_port, C1 => 
                           datapath_i_new_pc_value_decode_11_port, C2 => n1506,
                           ZN => n2277);
   U1855 : AOI222_X1 port map( A1 => n2567, A2 => n2550, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_27_port, C1 => 
                           datapath_i_new_pc_value_decode_27_port, C2 => n1758,
                           ZN => n2276);
   U1856 : AOI222_X1 port map( A1 => n2568, A2 => n2550, B1 => n1309, B2 => 
                           datapath_i_alu_output_val_i_29_port, C1 => 
                           datapath_i_new_pc_value_decode_29_port, C2 => n1758,
                           ZN => n2275);
   U1857 : MUX2_X1 port map( A => n1423, B => n1779, S => n719, Z => n2254);

end SYN_dlx_rtl;
