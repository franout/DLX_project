//
//					\\\ Sapere Aude ///
//
// -----------------------------------------------------------------------------
// Copyright (c) 2014-2020 All rights reserved
// -----------------------------------------------------------------------------
// Author : Angione Francesco s262620@studenti.polito.it franout@Github.com
// File   : property_def.svh
// Create : 2020-08-01 16:14:31
// Revise : 2020-08-01 16:14:31
// Editor : sublime text3, tab size (4)
// Description: Defintion of all propery and sequences for the DLX top level entity
// -----------------------------------------------------------------------------
`ifndef __PROPERTY_DEF_SVH
`define __PROPERTY_DEF_SVH




`endif //__PROPERTY_DEF_SVH