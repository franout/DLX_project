
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type TYPE_OP_ALU is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCLSL, FUNCLSR, 
   GE, LE, NE);
attribute ENUM_ENCODING of TYPE_OP_ALU : type is 
   "0000 0001 0010 0011 0100 0101 0110 0111 1000 1001 1010";
   
   -- Declarations for conversion functions.
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
               std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- enum type to std_logic_vector function
   function TYPE_OP_ALU_to_std_logic_vector(arg : in TYPE_OP_ALU) return 
   std_logic_vector is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when ADD => return "0000";
         when SUB => return "0001";
         when MULT => return "0010";
         when BITAND => return "0011";
         when BITOR => return "0100";
         when BITXOR => return "0101";
         when FUNCLSL => return "0110";
         when FUNCLSR => return "0111";
         when GE => return "1000";
         when LE => return "1001";
         when NE => return "1010";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "0000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity general_alu_N32 is

   port( clk : in std_logic;  zero_mul_detect, mul_exeception : out std_logic; 
         FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  cin, signed_notsigned : in std_logic;
         overflow : out std_logic;  OUTALU : out std_logic_vector (31 downto 0)
         ;  rst_BAR : in std_logic);

end general_alu_N32;

architecture SYN_behavioural of general_alu_N32 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal DATA2_I_31_port, DATA2_I_30_port, DATA2_I_29_port, DATA2_I_28_port, 
      DATA2_I_27_port, DATA2_I_26_port, DATA2_I_25_port, DATA2_I_24_port, 
      DATA2_I_23_port, DATA2_I_22_port, DATA2_I_21_port, DATA2_I_20_port, 
      DATA2_I_19_port, DATA2_I_18_port, DATA2_I_17_port, DATA2_I_16_port, 
      DATA2_I_15_port, DATA2_I_14_port, DATA2_I_13_port, DATA2_I_12_port, 
      DATA2_I_11_port, DATA2_I_10_port, DATA2_I_9_port, DATA2_I_8_port, 
      DATA2_I_7_port, DATA2_I_6_port, DATA2_I_5_port, DATA2_I_4_port, 
      DATA2_I_3_port, DATA2_I_2_port, DATA2_I_1_port, DATA2_I_0_port, 
      data1_mul_15_port, data1_mul_14_port, data1_mul_13_port, 
      data1_mul_12_port, data1_mul_11_port, data1_mul_10_port, data1_mul_9_port
      , data1_mul_8_port, data1_mul_7_port, data1_mul_6_port, data1_mul_5_port,
      data1_mul_4_port, data1_mul_3_port, data1_mul_2_port, data1_mul_1_port, 
      data1_mul_0_port, data2_mul_15_port, data2_mul_14_port, data2_mul_13_port
      , data2_mul_12_port, data2_mul_11_port, data2_mul_10_port, 
      data2_mul_9_port, data2_mul_8_port, data2_mul_7_port, data2_mul_6_port, 
      data2_mul_5_port, data2_mul_4_port, data2_mul_3_port, data2_mul_2_port, 
      data2_mul_1_port, dataout_mul_31_port, dataout_mul_30_port, 
      dataout_mul_29_port, dataout_mul_28_port, dataout_mul_27_port, 
      dataout_mul_26_port, dataout_mul_25_port, dataout_mul_24_port, 
      dataout_mul_23_port, dataout_mul_22_port, dataout_mul_21_port, 
      dataout_mul_20_port, dataout_mul_19_port, dataout_mul_18_port, 
      dataout_mul_17_port, dataout_mul_16_port, dataout_mul_15_port, 
      dataout_mul_13_port, dataout_mul_12_port, dataout_mul_11_port, 
      dataout_mul_10_port, dataout_mul_9_port, dataout_mul_8_port, 
      dataout_mul_7_port, dataout_mul_6_port, dataout_mul_5_port, 
      dataout_mul_4_port, dataout_mul_3_port, dataout_mul_2_port, 
      dataout_mul_1_port, dataout_mul_0_port, N2517, N2518, N2519, N2520, N2521
      , N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, 
      N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, 
      N2542, N2543, N2544, N2545, N2546, N2547, N2548, n553, 
      boothmul_pipelined_i_muxes_in_7_232_port, 
      boothmul_pipelined_i_muxes_in_7_231_port, 
      boothmul_pipelined_i_muxes_in_7_230_port, 
      boothmul_pipelined_i_muxes_in_7_229_port, 
      boothmul_pipelined_i_muxes_in_7_228_port, 
      boothmul_pipelined_i_muxes_in_7_227_port, 
      boothmul_pipelined_i_muxes_in_7_226_port, 
      boothmul_pipelined_i_muxes_in_7_225_port, 
      boothmul_pipelined_i_muxes_in_7_224_port, 
      boothmul_pipelined_i_muxes_in_7_223_port, 
      boothmul_pipelined_i_muxes_in_7_222_port, 
      boothmul_pipelined_i_muxes_in_7_221_port, 
      boothmul_pipelined_i_muxes_in_7_220_port, 
      boothmul_pipelined_i_muxes_in_7_219_port, 
      boothmul_pipelined_i_muxes_in_7_218_port, 
      boothmul_pipelined_i_muxes_in_7_217_port, 
      boothmul_pipelined_i_muxes_in_7_76_port, 
      boothmul_pipelined_i_muxes_in_7_75_port, 
      boothmul_pipelined_i_muxes_in_7_74_port, 
      boothmul_pipelined_i_muxes_in_7_73_port, 
      boothmul_pipelined_i_muxes_in_7_72_port, 
      boothmul_pipelined_i_muxes_in_7_71_port, 
      boothmul_pipelined_i_muxes_in_7_70_port, 
      boothmul_pipelined_i_muxes_in_7_69_port, 
      boothmul_pipelined_i_muxes_in_7_68_port, 
      boothmul_pipelined_i_muxes_in_7_67_port, 
      boothmul_pipelined_i_muxes_in_7_66_port, 
      boothmul_pipelined_i_muxes_in_7_65_port, 
      boothmul_pipelined_i_muxes_in_7_64_port, 
      boothmul_pipelined_i_muxes_in_7_63_port, 
      boothmul_pipelined_i_muxes_in_7_62_port, 
      boothmul_pipelined_i_muxes_in_6_218_port, 
      boothmul_pipelined_i_muxes_in_6_217_port, 
      boothmul_pipelined_i_muxes_in_6_216_port, 
      boothmul_pipelined_i_muxes_in_6_215_port, 
      boothmul_pipelined_i_muxes_in_6_214_port, 
      boothmul_pipelined_i_muxes_in_6_213_port, 
      boothmul_pipelined_i_muxes_in_6_212_port, 
      boothmul_pipelined_i_muxes_in_6_211_port, 
      boothmul_pipelined_i_muxes_in_6_210_port, 
      boothmul_pipelined_i_muxes_in_6_209_port, 
      boothmul_pipelined_i_muxes_in_6_208_port, 
      boothmul_pipelined_i_muxes_in_6_207_port, 
      boothmul_pipelined_i_muxes_in_6_206_port, 
      boothmul_pipelined_i_muxes_in_6_205_port, 
      boothmul_pipelined_i_muxes_in_6_204_port, 
      boothmul_pipelined_i_muxes_in_6_203_port, 
      boothmul_pipelined_i_muxes_in_6_73_port, 
      boothmul_pipelined_i_muxes_in_6_72_port, 
      boothmul_pipelined_i_muxes_in_6_71_port, 
      boothmul_pipelined_i_muxes_in_6_70_port, 
      boothmul_pipelined_i_muxes_in_6_69_port, 
      boothmul_pipelined_i_muxes_in_6_68_port, 
      boothmul_pipelined_i_muxes_in_6_67_port, 
      boothmul_pipelined_i_muxes_in_6_66_port, 
      boothmul_pipelined_i_muxes_in_6_65_port, 
      boothmul_pipelined_i_muxes_in_6_64_port, 
      boothmul_pipelined_i_muxes_in_6_63_port, 
      boothmul_pipelined_i_muxes_in_6_62_port, 
      boothmul_pipelined_i_muxes_in_6_61_port, 
      boothmul_pipelined_i_muxes_in_6_60_port, 
      boothmul_pipelined_i_muxes_in_6_59_port, 
      boothmul_pipelined_i_muxes_in_6_58_port, 
      boothmul_pipelined_i_muxes_in_5_205_port, 
      boothmul_pipelined_i_muxes_in_5_204_port, 
      boothmul_pipelined_i_muxes_in_5_203_port, 
      boothmul_pipelined_i_muxes_in_5_202_port, 
      boothmul_pipelined_i_muxes_in_5_201_port, 
      boothmul_pipelined_i_muxes_in_5_200_port, 
      boothmul_pipelined_i_muxes_in_5_199_port, 
      boothmul_pipelined_i_muxes_in_5_198_port, 
      boothmul_pipelined_i_muxes_in_5_197_port, 
      boothmul_pipelined_i_muxes_in_5_196_port, 
      boothmul_pipelined_i_muxes_in_5_195_port, 
      boothmul_pipelined_i_muxes_in_5_194_port, 
      boothmul_pipelined_i_muxes_in_5_193_port, 
      boothmul_pipelined_i_muxes_in_5_192_port, 
      boothmul_pipelined_i_muxes_in_5_191_port, 
      boothmul_pipelined_i_muxes_in_5_190_port, 
      boothmul_pipelined_i_muxes_in_5_189_port, 
      boothmul_pipelined_i_muxes_in_5_68_port, 
      boothmul_pipelined_i_muxes_in_5_67_port, 
      boothmul_pipelined_i_muxes_in_5_66_port, 
      boothmul_pipelined_i_muxes_in_5_65_port, 
      boothmul_pipelined_i_muxes_in_5_64_port, 
      boothmul_pipelined_i_muxes_in_5_63_port, 
      boothmul_pipelined_i_muxes_in_5_62_port, 
      boothmul_pipelined_i_muxes_in_5_61_port, 
      boothmul_pipelined_i_muxes_in_5_60_port, 
      boothmul_pipelined_i_muxes_in_5_59_port, 
      boothmul_pipelined_i_muxes_in_5_58_port, 
      boothmul_pipelined_i_muxes_in_5_57_port, 
      boothmul_pipelined_i_muxes_in_5_56_port, 
      boothmul_pipelined_i_muxes_in_5_55_port, 
      boothmul_pipelined_i_muxes_in_5_54_port, 
      boothmul_pipelined_i_muxes_in_4_190_port, 
      boothmul_pipelined_i_muxes_in_4_189_port, 
      boothmul_pipelined_i_muxes_in_4_188_port, 
      boothmul_pipelined_i_muxes_in_4_187_port, 
      boothmul_pipelined_i_muxes_in_4_186_port, 
      boothmul_pipelined_i_muxes_in_4_185_port, 
      boothmul_pipelined_i_muxes_in_4_184_port, 
      boothmul_pipelined_i_muxes_in_4_183_port, 
      boothmul_pipelined_i_muxes_in_4_182_port, 
      boothmul_pipelined_i_muxes_in_4_181_port, 
      boothmul_pipelined_i_muxes_in_4_180_port, 
      boothmul_pipelined_i_muxes_in_4_179_port, 
      boothmul_pipelined_i_muxes_in_4_178_port, 
      boothmul_pipelined_i_muxes_in_4_177_port, 
      boothmul_pipelined_i_muxes_in_4_176_port, 
      boothmul_pipelined_i_muxes_in_4_175_port, 
      boothmul_pipelined_i_muxes_in_4_65_port, 
      boothmul_pipelined_i_muxes_in_4_64_port, 
      boothmul_pipelined_i_muxes_in_4_63_port, 
      boothmul_pipelined_i_muxes_in_4_62_port, 
      boothmul_pipelined_i_muxes_in_4_61_port, 
      boothmul_pipelined_i_muxes_in_4_60_port, 
      boothmul_pipelined_i_muxes_in_4_59_port, 
      boothmul_pipelined_i_muxes_in_4_58_port, 
      boothmul_pipelined_i_muxes_in_4_57_port, 
      boothmul_pipelined_i_muxes_in_4_56_port, 
      boothmul_pipelined_i_muxes_in_4_55_port, 
      boothmul_pipelined_i_muxes_in_4_54_port, 
      boothmul_pipelined_i_muxes_in_4_53_port, 
      boothmul_pipelined_i_muxes_in_4_52_port, 
      boothmul_pipelined_i_muxes_in_4_51_port, 
      boothmul_pipelined_i_muxes_in_4_50_port, 
      boothmul_pipelined_i_muxes_in_3_177_port, 
      boothmul_pipelined_i_muxes_in_3_176_port, 
      boothmul_pipelined_i_muxes_in_3_175_port, 
      boothmul_pipelined_i_muxes_in_3_174_port, 
      boothmul_pipelined_i_muxes_in_3_173_port, 
      boothmul_pipelined_i_muxes_in_3_172_port, 
      boothmul_pipelined_i_muxes_in_3_171_port, 
      boothmul_pipelined_i_muxes_in_3_170_port, 
      boothmul_pipelined_i_muxes_in_3_169_port, 
      boothmul_pipelined_i_muxes_in_3_168_port, 
      boothmul_pipelined_i_muxes_in_3_167_port, 
      boothmul_pipelined_i_muxes_in_3_166_port, 
      boothmul_pipelined_i_muxes_in_3_165_port, 
      boothmul_pipelined_i_muxes_in_3_164_port, 
      boothmul_pipelined_i_muxes_in_3_163_port, 
      boothmul_pipelined_i_muxes_in_3_162_port, 
      boothmul_pipelined_i_muxes_in_3_161_port, 
      boothmul_pipelined_i_muxes_in_3_60_port, 
      boothmul_pipelined_i_muxes_in_3_59_port, 
      boothmul_pipelined_i_muxes_in_3_58_port, 
      boothmul_pipelined_i_muxes_in_3_57_port, 
      boothmul_pipelined_i_muxes_in_3_56_port, 
      boothmul_pipelined_i_muxes_in_3_55_port, 
      boothmul_pipelined_i_muxes_in_3_54_port, 
      boothmul_pipelined_i_muxes_in_3_53_port, 
      boothmul_pipelined_i_muxes_in_3_52_port, 
      boothmul_pipelined_i_muxes_in_3_51_port, 
      boothmul_pipelined_i_muxes_in_3_50_port, 
      boothmul_pipelined_i_muxes_in_3_49_port, 
      boothmul_pipelined_i_muxes_in_3_48_port, 
      boothmul_pipelined_i_muxes_in_3_47_port, 
      boothmul_pipelined_i_muxes_in_3_46_port, 
      boothmul_pipelined_i_sum_out_6_0_port, 
      boothmul_pipelined_i_sum_out_6_1_port, 
      boothmul_pipelined_i_sum_out_6_2_port, 
      boothmul_pipelined_i_sum_out_6_3_port, 
      boothmul_pipelined_i_sum_out_6_4_port, 
      boothmul_pipelined_i_sum_out_6_5_port, 
      boothmul_pipelined_i_sum_out_6_6_port, 
      boothmul_pipelined_i_sum_out_6_7_port, 
      boothmul_pipelined_i_sum_out_6_8_port, 
      boothmul_pipelined_i_sum_out_6_9_port, 
      boothmul_pipelined_i_sum_out_6_10_port, 
      boothmul_pipelined_i_sum_out_6_11_port, 
      boothmul_pipelined_i_sum_out_6_13_port, 
      boothmul_pipelined_i_sum_out_6_14_port, 
      boothmul_pipelined_i_sum_out_6_15_port, 
      boothmul_pipelined_i_sum_out_6_16_port, 
      boothmul_pipelined_i_sum_out_6_17_port, 
      boothmul_pipelined_i_sum_out_6_18_port, 
      boothmul_pipelined_i_sum_out_6_19_port, 
      boothmul_pipelined_i_sum_out_6_20_port, 
      boothmul_pipelined_i_sum_out_6_21_port, 
      boothmul_pipelined_i_sum_out_6_22_port, 
      boothmul_pipelined_i_sum_out_6_23_port, 
      boothmul_pipelined_i_sum_out_6_24_port, 
      boothmul_pipelined_i_sum_out_6_25_port, 
      boothmul_pipelined_i_sum_out_6_26_port, 
      boothmul_pipelined_i_sum_out_6_27_port, 
      boothmul_pipelined_i_sum_out_6_28_port, 
      boothmul_pipelined_i_sum_out_5_0_port, 
      boothmul_pipelined_i_sum_out_5_1_port, 
      boothmul_pipelined_i_sum_out_5_2_port, 
      boothmul_pipelined_i_sum_out_5_3_port, 
      boothmul_pipelined_i_sum_out_5_4_port, 
      boothmul_pipelined_i_sum_out_5_5_port, 
      boothmul_pipelined_i_sum_out_5_6_port, 
      boothmul_pipelined_i_sum_out_5_7_port, 
      boothmul_pipelined_i_sum_out_5_8_port, 
      boothmul_pipelined_i_sum_out_5_9_port, 
      boothmul_pipelined_i_sum_out_5_11_port, 
      boothmul_pipelined_i_sum_out_5_12_port, 
      boothmul_pipelined_i_sum_out_5_13_port, 
      boothmul_pipelined_i_sum_out_5_14_port, 
      boothmul_pipelined_i_sum_out_5_15_port, 
      boothmul_pipelined_i_sum_out_5_16_port, 
      boothmul_pipelined_i_sum_out_5_17_port, 
      boothmul_pipelined_i_sum_out_5_18_port, 
      boothmul_pipelined_i_sum_out_5_19_port, 
      boothmul_pipelined_i_sum_out_5_20_port, 
      boothmul_pipelined_i_sum_out_5_21_port, 
      boothmul_pipelined_i_sum_out_5_22_port, 
      boothmul_pipelined_i_sum_out_5_23_port, 
      boothmul_pipelined_i_sum_out_5_24_port, 
      boothmul_pipelined_i_sum_out_5_25_port, 
      boothmul_pipelined_i_sum_out_5_26_port, 
      boothmul_pipelined_i_sum_out_4_0_port, 
      boothmul_pipelined_i_sum_out_4_1_port, 
      boothmul_pipelined_i_sum_out_4_2_port, 
      boothmul_pipelined_i_sum_out_4_3_port, 
      boothmul_pipelined_i_sum_out_4_4_port, 
      boothmul_pipelined_i_sum_out_4_5_port, 
      boothmul_pipelined_i_sum_out_4_6_port, 
      boothmul_pipelined_i_sum_out_4_7_port, 
      boothmul_pipelined_i_sum_out_4_9_port, 
      boothmul_pipelined_i_sum_out_4_10_port, 
      boothmul_pipelined_i_sum_out_4_11_port, 
      boothmul_pipelined_i_sum_out_4_12_port, 
      boothmul_pipelined_i_sum_out_4_13_port, 
      boothmul_pipelined_i_sum_out_4_14_port, 
      boothmul_pipelined_i_sum_out_4_15_port, 
      boothmul_pipelined_i_sum_out_4_16_port, 
      boothmul_pipelined_i_sum_out_4_17_port, 
      boothmul_pipelined_i_sum_out_4_18_port, 
      boothmul_pipelined_i_sum_out_4_19_port, 
      boothmul_pipelined_i_sum_out_4_20_port, 
      boothmul_pipelined_i_sum_out_4_21_port, 
      boothmul_pipelined_i_sum_out_4_22_port, 
      boothmul_pipelined_i_sum_out_4_23_port, 
      boothmul_pipelined_i_sum_out_4_24_port, 
      boothmul_pipelined_i_sum_out_3_0_port, 
      boothmul_pipelined_i_sum_out_3_1_port, 
      boothmul_pipelined_i_sum_out_3_2_port, 
      boothmul_pipelined_i_sum_out_3_3_port, 
      boothmul_pipelined_i_sum_out_3_4_port, 
      boothmul_pipelined_i_sum_out_3_5_port, 
      boothmul_pipelined_i_sum_out_3_7_port, 
      boothmul_pipelined_i_sum_out_3_8_port, 
      boothmul_pipelined_i_sum_out_3_9_port, 
      boothmul_pipelined_i_sum_out_3_10_port, 
      boothmul_pipelined_i_sum_out_3_11_port, 
      boothmul_pipelined_i_sum_out_3_12_port, 
      boothmul_pipelined_i_sum_out_3_13_port, 
      boothmul_pipelined_i_sum_out_3_14_port, 
      boothmul_pipelined_i_sum_out_3_15_port, 
      boothmul_pipelined_i_sum_out_3_16_port, 
      boothmul_pipelined_i_sum_out_3_17_port, 
      boothmul_pipelined_i_sum_out_3_18_port, 
      boothmul_pipelined_i_sum_out_3_19_port, 
      boothmul_pipelined_i_sum_out_3_20_port, 
      boothmul_pipelined_i_sum_out_3_21_port, 
      boothmul_pipelined_i_sum_out_3_22_port, 
      boothmul_pipelined_i_sum_out_2_0_port, 
      boothmul_pipelined_i_sum_out_2_1_port, 
      boothmul_pipelined_i_sum_out_2_2_port, 
      boothmul_pipelined_i_sum_out_2_3_port, 
      boothmul_pipelined_i_sum_out_2_5_port, 
      boothmul_pipelined_i_sum_out_2_6_port, 
      boothmul_pipelined_i_sum_out_2_7_port, 
      boothmul_pipelined_i_sum_out_2_8_port, 
      boothmul_pipelined_i_sum_out_2_9_port, 
      boothmul_pipelined_i_sum_out_2_10_port, 
      boothmul_pipelined_i_sum_out_2_11_port, 
      boothmul_pipelined_i_sum_out_2_12_port, 
      boothmul_pipelined_i_sum_out_2_13_port, 
      boothmul_pipelined_i_sum_out_2_14_port, 
      boothmul_pipelined_i_sum_out_2_15_port, 
      boothmul_pipelined_i_sum_out_2_16_port, 
      boothmul_pipelined_i_sum_out_2_17_port, 
      boothmul_pipelined_i_sum_out_2_18_port, 
      boothmul_pipelined_i_sum_out_2_19_port, 
      boothmul_pipelined_i_sum_out_2_20_port, 
      boothmul_pipelined_i_sum_out_1_0_port, 
      boothmul_pipelined_i_sum_out_1_3_port, 
      boothmul_pipelined_i_sum_out_1_4_port, 
      boothmul_pipelined_i_sum_out_1_5_port, 
      boothmul_pipelined_i_sum_out_1_6_port, 
      boothmul_pipelined_i_sum_out_1_7_port, 
      boothmul_pipelined_i_sum_out_1_8_port, 
      boothmul_pipelined_i_sum_out_1_9_port, 
      boothmul_pipelined_i_sum_out_1_10_port, 
      boothmul_pipelined_i_sum_out_1_11_port, 
      boothmul_pipelined_i_sum_out_1_12_port, 
      boothmul_pipelined_i_sum_out_1_13_port, 
      boothmul_pipelined_i_sum_out_1_14_port, 
      boothmul_pipelined_i_sum_out_1_15_port, 
      boothmul_pipelined_i_sum_out_1_16_port, 
      boothmul_pipelined_i_sum_out_1_17_port, 
      boothmul_pipelined_i_sum_out_1_18_port, 
      boothmul_pipelined_i_sum_B_in_7_15_port, 
      boothmul_pipelined_i_sum_B_in_7_16_port, 
      boothmul_pipelined_i_sum_B_in_7_17_port, 
      boothmul_pipelined_i_sum_B_in_7_18_port, 
      boothmul_pipelined_i_sum_B_in_7_19_port, 
      boothmul_pipelined_i_sum_B_in_7_20_port, 
      boothmul_pipelined_i_sum_B_in_7_21_port, 
      boothmul_pipelined_i_sum_B_in_7_22_port, 
      boothmul_pipelined_i_sum_B_in_7_23_port, 
      boothmul_pipelined_i_sum_B_in_7_24_port, 
      boothmul_pipelined_i_sum_B_in_7_25_port, 
      boothmul_pipelined_i_sum_B_in_7_26_port, 
      boothmul_pipelined_i_sum_B_in_7_27_port, 
      boothmul_pipelined_i_sum_B_in_7_30_port, 
      boothmul_pipelined_i_sum_B_in_6_13_port, 
      boothmul_pipelined_i_sum_B_in_6_14_port, 
      boothmul_pipelined_i_sum_B_in_6_15_port, 
      boothmul_pipelined_i_sum_B_in_6_16_port, 
      boothmul_pipelined_i_sum_B_in_6_17_port, 
      boothmul_pipelined_i_sum_B_in_6_18_port, 
      boothmul_pipelined_i_sum_B_in_6_19_port, 
      boothmul_pipelined_i_sum_B_in_6_20_port, 
      boothmul_pipelined_i_sum_B_in_6_21_port, 
      boothmul_pipelined_i_sum_B_in_6_22_port, 
      boothmul_pipelined_i_sum_B_in_6_23_port, 
      boothmul_pipelined_i_sum_B_in_6_24_port, 
      boothmul_pipelined_i_sum_B_in_6_25_port, 
      boothmul_pipelined_i_sum_B_in_6_28_port, 
      boothmul_pipelined_i_sum_B_in_5_11_port, 
      boothmul_pipelined_i_sum_B_in_5_12_port, 
      boothmul_pipelined_i_sum_B_in_5_13_port, 
      boothmul_pipelined_i_sum_B_in_5_14_port, 
      boothmul_pipelined_i_sum_B_in_5_15_port, 
      boothmul_pipelined_i_sum_B_in_5_16_port, 
      boothmul_pipelined_i_sum_B_in_5_17_port, 
      boothmul_pipelined_i_sum_B_in_5_18_port, 
      boothmul_pipelined_i_sum_B_in_5_19_port, 
      boothmul_pipelined_i_sum_B_in_5_20_port, 
      boothmul_pipelined_i_sum_B_in_5_21_port, 
      boothmul_pipelined_i_sum_B_in_5_22_port, 
      boothmul_pipelined_i_sum_B_in_5_23_port, 
      boothmul_pipelined_i_sum_B_in_5_26_port, 
      boothmul_pipelined_i_sum_B_in_4_9_port, 
      boothmul_pipelined_i_sum_B_in_4_10_port, 
      boothmul_pipelined_i_sum_B_in_4_11_port, 
      boothmul_pipelined_i_sum_B_in_4_12_port, 
      boothmul_pipelined_i_sum_B_in_4_13_port, 
      boothmul_pipelined_i_sum_B_in_4_14_port, 
      boothmul_pipelined_i_sum_B_in_4_15_port, 
      boothmul_pipelined_i_sum_B_in_4_16_port, 
      boothmul_pipelined_i_sum_B_in_4_17_port, 
      boothmul_pipelined_i_sum_B_in_4_18_port, 
      boothmul_pipelined_i_sum_B_in_4_19_port, 
      boothmul_pipelined_i_sum_B_in_4_20_port, 
      boothmul_pipelined_i_sum_B_in_4_21_port, 
      boothmul_pipelined_i_sum_B_in_4_24_port, 
      boothmul_pipelined_i_sum_B_in_3_7_port, 
      boothmul_pipelined_i_sum_B_in_3_8_port, 
      boothmul_pipelined_i_sum_B_in_3_9_port, 
      boothmul_pipelined_i_sum_B_in_3_10_port, 
      boothmul_pipelined_i_sum_B_in_3_11_port, 
      boothmul_pipelined_i_sum_B_in_3_12_port, 
      boothmul_pipelined_i_sum_B_in_3_13_port, 
      boothmul_pipelined_i_sum_B_in_3_14_port, 
      boothmul_pipelined_i_sum_B_in_3_15_port, 
      boothmul_pipelined_i_sum_B_in_3_16_port, 
      boothmul_pipelined_i_sum_B_in_3_17_port, 
      boothmul_pipelined_i_sum_B_in_3_18_port, 
      boothmul_pipelined_i_sum_B_in_3_19_port, 
      boothmul_pipelined_i_sum_B_in_3_22_port, 
      boothmul_pipelined_i_sum_B_in_2_5_port, 
      boothmul_pipelined_i_sum_B_in_2_6_port, 
      boothmul_pipelined_i_sum_B_in_2_7_port, 
      boothmul_pipelined_i_sum_B_in_2_8_port, 
      boothmul_pipelined_i_sum_B_in_2_9_port, 
      boothmul_pipelined_i_sum_B_in_2_10_port, 
      boothmul_pipelined_i_sum_B_in_2_11_port, 
      boothmul_pipelined_i_sum_B_in_2_12_port, 
      boothmul_pipelined_i_sum_B_in_2_13_port, 
      boothmul_pipelined_i_sum_B_in_2_14_port, 
      boothmul_pipelined_i_sum_B_in_2_15_port, 
      boothmul_pipelined_i_sum_B_in_2_16_port, 
      boothmul_pipelined_i_sum_B_in_2_17_port, 
      boothmul_pipelined_i_sum_B_in_2_20_port, 
      boothmul_pipelined_i_sum_B_in_1_15_port, 
      boothmul_pipelined_i_sum_B_in_1_18_port, 
      boothmul_pipelined_i_mux_out_7_15_port, 
      boothmul_pipelined_i_mux_out_7_16_port, 
      boothmul_pipelined_i_mux_out_7_17_port, 
      boothmul_pipelined_i_mux_out_7_18_port, 
      boothmul_pipelined_i_mux_out_7_19_port, 
      boothmul_pipelined_i_mux_out_7_20_port, 
      boothmul_pipelined_i_mux_out_7_21_port, 
      boothmul_pipelined_i_mux_out_7_22_port, 
      boothmul_pipelined_i_mux_out_7_23_port, 
      boothmul_pipelined_i_mux_out_7_24_port, 
      boothmul_pipelined_i_mux_out_7_25_port, 
      boothmul_pipelined_i_mux_out_7_26_port, 
      boothmul_pipelined_i_mux_out_7_27_port, 
      boothmul_pipelined_i_mux_out_7_28_port, 
      boothmul_pipelined_i_mux_out_7_29_port, 
      boothmul_pipelined_i_mux_out_7_30_port, 
      boothmul_pipelined_i_mux_out_6_13_port, 
      boothmul_pipelined_i_mux_out_6_14_port, 
      boothmul_pipelined_i_mux_out_6_15_port, 
      boothmul_pipelined_i_mux_out_6_16_port, 
      boothmul_pipelined_i_mux_out_6_17_port, 
      boothmul_pipelined_i_mux_out_6_18_port, 
      boothmul_pipelined_i_mux_out_6_19_port, 
      boothmul_pipelined_i_mux_out_6_20_port, 
      boothmul_pipelined_i_mux_out_6_21_port, 
      boothmul_pipelined_i_mux_out_6_22_port, 
      boothmul_pipelined_i_mux_out_6_23_port, 
      boothmul_pipelined_i_mux_out_6_24_port, 
      boothmul_pipelined_i_mux_out_6_25_port, 
      boothmul_pipelined_i_mux_out_6_26_port, 
      boothmul_pipelined_i_mux_out_6_27_port, 
      boothmul_pipelined_i_mux_out_5_11_port, 
      boothmul_pipelined_i_mux_out_5_12_port, 
      boothmul_pipelined_i_mux_out_5_13_port, 
      boothmul_pipelined_i_mux_out_5_14_port, 
      boothmul_pipelined_i_mux_out_5_15_port, 
      boothmul_pipelined_i_mux_out_5_16_port, 
      boothmul_pipelined_i_mux_out_5_17_port, 
      boothmul_pipelined_i_mux_out_5_18_port, 
      boothmul_pipelined_i_mux_out_5_19_port, 
      boothmul_pipelined_i_mux_out_5_20_port, 
      boothmul_pipelined_i_mux_out_5_21_port, 
      boothmul_pipelined_i_mux_out_5_22_port, 
      boothmul_pipelined_i_mux_out_5_23_port, 
      boothmul_pipelined_i_mux_out_5_24_port, 
      boothmul_pipelined_i_mux_out_5_25_port, 
      boothmul_pipelined_i_mux_out_4_9_port, 
      boothmul_pipelined_i_mux_out_4_10_port, 
      boothmul_pipelined_i_mux_out_4_11_port, 
      boothmul_pipelined_i_mux_out_4_12_port, 
      boothmul_pipelined_i_mux_out_4_13_port, 
      boothmul_pipelined_i_mux_out_4_14_port, 
      boothmul_pipelined_i_mux_out_4_15_port, 
      boothmul_pipelined_i_mux_out_4_16_port, 
      boothmul_pipelined_i_mux_out_4_17_port, 
      boothmul_pipelined_i_mux_out_4_18_port, 
      boothmul_pipelined_i_mux_out_4_19_port, 
      boothmul_pipelined_i_mux_out_4_20_port, 
      boothmul_pipelined_i_mux_out_4_21_port, 
      boothmul_pipelined_i_mux_out_4_22_port, 
      boothmul_pipelined_i_mux_out_4_23_port, 
      boothmul_pipelined_i_mux_out_3_7_port, 
      boothmul_pipelined_i_mux_out_3_8_port, 
      boothmul_pipelined_i_mux_out_3_9_port, 
      boothmul_pipelined_i_mux_out_3_10_port, 
      boothmul_pipelined_i_mux_out_3_11_port, 
      boothmul_pipelined_i_mux_out_3_12_port, 
      boothmul_pipelined_i_mux_out_3_13_port, 
      boothmul_pipelined_i_mux_out_3_14_port, 
      boothmul_pipelined_i_mux_out_3_15_port, 
      boothmul_pipelined_i_mux_out_3_16_port, 
      boothmul_pipelined_i_mux_out_3_17_port, 
      boothmul_pipelined_i_mux_out_3_18_port, 
      boothmul_pipelined_i_mux_out_3_19_port, 
      boothmul_pipelined_i_mux_out_3_20_port, 
      boothmul_pipelined_i_mux_out_3_21_port, 
      boothmul_pipelined_i_mux_out_2_5_port, 
      boothmul_pipelined_i_mux_out_2_6_port, 
      boothmul_pipelined_i_mux_out_2_7_port, 
      boothmul_pipelined_i_mux_out_2_8_port, 
      boothmul_pipelined_i_mux_out_2_9_port, 
      boothmul_pipelined_i_mux_out_2_10_port, 
      boothmul_pipelined_i_mux_out_2_11_port, 
      boothmul_pipelined_i_mux_out_2_12_port, 
      boothmul_pipelined_i_mux_out_2_13_port, 
      boothmul_pipelined_i_mux_out_2_14_port, 
      boothmul_pipelined_i_mux_out_2_15_port, 
      boothmul_pipelined_i_mux_out_2_16_port, 
      boothmul_pipelined_i_mux_out_2_17_port, 
      boothmul_pipelined_i_mux_out_2_18_port, 
      boothmul_pipelined_i_mux_out_2_19_port, 
      boothmul_pipelined_i_mux_out_2_20_port, 
      boothmul_pipelined_i_mux_out_1_3_port, 
      boothmul_pipelined_i_mux_out_1_4_port, 
      boothmul_pipelined_i_mux_out_1_5_port, 
      boothmul_pipelined_i_mux_out_1_6_port, 
      boothmul_pipelined_i_mux_out_1_7_port, 
      boothmul_pipelined_i_mux_out_1_8_port, 
      boothmul_pipelined_i_mux_out_1_9_port, 
      boothmul_pipelined_i_mux_out_1_10_port, 
      boothmul_pipelined_i_mux_out_1_11_port, 
      boothmul_pipelined_i_mux_out_1_12_port, 
      boothmul_pipelined_i_mux_out_1_13_port, 
      boothmul_pipelined_i_mux_out_1_14_port, 
      boothmul_pipelined_i_mux_out_1_15_port, 
      boothmul_pipelined_i_mux_out_1_16_port, 
      boothmul_pipelined_i_mux_out_1_17_port, 
      boothmul_pipelined_i_mux_out_1_18_port, 
      boothmul_pipelined_i_encoder_out_0_0_port, 
      boothmul_pipelined_i_multiplicand_pip_7_13_port, 
      boothmul_pipelined_i_multiplicand_pip_7_14_port, 
      boothmul_pipelined_i_multiplicand_pip_7_15_port, 
      boothmul_pipelined_i_multiplicand_pip_6_11_port, 
      boothmul_pipelined_i_multiplicand_pip_6_12_port, 
      boothmul_pipelined_i_multiplicand_pip_6_13_port, 
      boothmul_pipelined_i_multiplicand_pip_6_14_port, 
      boothmul_pipelined_i_multiplicand_pip_6_15_port, 
      boothmul_pipelined_i_multiplicand_pip_5_9_port, 
      boothmul_pipelined_i_multiplicand_pip_5_10_port, 
      boothmul_pipelined_i_multiplicand_pip_5_11_port, 
      boothmul_pipelined_i_multiplicand_pip_5_12_port, 
      boothmul_pipelined_i_multiplicand_pip_5_13_port, 
      boothmul_pipelined_i_multiplicand_pip_5_14_port, 
      boothmul_pipelined_i_multiplicand_pip_5_15_port, 
      boothmul_pipelined_i_multiplicand_pip_4_7_port, 
      boothmul_pipelined_i_multiplicand_pip_4_8_port, 
      boothmul_pipelined_i_multiplicand_pip_4_9_port, 
      boothmul_pipelined_i_multiplicand_pip_4_10_port, 
      boothmul_pipelined_i_multiplicand_pip_4_11_port, 
      boothmul_pipelined_i_multiplicand_pip_4_12_port, 
      boothmul_pipelined_i_multiplicand_pip_4_13_port, 
      boothmul_pipelined_i_multiplicand_pip_4_14_port, 
      boothmul_pipelined_i_multiplicand_pip_4_15_port, 
      boothmul_pipelined_i_multiplicand_pip_3_5_port, 
      boothmul_pipelined_i_multiplicand_pip_3_6_port, 
      boothmul_pipelined_i_multiplicand_pip_3_7_port, 
      boothmul_pipelined_i_multiplicand_pip_3_8_port, 
      boothmul_pipelined_i_multiplicand_pip_3_9_port, 
      boothmul_pipelined_i_multiplicand_pip_3_10_port, 
      boothmul_pipelined_i_multiplicand_pip_3_11_port, 
      boothmul_pipelined_i_multiplicand_pip_3_12_port, 
      boothmul_pipelined_i_multiplicand_pip_3_13_port, 
      boothmul_pipelined_i_multiplicand_pip_3_14_port, 
      boothmul_pipelined_i_multiplicand_pip_3_15_port, 
      boothmul_pipelined_i_multiplicand_pip_2_3_port, 
      boothmul_pipelined_i_multiplicand_pip_2_4_port, 
      boothmul_pipelined_i_multiplicand_pip_2_5_port, 
      boothmul_pipelined_i_multiplicand_pip_2_6_port, 
      boothmul_pipelined_i_multiplicand_pip_2_7_port, 
      boothmul_pipelined_i_multiplicand_pip_2_8_port, 
      boothmul_pipelined_i_multiplicand_pip_2_9_port, 
      boothmul_pipelined_i_multiplicand_pip_2_10_port, 
      boothmul_pipelined_i_multiplicand_pip_2_11_port, 
      boothmul_pipelined_i_multiplicand_pip_2_12_port, 
      boothmul_pipelined_i_multiplicand_pip_2_13_port, 
      boothmul_pipelined_i_multiplicand_pip_2_14_port, 
      boothmul_pipelined_i_multiplicand_pip_2_15_port, 
      boothmul_pipelined_i_muxes_in_0_119_port, 
      boothmul_pipelined_i_muxes_in_0_116_port, 
      boothmul_pipelined_i_muxes_in_0_115_port, 
      boothmul_pipelined_i_muxes_in_0_114_port, 
      boothmul_pipelined_i_muxes_in_0_113_port, 
      boothmul_pipelined_i_muxes_in_0_112_port, 
      boothmul_pipelined_i_muxes_in_0_111_port, 
      boothmul_pipelined_i_muxes_in_0_110_port, 
      boothmul_pipelined_i_muxes_in_0_109_port, 
      boothmul_pipelined_i_muxes_in_0_108_port, 
      boothmul_pipelined_i_muxes_in_0_107_port, 
      boothmul_pipelined_i_muxes_in_0_106_port, 
      boothmul_pipelined_i_muxes_in_0_105_port, 
      boothmul_pipelined_i_muxes_in_0_104_port, 
      boothmul_pipelined_i_muxes_in_0_103_port, 
      boothmul_pipelined_i_muxes_in_0_102_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
      boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
      boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, n3076, 
      n3077, n3078, n3079, n3080, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n1995, n1996, 
      n1997, n5121, n5122, n5123, n5124, n5126, n5127, n5128, n5129, n5130, 
      n5131, n5132, n5133, n5134, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n5141, n5142, n5143, n5144, n5145, 
      n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, 
      n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, 
      n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, 
      n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, 
      n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, 
      n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, 
      n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, 
      n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, 
      n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, 
      n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, 
      n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, 
      n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, 
      n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, 
      n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, 
      n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, 
      n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, 
      n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, 
      n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, 
      n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, 
      n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, 
      n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, 
      n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, 
      n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, 
      n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, 
      n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, 
      n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, 
      n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, 
      n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, 
      n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, 
      n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, 
      n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, 
      n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, 
      n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, 
      n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, 
      n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, 
      n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, 
      n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, 
      n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, 
      n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, 
      n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, 
      n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, 
      n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, 
      n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, 
      n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, 
      n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, 
      n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, 
      n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, 
      n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, 
      n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, 
      n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, 
      n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, 
      n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, 
      n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, 
      n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, 
      n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, 
      n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, 
      n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, 
      n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, 
      n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, 
      n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, 
      n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, 
      n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, 
      n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, 
      n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, 
      n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, 
      n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, 
      n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, 
      n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, 
      n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, 
      n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, 
      n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, 
      n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, 
      n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, 
      n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, 
      n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, 
      n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, 
      n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, 
      n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, 
      n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, 
      n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, 
      n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, 
      n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, 
      n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, 
      n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, 
      n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, 
      n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, 
      n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, 
      n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, 
      n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, 
      n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, 
      n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, 
      n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, 
      n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, 
      n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, 
      n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, 
      n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, 
      n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, 
      n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, 
      n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, 
      n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, 
      n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, 
      n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, 
      n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, 
      n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, 
      n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, 
      n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, 
      n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, 
      n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, 
      n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, 
      n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, 
      n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, 
      n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, 
      n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, 
      n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, 
      n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, 
      n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, 
      n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
      n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, 
      n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, 
      n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, 
      n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
      n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, 
      n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, 
      n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, 
      n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, 
      n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, 
      n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, 
      n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, 
      n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, 
      n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, 
      n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, 
      n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, 
      n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, 
      n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, 
      n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, 
      n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, 
      n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, 
      n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, 
      n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, 
      n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, 
      n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, 
      n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, 
      n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, 
      n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, 
      n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, 
      n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, 
      n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, 
      n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, 
      n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, 
      n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, 
      n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, 
      n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, 
      n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, 
      n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, 
      n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, 
      n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, 
      n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, 
      n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, 
      n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, 
      n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, 
      n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, 
      n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, 
      n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, 
      n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, 
      n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
      n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, 
      n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, 
      n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, 
      n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, 
      n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, 
      n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, 
      n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, 
      n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, 
      n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, 
      n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
      n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, 
      n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, 
      n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, 
      n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
      n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, 
      n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, 
      n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, 
      n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
      n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, 
      n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, 
      n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, 
      n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, 
      n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, 
      n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, 
      n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, 
      n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, 
      n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, 
      n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, 
      n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, 
      n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, 
      n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, 
      n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, 
      n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, 
      n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, 
      n7166, n7167, n7168, n7169, n_1004, n_1005, n_1006, n_1007, n_1008, 
      n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, 
      n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, 
      n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, 
      n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, 
      n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, 
      n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, 
      n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, 
      n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, 
      n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, 
      n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, 
      n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, 
      n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, 
      n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, 
      n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, 
      n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, 
      n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, 
      n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, 
      n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, 
      n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, 
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, 
      n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, 
      n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, 
      n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, 
      n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, 
      n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, 
      n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, 
      n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, 
      n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, 
      n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, 
      n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, 
      n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, 
      n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, 
      n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, 
      n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, 
      n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, 
      n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, 
      n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348 : std_logic;

begin
   
   DATA2_I_reg_28_inst : DLL_X1 port map( D => N2545, GN => n7166, Q => 
                           DATA2_I_28_port);
   DATA2_I_reg_27_inst : DLL_X1 port map( D => N2544, GN => n1992, Q => 
                           DATA2_I_27_port);
   DATA2_I_reg_26_inst : DLL_X1 port map( D => N2543, GN => n1992, Q => 
                           DATA2_I_26_port);
   DATA2_I_reg_25_inst : DLL_X1 port map( D => N2542, GN => n1992, Q => 
                           DATA2_I_25_port);
   DATA2_I_reg_24_inst : DLL_X1 port map( D => N2541, GN => n1992, Q => 
                           DATA2_I_24_port);
   DATA2_I_reg_23_inst : DLL_X1 port map( D => N2540, GN => n1992, Q => 
                           DATA2_I_23_port);
   DATA2_I_reg_22_inst : DLL_X1 port map( D => N2539, GN => n7166, Q => 
                           DATA2_I_22_port);
   DATA2_I_reg_21_inst : DLL_X1 port map( D => N2538, GN => n7166, Q => 
                           DATA2_I_21_port);
   DATA2_I_reg_20_inst : DLL_X1 port map( D => N2537, GN => n1992, Q => 
                           DATA2_I_20_port);
   DATA2_I_reg_19_inst : DLL_X1 port map( D => N2536, GN => n7166, Q => 
                           DATA2_I_19_port);
   DATA2_I_reg_18_inst : DLL_X1 port map( D => N2535, GN => n1992, Q => 
                           DATA2_I_18_port);
   DATA2_I_reg_17_inst : DLL_X1 port map( D => N2534, GN => n1992, Q => 
                           DATA2_I_17_port);
   DATA2_I_reg_16_inst : DLL_X1 port map( D => N2533, GN => n1992, Q => 
                           DATA2_I_16_port);
   DATA2_I_reg_15_inst : DLL_X1 port map( D => N2532, GN => n7166, Q => 
                           DATA2_I_15_port);
   DATA2_I_reg_14_inst : DLL_X1 port map( D => N2531, GN => n1992, Q => 
                           DATA2_I_14_port);
   DATA2_I_reg_13_inst : DLL_X1 port map( D => N2530, GN => n7166, Q => 
                           DATA2_I_13_port);
   DATA2_I_reg_12_inst : DLL_X1 port map( D => N2529, GN => n1992, Q => 
                           DATA2_I_12_port);
   DATA2_I_reg_11_inst : DLL_X1 port map( D => N2528, GN => n7166, Q => 
                           DATA2_I_11_port);
   DATA2_I_reg_10_inst : DLL_X1 port map( D => N2527, GN => n1992, Q => 
                           DATA2_I_10_port);
   DATA2_I_reg_9_inst : DLL_X1 port map( D => N2526, GN => n7166, Q => 
                           DATA2_I_9_port);
   DATA2_I_reg_8_inst : DLL_X1 port map( D => N2525, GN => n7166, Q => 
                           DATA2_I_8_port);
   DATA2_I_reg_7_inst : DLL_X1 port map( D => N2524, GN => n1992, Q => 
                           DATA2_I_7_port);
   DATA2_I_reg_6_inst : DLL_X1 port map( D => N2523, GN => n7166, Q => 
                           DATA2_I_6_port);
   DATA2_I_reg_5_inst : DLL_X1 port map( D => N2522, GN => n7166, Q => 
                           DATA2_I_5_port);
   DATA2_I_reg_4_inst : DLL_X1 port map( D => N2521, GN => n7166, Q => 
                           DATA2_I_4_port);
   DATA2_I_reg_3_inst : DLL_X1 port map( D => N2520, GN => n1992, Q => 
                           DATA2_I_3_port);
   DATA2_I_reg_2_inst : DLL_X1 port map( D => N2519, GN => n1992, Q => 
                           DATA2_I_2_port);
   DATA2_I_reg_1_inst : DLL_X1 port map( D => N2518, GN => n7166, Q => 
                           DATA2_I_1_port);
   DATA2_I_reg_0_inst : DLL_X1 port map( D => N2517, GN => n7166, Q => 
                           DATA2_I_0_port);
   data1_mul_reg_15_inst : DLL_X1 port map( D => DATA1(15), GN => n553, Q => 
                           data1_mul_15_port);
   data1_mul_reg_14_inst : DLL_X1 port map( D => n7169, GN => n553, Q => 
                           data1_mul_14_port);
   data1_mul_reg_13_inst : DLL_X1 port map( D => DATA1(13), GN => n553, Q => 
                           data1_mul_13_port);
   data1_mul_reg_12_inst : DLL_X1 port map( D => n7168, GN => n553, Q => 
                           data1_mul_12_port);
   data1_mul_reg_11_inst : DLL_X1 port map( D => DATA1(11), GN => n553, Q => 
                           data1_mul_11_port);
   data1_mul_reg_10_inst : DLL_X1 port map( D => n7167, GN => n553, Q => 
                           data1_mul_10_port);
   data1_mul_reg_9_inst : DLL_X1 port map( D => DATA1(9), GN => n553, Q => 
                           data1_mul_9_port);
   data1_mul_reg_8_inst : DLL_X1 port map( D => DATA1(8), GN => n553, Q => 
                           data1_mul_8_port);
   data1_mul_reg_7_inst : DLL_X1 port map( D => DATA1(7), GN => n553, Q => 
                           data1_mul_7_port);
   data1_mul_reg_6_inst : DLL_X1 port map( D => DATA1(6), GN => n553, Q => 
                           data1_mul_6_port);
   data1_mul_reg_5_inst : DLL_X1 port map( D => DATA1(5), GN => n553, Q => 
                           data1_mul_5_port);
   data1_mul_reg_4_inst : DLL_X1 port map( D => DATA1(4), GN => n553, Q => 
                           data1_mul_4_port);
   data1_mul_reg_3_inst : DLL_X1 port map( D => DATA1(3), GN => n553, Q => 
                           data1_mul_3_port);
   data1_mul_reg_2_inst : DLL_X1 port map( D => DATA1(2), GN => n553, Q => 
                           data1_mul_2_port);
   data1_mul_reg_1_inst : DLL_X1 port map( D => DATA1(1), GN => n553, Q => 
                           data1_mul_1_port);
   data1_mul_reg_0_inst : DLL_X1 port map( D => DATA1(0), GN => n553, Q => 
                           data1_mul_0_port);
   data2_mul_reg_15_inst : DLL_X1 port map( D => DATA2(15), GN => n553, Q => 
                           data2_mul_15_port);
   data2_mul_reg_14_inst : DLL_X1 port map( D => DATA2(14), GN => n553, Q => 
                           data2_mul_14_port);
   data2_mul_reg_13_inst : DLL_X1 port map( D => DATA2(13), GN => n553, Q => 
                           data2_mul_13_port);
   data2_mul_reg_12_inst : DLL_X1 port map( D => DATA2(12), GN => n553, Q => 
                           data2_mul_12_port);
   data2_mul_reg_11_inst : DLL_X1 port map( D => DATA2(11), GN => n553, Q => 
                           data2_mul_11_port);
   data2_mul_reg_10_inst : DLL_X1 port map( D => DATA2(10), GN => n553, Q => 
                           data2_mul_10_port);
   data2_mul_reg_9_inst : DLL_X1 port map( D => DATA2(9), GN => n553, Q => 
                           data2_mul_9_port);
   data2_mul_reg_8_inst : DLL_X1 port map( D => DATA2(8), GN => n553, Q => 
                           data2_mul_8_port);
   data2_mul_reg_7_inst : DLL_X1 port map( D => DATA2(7), GN => n553, Q => 
                           data2_mul_7_port);
   data2_mul_reg_6_inst : DLL_X1 port map( D => DATA2(6), GN => n553, Q => 
                           data2_mul_6_port);
   data2_mul_reg_5_inst : DLL_X1 port map( D => DATA2(5), GN => n553, Q => 
                           data2_mul_5_port);
   data2_mul_reg_4_inst : DLL_X1 port map( D => DATA2(4), GN => n553, Q => 
                           data2_mul_4_port);
   data2_mul_reg_3_inst : DLL_X1 port map( D => DATA2(3), GN => n553, Q => 
                           data2_mul_3_port);
   data2_mul_reg_2_inst : DLL_X1 port map( D => DATA2(2), GN => n553, Q => 
                           data2_mul_2_port);
   data2_mul_reg_0_inst : DLL_X1 port map( D => DATA2(0), GN => n553, Q => 
                           boothmul_pipelined_i_encoder_out_0_0_port);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, CK 
                           => clk, RN => n5146, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, QN 
                           => n7165);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, CK 
                           => clk, RN => n5147, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_14_port, QN 
                           => n_1004);
   boothmul_pipelined_i_pip_del_reg_i_7_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, QN 
                           => n_1005);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, CK 
                           => clk, RN => n5154, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_15_port, QN 
                           => n_1006);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, CK 
                           => clk, RN => n5143, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_14_port, QN 
                           => n_1007);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, CK 
                           => clk, RN => n5145, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_13_port, QN 
                           => n3080);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, CK 
                           => clk, RN => n5142, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, QN 
                           => n_1008);
   boothmul_pipelined_i_pip_del_reg_i_6_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, CK 
                           => clk, RN => n5145, Q => 
                           boothmul_pipelined_i_multiplicand_pip_6_11_port, QN 
                           => n_1009);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_15_port, QN 
                           => n_1010);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, CK 
                           => clk, RN => n5142, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_14_port, QN 
                           => n_1011);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, CK 
                           => clk, RN => n5152, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_13_port, QN 
                           => n_1012);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, CK 
                           => clk, RN => n5150, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_12_port, QN 
                           => n_1013);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, CK 
                           => clk, RN => n5147, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_11_port, QN 
                           => n3079);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, CK 
                           => clk, RN => n5148, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, QN 
                           => n_1014);
   boothmul_pipelined_i_pip_del_reg_i_5_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, CK 
                           => clk, RN => n5155, Q => 
                           boothmul_pipelined_i_multiplicand_pip_5_9_port, QN 
                           => n_1015);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, CK 
                           => clk, RN => n5143, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_15_port, QN 
                           => n_1016);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, CK 
                           => clk, RN => n5151, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_14_port, QN 
                           => n_1017);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, CK 
                           => clk, RN => n5152, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_13_port, QN 
                           => n_1018);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, CK 
                           => clk, RN => n5141, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_12_port, QN 
                           => n_1019);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, CK 
                           => clk, RN => n5153, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_11_port, QN 
                           => n_1020);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, CK 
                           => clk, RN => n5145, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_10_port, QN 
                           => n_1021);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, CK 
                           => clk, RN => n5153, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_9_port, QN 
                           => n3078);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, QN 
                           => n_1022);
   boothmul_pipelined_i_pip_del_reg_i_4_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, CK 
                           => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_4_7_port, QN 
                           => n_1023);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, CK 
                           => clk, RN => n5152, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_15_port, QN 
                           => n_1024);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, CK 
                           => clk, RN => n5151, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_14_port, QN 
                           => n_1025);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, CK 
                           => clk, RN => n5147, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_13_port, QN 
                           => n_1026);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, CK 
                           => clk, RN => n5151, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_12_port, QN 
                           => n_1027);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, CK 
                           => clk, RN => n5146, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_11_port, QN 
                           => n_1028);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, CK 
                           => clk, RN => n5145, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_10_port, QN 
                           => n_1029);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, CK 
                           => clk, RN => n5154, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_9_port, QN 
                           => n_1030);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, CK 
                           => clk, RN => n5152, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_8_port, QN 
                           => n_1031);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, CK 
                           => clk, RN => n5150, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, QN 
                           => n3082);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, CK 
                           => clk, RN => n5144, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, QN 
                           => n_1032);
   boothmul_pipelined_i_pip_del_reg_i_3_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, CK 
                           => clk, RN => n5149, Q => 
                           boothmul_pipelined_i_multiplicand_pip_3_5_port, QN 
                           => n_1033);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_15_port, CK => clk, RN => n5143, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_15_port, QN 
                           => n_1034);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_14_port, CK => clk, RN => n5148, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_14_port, QN 
                           => n_1035);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_13_port, CK => clk, RN => n5155, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_13_port, QN 
                           => n_1036);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_12_port, CK => clk, RN => n5144, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_12_port, QN 
                           => n_1037);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_11_port, CK => clk, RN => n5155, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_11_port, QN 
                           => n_1038);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_10_port, CK => clk, RN => n5146, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_10_port, QN 
                           => n_1039);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_9_port, CK => clk, RN => n5148, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_9_port, QN 
                           => n_1040);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_8_port, CK => clk, RN => n5148, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_8_port, QN 
                           => n_1041);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_7_port, CK => clk, RN => n5152, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_7_port, QN 
                           => n_1042);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_6_port, CK => clk, RN => n5142, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_6_port, QN 
                           => n_1043);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_5_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, QN 
                           => n3076);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_4_port, CK => clk, RN => n5155, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, QN 
                           => n_1044);
   boothmul_pipelined_i_pip_del_reg_i_2_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           data2_mul_3_port, CK => clk, RN => n5148, Q => 
                           boothmul_pipelined_i_multiplicand_pip_2_3_port, QN 
                           => n_1045);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_28_port, CK => clk
                           , RN => n5155, Q => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, QN => 
                           n_1046);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_27_port, CK => clk
                           , RN => n5144, Q => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, QN => 
                           n_1047);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_26_port, CK => clk
                           , RN => n5144, Q => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, QN => 
                           n_1048);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_25_port, CK => clk
                           , RN => n5150, Q => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, QN => 
                           n_1049);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_24_port, CK => clk
                           , RN => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, QN => 
                           n_1050);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_23_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, QN => 
                           n_1051);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_22_port, CK => clk
                           , RN => n5150, Q => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, QN => 
                           n_1052);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_21_port, CK => clk
                           , RN => n5143, Q => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, QN => 
                           n_1053);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_20_port, CK => clk
                           , RN => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, QN => 
                           n_1054);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_19_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, QN => 
                           n_1055);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_18_port, CK => clk
                           , RN => n5154, Q => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, QN => 
                           n_1056);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_17_port, CK => clk
                           , RN => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, QN => 
                           n_1057);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_16_port, CK => clk
                           , RN => n5147, Q => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, QN => 
                           n_1058);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_15_port, CK => clk
                           , RN => n5145, Q => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, QN => 
                           n_1059);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_14_port, CK => clk
                           , RN => n5146, Q => n_1060, QN => n5126);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_13_port, CK => clk
                           , RN => n5152, Q => dataout_mul_13_port, QN => 
                           n_1061);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => n3095, CK => clk, RN => n5142, Q => 
                           dataout_mul_12_port, QN => n_1062);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_11_port, CK => clk
                           , RN => n5150, Q => dataout_mul_11_port, QN => 
                           n_1063);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_6_10_port, CK => clk
                           , RN => n5152, Q => dataout_mul_10_port, QN => 
                           n_1064);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_9_port, CK => clk, RN
                           => n5146, Q => dataout_mul_9_port, QN => n_1065);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_8_port, CK => clk, RN
                           => n5155, Q => dataout_mul_8_port, QN => n_1066);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_7_port, CK => clk, RN
                           => n5155, Q => dataout_mul_7_port, QN => n_1067);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_6_port, CK => clk, RN
                           => n5153, Q => dataout_mul_6_port, QN => n_1068);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_5_port, CK => clk, RN
                           => n5142, Q => dataout_mul_5_port, QN => n_1069);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_4_port, CK => clk, RN
                           => n5145, Q => dataout_mul_4_port, QN => n_1070);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_3_port, CK => clk, RN
                           => n5151, Q => dataout_mul_3_port, QN => n_1071);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_2_port, CK => clk, RN
                           => n5142, Q => dataout_mul_2_port, QN => n_1072);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_1_port, CK => clk, RN
                           => n5151, Q => dataout_mul_1_port, QN => n_1073);
   boothmul_pipelined_i_pip_del_reg_addi_6_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_6_0_port, CK => clk, RN
                           => n5153, Q => dataout_mul_0_port, QN => n_1074);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_58_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_7_62_port, QN => 
                           n_1075);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_59_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_7_63_port, QN => 
                           n_1076);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_60_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_7_64_port, QN => 
                           n_1077);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_61_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_7_65_port, QN => 
                           n_1078);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_62_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_7_66_port, QN => 
                           n_1079);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_63_port, CK => 
                           clk, RN => n5142, Q => 
                           boothmul_pipelined_i_muxes_in_7_67_port, QN => 
                           n_1080);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_64_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_7_68_port, QN => 
                           n_1081);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_65_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_7_69_port, QN => 
                           n_1082);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_66_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_7_70_port, QN => 
                           n_1083);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_67_port, CK => 
                           clk, RN => n5143, Q => 
                           boothmul_pipelined_i_muxes_in_7_71_port, QN => 
                           n_1084);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_68_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_7_72_port, QN => 
                           n_1085);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_69_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_7_73_port, QN => 
                           n_1086);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_178_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_70_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_7_74_port, QN => 
                           n_1087);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_177_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_71_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_7_75_port, QN => 
                           n_1088);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_176_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_72_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_7_76_port, QN => 
                           n_1089);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_203_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_7_217_port, QN => 
                           n_1090);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_204_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_7_218_port, QN => 
                           n_1091);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_43_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_205_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_7_219_port, QN => 
                           n_1092);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_42_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_206_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_7_220_port, QN => 
                           n_1093);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_41_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_207_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_7_221_port, QN => 
                           n_1094);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_40_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_208_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_7_222_port, QN => 
                           n_1095);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_39_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_209_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_7_223_port, QN => 
                           n_1096);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_38_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_210_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_7_224_port, QN => 
                           n_1097);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_37_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_211_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_7_225_port, QN => 
                           n_1098);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_36_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_212_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_7_226_port, QN => 
                           n_1099);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_35_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_213_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_7_227_port, QN => 
                           n_1100);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_34_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_214_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_7_228_port, QN => 
                           n_1101);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_33_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_215_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_7_229_port, QN => 
                           n_1102);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_216_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_7_230_port, QN => 
                           n_1103);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_217_port, CK => 
                           clk, RN => n5152, Q => 
                           boothmul_pipelined_i_muxes_in_7_231_port, QN => 
                           n_1104);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_218_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_7_232_port, QN => 
                           n_1105);
   boothmul_pipelined_i_pip_del_reg_muxi_6_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_6_73_port, CK => 
                           clk, RN => n5147, Q => n_1106, QN => n5134);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_26_port, CK => clk
                           , RN => n5152, Q => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, QN => 
                           n_1107);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_25_port, CK => clk
                           , RN => n5142, Q => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, QN => 
                           n_1108);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_24_port, CK => clk
                           , RN => n5151, Q => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, QN => 
                           n_1109);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_23_port, CK => clk
                           , RN => n5150, Q => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, QN => 
                           n_1110);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_22_port, CK => clk
                           , RN => n5143, Q => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, QN => 
                           n_1111);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_21_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, QN => 
                           n_1112);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_20_port, CK => clk
                           , RN => n5151, Q => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, QN => 
                           n_1113);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_19_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, QN => 
                           n_1114);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_18_port, CK => clk
                           , RN => n5146, Q => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, QN => 
                           n_1115);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_17_port, CK => clk
                           , RN => n5154, Q => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, QN => 
                           n_1116);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_16_port, CK => clk
                           , RN => n5147, Q => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, QN => 
                           n_1117);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_15_port, CK => clk
                           , RN => n5151, Q => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, QN => 
                           n_1118);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_14_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, QN => 
                           n_1119);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_13_port, CK => clk
                           , RN => n5155, Q => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, QN => 
                           n_1120);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_12_port, CK => clk
                           , RN => n5146, Q => n_1121, QN => n5133);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_5_11_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_out_6_11_port, QN => n_1122
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => n3094, CK => clk, RN => n5150, Q => 
                           boothmul_pipelined_i_sum_out_6_10_port, QN => n_1123
                           );
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_9_port, CK => clk, RN
                           => n5149, Q => boothmul_pipelined_i_sum_out_6_9_port
                           , QN => n_1124);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_8_port, CK => clk, RN
                           => n5150, Q => boothmul_pipelined_i_sum_out_6_8_port
                           , QN => n_1125);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_7_port, CK => clk, RN
                           => n5143, Q => boothmul_pipelined_i_sum_out_6_7_port
                           , QN => n_1126);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_6_port, CK => clk, RN
                           => n5154, Q => boothmul_pipelined_i_sum_out_6_6_port
                           , QN => n_1127);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_5_port, CK => clk, RN
                           => n5145, Q => boothmul_pipelined_i_sum_out_6_5_port
                           , QN => n_1128);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_4_port, CK => clk, RN
                           => n5148, Q => boothmul_pipelined_i_sum_out_6_4_port
                           , QN => n_1129);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_3_port, CK => clk, RN
                           => n5149, Q => boothmul_pipelined_i_sum_out_6_3_port
                           , QN => n_1130);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_2_port, CK => clk, RN
                           => n5145, Q => boothmul_pipelined_i_sum_out_6_2_port
                           , QN => n_1131);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_1_port, CK => clk, RN
                           => n5154, Q => boothmul_pipelined_i_sum_out_6_1_port
                           , QN => n_1132);
   boothmul_pipelined_i_pip_del_reg_addi_5_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_5_0_port, CK => clk, RN
                           => n5142, Q => boothmul_pipelined_i_sum_out_6_0_port
                           , QN => n_1133);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_54_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_6_58_port, QN => n5129
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_55_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_6_59_port, QN => 
                           n_1134);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_56_port, CK => 
                           clk, RN => n5152, Q => 
                           boothmul_pipelined_i_muxes_in_6_60_port, QN => 
                           n_1135);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_57_port, CK => 
                           clk, RN => n5143, Q => 
                           boothmul_pipelined_i_muxes_in_6_61_port, QN => 
                           n_1136);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_58_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_6_62_port, QN => 
                           n_1137);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_59_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_6_63_port, QN => 
                           n_1138);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_60_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_6_64_port, QN => 
                           n_1139);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_61_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_6_65_port, QN => 
                           n_1140);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_62_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_6_66_port, QN => 
                           n_1141);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_63_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_6_67_port, QN => 
                           n_1142);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_64_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_6_68_port, QN => 
                           n_1143);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_183_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_65_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_6_69_port, QN => 
                           n_1144);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_182_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_66_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_6_70_port, QN => 
                           n_1145);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_181_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_67_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_6_71_port, QN => 
                           n_1146);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_180_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_68_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_6_72_port, QN => 
                           n_1147);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_179_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_205_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_6_73_port, QN => n5123
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_189_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_6_203_port, QN => 
                           n_1148);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_190_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_6_204_port, QN => 
                           n_1149);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_191_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_6_205_port, QN => 
                           n_1150);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_56_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_192_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_6_206_port, QN => 
                           n_1151);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_55_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_193_port, CK => 
                           clk, RN => n5142, Q => 
                           boothmul_pipelined_i_muxes_in_6_207_port, QN => 
                           n_1152);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_54_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_194_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_6_208_port, QN => 
                           n_1153);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_53_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_195_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_6_209_port, QN => 
                           n_1154);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_52_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_196_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_6_210_port, QN => 
                           n_1155);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_51_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_197_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_6_211_port, QN => 
                           n_1156);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_50_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_198_port, CK => 
                           clk, RN => n5142, Q => 
                           boothmul_pipelined_i_muxes_in_6_212_port, QN => 
                           n_1157);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_49_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_199_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_6_213_port, QN => 
                           n_1158);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_48_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_200_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_6_214_port, QN => 
                           n_1159);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_47_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_201_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_6_215_port, QN => 
                           n_1160);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_46_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_202_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_6_216_port, QN => 
                           n_1161);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_45_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_203_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_6_217_port, QN => 
                           n_1162);
   boothmul_pipelined_i_pip_del_reg_muxi_5_D_I_44_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_5_204_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_6_218_port, QN => 
                           n_1163);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_24_port, CK => clk
                           , RN => n5143, Q => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, QN => 
                           n_1164);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_23_port, CK => clk
                           , RN => n5150, Q => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, QN => 
                           n_1165);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_22_port, CK => clk
                           , RN => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, QN => 
                           n_1166);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_21_port, CK => clk
                           , RN => n5145, Q => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, QN => 
                           n_1167);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_20_port, CK => clk
                           , RN => n5144, Q => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, QN => 
                           n_1168);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_19_port, CK => clk
                           , RN => n5145, Q => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, QN => 
                           n_1169);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_18_port, CK => clk
                           , RN => n5145, Q => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, QN => 
                           n_1170);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_17_port, CK => clk
                           , RN => n5146, Q => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, QN => 
                           n_1171);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_16_port, CK => clk
                           , RN => n5143, Q => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, QN => 
                           n_1172);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_15_port, CK => clk
                           , RN => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, QN => 
                           n_1173);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_14_port, CK => clk
                           , RN => n5148, Q => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, QN => 
                           n_1174);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_13_port, CK => clk
                           , RN => n5154, Q => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, QN => 
                           n_1175);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_12_port, CK => clk
                           , RN => n5148, Q => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, QN => 
                           n_1176);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_11_port, CK => clk
                           , RN => n5142, Q => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, QN => 
                           n_1177);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_4_10_port, CK => clk
                           , RN => n5146, Q => n_1178, QN => n5132);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_9_port, CK => clk, RN
                           => n5152, Q => boothmul_pipelined_i_sum_out_5_9_port
                           , QN => n_1179);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           n3093, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_5_8_port, QN => n_1180)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_7_port, CK => clk, RN
                           => n5144, Q => boothmul_pipelined_i_sum_out_5_7_port
                           , QN => n_1181);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_6_port, CK => clk, RN
                           => n5152, Q => boothmul_pipelined_i_sum_out_5_6_port
                           , QN => n_1182);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_5_port, CK => clk, RN
                           => n5154, Q => boothmul_pipelined_i_sum_out_5_5_port
                           , QN => n_1183);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_4_port, CK => clk, RN
                           => n5152, Q => boothmul_pipelined_i_sum_out_5_4_port
                           , QN => n_1184);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_3_port, CK => clk, RN
                           => n5154, Q => boothmul_pipelined_i_sum_out_5_3_port
                           , QN => n_1185);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_2_port, CK => clk, RN
                           => n5154, Q => boothmul_pipelined_i_sum_out_5_2_port
                           , QN => n_1186);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_1_port, CK => clk, RN
                           => n5152, Q => boothmul_pipelined_i_sum_out_5_1_port
                           , QN => n_1187);
   boothmul_pipelined_i_pip_del_reg_addi_4_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_4_0_port, CK => clk, RN
                           => n5146, Q => boothmul_pipelined_i_sum_out_5_0_port
                           , QN => n_1188);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_50_port, CK => 
                           clk, RN => n5142, Q => 
                           boothmul_pipelined_i_muxes_in_5_54_port, QN => n5128
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_51_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_5_55_port, QN => 
                           n_1189);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_52_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_56_port, QN => 
                           n_1190);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_53_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_5_57_port, QN => 
                           n_1191);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_54_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_5_58_port, QN => 
                           n_1192);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_55_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_5_59_port, QN => 
                           n_1193);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_56_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_5_60_port, QN => 
                           n_1194);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_57_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_5_61_port, QN => 
                           n_1195);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_58_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_5_62_port, QN => 
                           n_1196);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_59_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_5_63_port, QN => 
                           n_1197);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_60_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_5_64_port, QN => 
                           n_1198);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_61_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_5_65_port, QN => 
                           n_1199);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_186_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_62_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_5_66_port, QN => 
                           n_1200);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_185_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_63_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_5_67_port, QN => 
                           n_1201);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_184_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_64_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_5_68_port, QN => 
                           n_1202);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_175_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_5_189_port, QN => 
                           n_1203);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_176_port, CK => 
                           clk, RN => n5142, Q => 
                           boothmul_pipelined_i_muxes_in_5_190_port, QN => 
                           n_1204);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_71_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_177_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_5_191_port, QN => 
                           n_1205);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_70_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_178_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_5_192_port, QN => 
                           n_1206);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_69_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_179_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_5_193_port, QN => 
                           n_1207);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_68_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_180_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_5_194_port, QN => 
                           n_1208);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_67_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_181_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_5_195_port, QN => 
                           n_1209);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_66_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_182_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_5_196_port, QN => 
                           n_1210);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_65_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_183_port, CK => 
                           clk, RN => n5152, Q => 
                           boothmul_pipelined_i_muxes_in_5_197_port, QN => 
                           n_1211);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_64_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_184_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_5_198_port, QN => 
                           n_1212);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_63_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_185_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_5_199_port, QN => 
                           n_1213);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_62_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_186_port, CK => 
                           clk, RN => n5143, Q => 
                           boothmul_pipelined_i_muxes_in_5_200_port, QN => 
                           n_1214);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_61_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_187_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_5_201_port, QN => 
                           n_1215);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_60_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_188_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_5_202_port, QN => 
                           n_1216);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_59_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_189_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_5_203_port, QN => 
                           n_1217);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_58_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_190_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_5_204_port, QN => 
                           n_1218);
   boothmul_pipelined_i_pip_del_reg_muxi_4_D_I_57_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_4_65_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_5_205_port, QN => 
                           n5122);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_22_port, CK => clk
                           , RN => n5146, Q => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, QN => 
                           n_1219);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_21_port, CK => clk
                           , RN => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, QN => 
                           n_1220);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_20_port, CK => clk
                           , RN => n5151, Q => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, QN => 
                           n_1221);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_19_port, CK => clk
                           , RN => n5151, Q => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, QN => 
                           n_1222);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_18_port, CK => clk
                           , RN => n5143, Q => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, QN => 
                           n_1223);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_17_port, CK => clk
                           , RN => n5148, Q => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, QN => 
                           n_1224);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_16_port, CK => clk
                           , RN => n5155, Q => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, QN => 
                           n_1225);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_15_port, CK => clk
                           , RN => n5152, Q => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, QN => 
                           n_1226);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_14_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, QN => 
                           n_1227);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_13_port, CK => clk
                           , RN => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, QN => 
                           n_1228);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_12_port, CK => clk
                           , RN => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, QN => 
                           n_1229);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_11_port, CK => clk
                           , RN => n5144, Q => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, QN => 
                           n_1230);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_3_10_port, CK => clk
                           , RN => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, QN => 
                           n_1231);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_9_port, CK => clk, RN
                           => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, QN => n_1232
                           );
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_8_port, CK => clk, RN
                           => n5147, Q => n_1233, QN => n5131);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_7_port, CK => clk, RN
                           => n5149, Q => boothmul_pipelined_i_sum_out_4_7_port
                           , QN => n_1234);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           n3092, CK => clk, RN => n5149, Q => 
                           boothmul_pipelined_i_sum_out_4_6_port, QN => n_1235)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_5_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_out_4_5_port, QN => n_1236)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_4_port, CK => clk, RN
                           => n5146, Q => boothmul_pipelined_i_sum_out_4_4_port
                           , QN => n_1237);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_3_port, CK => clk, RN
                           => n5152, Q => boothmul_pipelined_i_sum_out_4_3_port
                           , QN => n_1238);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_2_port, CK => clk, RN
                           => n5147, Q => boothmul_pipelined_i_sum_out_4_2_port
                           , QN => n_1239);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_1_port, CK => clk, RN
                           => n5143, Q => boothmul_pipelined_i_sum_out_4_1_port
                           , QN => n_1240);
   boothmul_pipelined_i_pip_del_reg_addi_3_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_3_0_port, CK => clk, RN
                           => n5141, Q => boothmul_pipelined_i_sum_out_4_0_port
                           , QN => n_1241);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_46_port, CK => 
                           clk, RN => n5152, Q => 
                           boothmul_pipelined_i_muxes_in_4_50_port, QN => n5127
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_47_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_4_51_port, QN => 
                           n_1242);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_48_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_4_52_port, QN => 
                           n_1243);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_49_port, CK => 
                           clk, RN => n5143, Q => 
                           boothmul_pipelined_i_muxes_in_4_53_port, QN => 
                           n_1244);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_50_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_4_54_port, QN => 
                           n_1245);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_51_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_4_55_port, QN => 
                           n_1246);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_52_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_4_56_port, QN => 
                           n_1247);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_53_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_4_57_port, QN => 
                           n_1248);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_54_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_4_58_port, QN => 
                           n_1249);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_55_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_4_59_port, QN => 
                           n_1250);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_56_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_4_60_port, QN => 
                           n_1251);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_191_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_57_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_4_61_port, QN => 
                           n_1252);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_190_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_58_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_4_62_port, QN => 
                           n_1253);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_189_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_59_port, CK => 
                           clk, RN => n5142, Q => 
                           boothmul_pipelined_i_muxes_in_4_63_port, QN => 
                           n_1254);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_188_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_60_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_4_64_port, QN => 
                           n_1255);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_187_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_177_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_4_65_port, QN => n5121
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_161_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_4_175_port, QN => 
                           n_1256);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_162_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_4_176_port, QN => 
                           n_1257);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_163_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_4_177_port, QN => 
                           n_1258);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_84_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_164_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_4_178_port, QN => 
                           n_1259);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_83_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_165_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_4_179_port, QN => 
                           n_1260);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_82_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_166_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_4_180_port, QN => 
                           n_1261);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_81_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_167_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_4_181_port, QN => 
                           n_1262);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_80_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_168_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_4_182_port, QN => 
                           n_1263);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_79_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_169_port, CK => 
                           clk, RN => n5143, Q => 
                           boothmul_pipelined_i_muxes_in_4_183_port, QN => 
                           n_1264);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_78_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_170_port, CK => 
                           clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_4_184_port, QN => 
                           n_1265);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_77_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_171_port, CK => 
                           clk, RN => n5143, Q => 
                           boothmul_pipelined_i_muxes_in_4_185_port, QN => 
                           n_1266);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_76_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_172_port, CK => 
                           clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_4_186_port, QN => 
                           n_1267);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_75_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_173_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_4_187_port, QN => 
                           n_1268);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_74_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_174_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_4_188_port, QN => 
                           n_1269);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_73_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_175_port, CK => 
                           clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_4_189_port, QN => 
                           n_1270);
   boothmul_pipelined_i_pip_del_reg_muxi_3_D_I_72_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_3_176_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_4_190_port, QN => 
                           n_1271);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_20_port, CK => clk
                           , RN => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, QN => 
                           n_1272);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_19_port, CK => clk
                           , RN => n5152, Q => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, QN => 
                           n_1273);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_18_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, QN => 
                           n_1274);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_17_port, CK => clk
                           , RN => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, QN => 
                           n_1275);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_16_port, CK => clk
                           , RN => n5150, Q => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, QN => 
                           n_1276);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_15_port, CK => clk
                           , RN => n5147, Q => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, QN => 
                           n_1277);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_14_port, CK => clk
                           , RN => n5144, Q => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, QN => 
                           n_1278);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_13_port, CK => clk
                           , RN => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, QN => 
                           n_1279);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_12_port, CK => clk
                           , RN => n5152, Q => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, QN => 
                           n_1280);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_11_port, CK => clk
                           , RN => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, QN => 
                           n_1281);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_2_10_port, CK => clk
                           , RN => n5143, Q => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, QN => 
                           n_1282);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_9_port, CK => clk, RN
                           => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, QN => n_1283
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_8_port, CK => clk, RN
                           => n5148, Q => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, QN => n_1284
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_7_port, CK => clk, RN
                           => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, QN => n_1285
                           );
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_6_port, CK => clk, RN
                           => n5149, Q => n_1286, QN => n5124);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_5_port, CK => clk, RN
                           => n5148, Q => boothmul_pipelined_i_sum_out_3_5_port
                           , QN => n_1287);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           n3091, CK => clk, RN => n5147, Q => 
                           boothmul_pipelined_i_sum_out_3_4_port, QN => n_1288)
                           ;
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_3_port, CK => clk, RN
                           => n5146, Q => boothmul_pipelined_i_sum_out_3_3_port
                           , QN => n_1289);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_2_port, CK => clk, RN
                           => n5152, Q => boothmul_pipelined_i_sum_out_3_2_port
                           , QN => n_1290);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_1_port, CK => clk, RN
                           => n5148, Q => boothmul_pipelined_i_sum_out_3_1_port
                           , QN => n_1291);
   boothmul_pipelined_i_pip_del_reg_addi_2_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_2_0_port, CK => clk, RN
                           => n5142, Q => boothmul_pipelined_i_sum_out_3_0_port
                           , QN => n_1292);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_206_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_15_port, CK => clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_3_46_port, QN => n7164
                           );
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_205_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_14_port, CK => clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_3_47_port, QN => 
                           n_1293);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_204_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_13_port, CK => clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_3_48_port, QN => 
                           n_1294);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_203_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_12_port, CK => clk, RN => n5152, Q => 
                           boothmul_pipelined_i_muxes_in_3_49_port, QN => 
                           n_1295);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_202_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_11_port, CK => clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_3_50_port, QN => 
                           n_1296);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_201_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_10_port, CK => clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_3_51_port, QN => 
                           n_1297);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_200_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_9_port, CK => clk, RN => n5151, Q => 
                           boothmul_pipelined_i_muxes_in_3_52_port, QN => 
                           n_1298);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_199_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_8_port, CK => clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_3_53_port, QN => 
                           n_1299);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_198_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_7_port, CK => clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_3_54_port, QN => 
                           n_1300);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_197_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_6_port, CK => clk, RN => n5144, Q => 
                           boothmul_pipelined_i_muxes_in_3_55_port, QN => 
                           n_1301);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_196_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_5_port, CK => clk, RN => n5146, Q => 
                           boothmul_pipelined_i_muxes_in_3_56_port, QN => 
                           n_1302);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_195_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_4_port, CK => clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_3_57_port, QN => 
                           n_1303);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_194_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_3_port, CK => clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_58_port, QN => 
                           n_1304);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_193_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_2_port, CK => clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_3_59_port, QN => 
                           n_1305);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_192_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_1_port, CK => clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_3_60_port, QN => 
                           n_1306);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_101_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_119_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_3_161_port, QN => 
                           n_1307);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_100_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_102_port, CK => 
                           clk, RN => n5152, Q => 
                           boothmul_pipelined_i_muxes_in_3_162_port, QN => 
                           n_1308);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_99_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_103_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_3_163_port, QN => 
                           n_1309);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_98_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_104_port, CK => 
                           clk, RN => n5143, Q => 
                           boothmul_pipelined_i_muxes_in_3_164_port, QN => 
                           n_1310);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_97_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_105_port, CK => 
                           clk, RN => n5149, Q => 
                           boothmul_pipelined_i_muxes_in_3_165_port, QN => 
                           n_1311);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_96_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_106_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_3_166_port, QN => 
                           n_1312);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_95_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_107_port, CK => 
                           clk, RN => n5147, Q => 
                           boothmul_pipelined_i_muxes_in_3_167_port, QN => 
                           n_1313);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_94_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_108_port, CK => 
                           clk, RN => n5148, Q => 
                           boothmul_pipelined_i_muxes_in_3_168_port, QN => 
                           n_1314);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_93_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_109_port, CK => 
                           clk, RN => n5154, Q => 
                           boothmul_pipelined_i_muxes_in_3_169_port, QN => 
                           n_1315);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_92_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_110_port, CK => 
                           clk, RN => n5155, Q => 
                           boothmul_pipelined_i_muxes_in_3_170_port, QN => 
                           n_1316);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_91_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_111_port, CK => 
                           clk, RN => n5150, Q => 
                           boothmul_pipelined_i_muxes_in_3_171_port, QN => 
                           n_1317);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_90_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_112_port, CK => 
                           clk, RN => n5145, Q => 
                           boothmul_pipelined_i_muxes_in_3_172_port, QN => 
                           n_1318);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_89_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_113_port, CK => 
                           clk, RN => rst_BAR, Q => 
                           boothmul_pipelined_i_muxes_in_3_173_port, QN => 
                           n_1319);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_88_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_114_port, CK => 
                           clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_3_174_port, QN => 
                           n_1320);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_87_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_115_port, CK => 
                           clk, RN => n5142, Q => 
                           boothmul_pipelined_i_muxes_in_3_175_port, QN => 
                           n_1321);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_86_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_muxes_in_0_116_port, CK => 
                           clk, RN => n5153, Q => 
                           boothmul_pipelined_i_muxes_in_3_176_port, QN => 
                           n_1322);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_18_port, CK => clk
                           , RN => n5148, Q => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, QN => 
                           n_1323);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_17_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, QN => 
                           n_1324);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_16_port, CK => clk
                           , RN => n5149, Q => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, QN => 
                           n_1325);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_15_port, CK => clk
                           , RN => n5154, Q => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, QN => 
                           n_1326);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_14_port, CK => clk
                           , RN => n5155, Q => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, QN => 
                           n_1327);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_13_port, CK => clk
                           , RN => n5151, Q => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, QN => 
                           n_1328);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_12_port, CK => clk
                           , RN => n5145, Q => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, QN => 
                           n_1329);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_11_port, CK => clk
                           , RN => n5150, Q => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, QN => 
                           n_1330);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => boothmul_pipelined_i_sum_out_1_10_port, CK => clk
                           , RN => n5150, Q => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, QN => 
                           n_1331);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_9_port, CK => clk, RN
                           => n5141, Q => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, QN => n_1332
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_8_port, CK => clk, RN
                           => rst_BAR, Q => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, QN => n_1333
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_7_port, CK => clk, RN
                           => n5153, Q => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, QN => n_1334
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_6_port, CK => clk, RN
                           => n5147, Q => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, QN => n_1335
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_5_port, CK => clk, RN
                           => n5142, Q => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, QN => n_1336
                           );
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_4_port, CK => clk, RN
                           => n5142, Q => n_1337, QN => n5130);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_3_port, CK => clk, RN
                           => n5143, Q => boothmul_pipelined_i_sum_out_2_3_port
                           , QN => n_1338);
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           n3086, CK => clk, RN => n5142, Q => 
                           boothmul_pipelined_i_sum_out_2_2_port, QN => n_1339)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           n1988, CK => clk, RN => n5151, Q => 
                           boothmul_pipelined_i_sum_out_2_1_port, QN => n_1340)
                           ;
   boothmul_pipelined_i_pip_del_reg_add1_1_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           boothmul_pipelined_i_sum_out_1_0_port, CK => clk, RN
                           => n5143, Q => boothmul_pipelined_i_sum_out_2_0_port
                           , QN => n_1341);
   boothmul_pipelined_i_pip_del_reg_muxi_2_D_I_85_Q_reg : DFFR_X1 port map( D 
                           => data1_mul_0_port, CK => clk, RN => n5141, Q => 
                           boothmul_pipelined_i_muxes_in_3_177_port, QN => 
                           n3077);
   DATA2_I_reg_31_inst : DLL_X1 port map( D => N2548, GN => n1992, Q => 
                           DATA2_I_31_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_1 : HA_X1 port map( 
                           A => n1989, B => n1990, CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, S 
                           => boothmul_pipelined_i_muxes_in_0_116_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_2 : HA_X1 port map( 
                           A => n1987, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_2_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, S 
                           => boothmul_pipelined_i_muxes_in_0_115_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_3 : HA_X1 port map( 
                           A => n1986, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_3_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, S 
                           => boothmul_pipelined_i_muxes_in_0_114_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_4 : HA_X1 port map( 
                           A => n1984, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, S 
                           => boothmul_pipelined_i_muxes_in_0_113_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_5 : HA_X1 port map( 
                           A => n1982, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, S 
                           => boothmul_pipelined_i_muxes_in_0_112_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_6 : HA_X1 port map( 
                           A => n1980, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, S 
                           => boothmul_pipelined_i_muxes_in_0_111_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_7 : HA_X1 port map( 
                           A => n1978, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, S 
                           => boothmul_pipelined_i_muxes_in_0_110_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_8 : HA_X1 port map( 
                           A => n1976, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, S 
                           => boothmul_pipelined_i_muxes_in_0_109_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_9 : HA_X1 port map( 
                           A => n1974, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, S 
                           => boothmul_pipelined_i_muxes_in_0_108_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_10 : HA_X1 port map(
                           A => n1972, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, S 
                           => boothmul_pipelined_i_muxes_in_0_107_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_11 : HA_X1 port map(
                           A => n1970, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, S 
                           => boothmul_pipelined_i_muxes_in_0_106_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_12 : HA_X1 port map(
                           A => n1968, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, S 
                           => boothmul_pipelined_i_muxes_in_0_105_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_13 : HA_X1 port map(
                           A => n1966, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, S 
                           => boothmul_pipelined_i_muxes_in_0_104_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_14 : HA_X1 port map(
                           A => n1964, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, S 
                           => boothmul_pipelined_i_muxes_in_0_103_port);
   boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_U1_1_15 : HA_X1 port map(
                           A => n1962, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, S 
                           => boothmul_pipelined_i_muxes_in_0_102_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_3 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_3_port, B => n1985, 
                           CI => n3083, CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, S 
                           => boothmul_pipelined_i_sum_out_1_3_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_4 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_4_port, B => n1983, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_4_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, S 
                           => boothmul_pipelined_i_sum_out_1_4_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_5_port, B => n1981, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_5_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_1_5_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_6_port, B => n1979, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_1_6_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_7_port, B => n1977, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_1_7_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_8_port, B => n1975, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_1_8_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_1_9_port, B => n1973, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_1_9_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_10_port, B => n1971, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_1_10_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_11_port, B => n1969, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_1_11_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_12_port, B => n1967, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_1_12_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_13_port, B => n1965, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_1_13_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_14_port, B => n1963, 
                           CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_1_14_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_15_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_1_15_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_1_16_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_1_17_port);
   boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_1_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_1_18_port, CI => 
                           boothmul_pipelined_i_ADD1_1_add_1_root_add_21_2_carry_18_port, 
                           CO => n_1342, S => 
                           boothmul_pipelined_i_sum_out_1_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_5 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_5_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_5_port, CI => n3085,
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, S 
                           => boothmul_pipelined_i_sum_out_2_5_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_6 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_6_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_6_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_6_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, S 
                           => boothmul_pipelined_i_sum_out_2_6_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_7_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_7_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_2_7_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_8_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_2_8_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_2_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_9_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_2_9_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_10_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_2_10_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_11_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_2_11_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_12_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_2_12_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_13_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_2_13_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_14_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_2_14_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_15_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_2_15_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_16_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_2_16_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_17_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_2_17_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_2_18_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_2_19_port);
   boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_2_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_2_20_port, CI => 
                           boothmul_pipelined_i_ADDi_2_add_1_root_add_21_2_carry_20_port, 
                           CO => n_1343, S => 
                           boothmul_pipelined_i_sum_out_2_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_7 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_7_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_7_port, CI => n3084,
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, S 
                           => boothmul_pipelined_i_sum_out_3_7_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_8 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_8_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_8_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_8_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, S 
                           => boothmul_pipelined_i_sum_out_3_8_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_3_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_9_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_9_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_3_9_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_10_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_3_10_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_11_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_3_11_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_12_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_3_12_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_13_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_3_13_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_14_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_3_14_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_15_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_3_15_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_16_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_3_16_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_17_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_3_17_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_18_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_3_18_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_19_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_3_19_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_3_20_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_3_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_3_22_port, CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_3_21_port);
   boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           n1991, B => boothmul_pipelined_i_sum_B_in_3_22_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_3_add_1_root_add_21_2_carry_22_port, 
                           CO => n_1344, S => 
                           boothmul_pipelined_i_sum_out_3_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_9 : FA_X1 port map( A => 
                           boothmul_pipelined_i_mux_out_4_9_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_9_port, CI => n3090,
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, S 
                           => boothmul_pipelined_i_sum_out_4_9_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_10 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_10_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_10_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_10_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, S 
                           => boothmul_pipelined_i_sum_out_4_10_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_11_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_11_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_4_11_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_12_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_4_12_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_13_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_4_13_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_14_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_4_14_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_15_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_4_15_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_16_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_4_16_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_17_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_4_17_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_18_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_4_18_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_19_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_4_19_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_20_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_4_20_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_21_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_4_21_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_4_22_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_4_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_4_24_port, CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_4_23_port);
   boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           n1997, B => boothmul_pipelined_i_sum_B_in_4_24_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_4_add_1_root_add_21_2_carry_24_port, 
                           CO => n_1345, S => 
                           boothmul_pipelined_i_sum_out_4_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_11 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_11_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_11_port, CI => n3089
                           , CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, S 
                           => boothmul_pipelined_i_sum_out_5_11_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_12 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_12_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_12_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_12_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, S 
                           => boothmul_pipelined_i_sum_out_5_12_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_13_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_13_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_5_13_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_14_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_5_14_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_15_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_5_15_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_16_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_5_16_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_17_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_5_17_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_18_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_5_18_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_19_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_5_19_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_20_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_5_20_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_21_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_5_21_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_22_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_5_22_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_23_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_5_23_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_5_24_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_5_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_5_26_port, CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_5_25_port);
   boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           n1996, B => boothmul_pipelined_i_sum_B_in_5_26_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_5_add_1_root_add_21_2_carry_26_port, 
                           CO => n_1346, S => 
                           boothmul_pipelined_i_sum_out_5_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_13 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_13_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_13_port, CI => n3088
                           , CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, S 
                           => boothmul_pipelined_i_sum_out_6_13_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_14 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_14_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_14_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_14_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, S 
                           => boothmul_pipelined_i_sum_out_6_14_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_15_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_15_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, S 
                           => boothmul_pipelined_i_sum_out_6_15_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_16_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, S 
                           => boothmul_pipelined_i_sum_out_6_16_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_17_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, S 
                           => boothmul_pipelined_i_sum_out_6_17_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_18_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, S 
                           => boothmul_pipelined_i_sum_out_6_18_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_19_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, S 
                           => boothmul_pipelined_i_sum_out_6_19_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_20_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, S 
                           => boothmul_pipelined_i_sum_out_6_20_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_21_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, S 
                           => boothmul_pipelined_i_sum_out_6_21_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_22_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, S 
                           => boothmul_pipelined_i_sum_out_6_22_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_23_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, S 
                           => boothmul_pipelined_i_sum_out_6_23_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_24_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, S 
                           => boothmul_pipelined_i_sum_out_6_24_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_25_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, S 
                           => boothmul_pipelined_i_sum_out_6_25_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, S 
                           => boothmul_pipelined_i_sum_out_6_26_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_6_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_6_28_port, CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, S 
                           => boothmul_pipelined_i_sum_out_6_27_port);
   boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           n1995, B => boothmul_pipelined_i_sum_B_in_6_28_port,
                           CI => 
                           boothmul_pipelined_i_ADDi_6_add_1_root_add_21_2_carry_28_port, 
                           CO => n_1347, S => 
                           boothmul_pipelined_i_sum_out_6_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_15 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_15_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_15_port, CI => n3087
                           , CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, S 
                           => dataout_mul_15_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_16 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_16_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_16_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_16_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, S 
                           => dataout_mul_16_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_17 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_17_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_17_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_17_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, S 
                           => dataout_mul_17_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_18 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_18_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_18_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_18_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, S 
                           => dataout_mul_18_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_19 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_19_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_19_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_19_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, S 
                           => dataout_mul_19_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_20 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_20_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_20_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_20_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, S 
                           => dataout_mul_20_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_21 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_21_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_21_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_21_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, S 
                           => dataout_mul_21_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_22 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_22_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_22_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_22_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, S 
                           => dataout_mul_22_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_23 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_23_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_23_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_23_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, S 
                           => dataout_mul_23_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_24 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_24_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_24_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_24_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, S 
                           => dataout_mul_24_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_25 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_25_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_25_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_25_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, S 
                           => dataout_mul_25_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_26 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_26_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_26_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_26_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, S 
                           => dataout_mul_26_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_27 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_27_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_27_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_27_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, S 
                           => dataout_mul_27_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_28 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_28_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_28_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, S 
                           => dataout_mul_28_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_29 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_29_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_29_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, S 
                           => dataout_mul_29_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_30 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_30_port, 
                           CO => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, S 
                           => dataout_mul_30_port);
   boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_U1_31 : FA_X1 port map( A =>
                           boothmul_pipelined_i_mux_out_7_30_port, B => 
                           boothmul_pipelined_i_sum_B_in_7_30_port, CI => 
                           boothmul_pipelined_i_ADDn_7_add_1_root_add_21_2_carry_31_port, 
                           CO => n_1348, S => dataout_mul_31_port);
   data2_mul_reg_1_inst : DLL_X1 port map( D => DATA2(1), GN => n553, Q => 
                           data2_mul_1_port);
   DATA2_I_reg_30_inst : DLL_X1 port map( D => N2547, GN => n1992, Q => 
                           DATA2_I_30_port);
   DATA2_I_reg_29_inst : DLL_X1 port map( D => N2546, GN => n1992, Q => 
                           DATA2_I_29_port);
   U3 : CLKBUF_X1 port map( A => n5144, Z => n5141);
   U4 : CLKBUF_X1 port map( A => n5144, Z => n5142);
   U5 : CLKBUF_X1 port map( A => n5144, Z => n5143);
   U6 : CLKBUF_X1 port map( A => rst_BAR, Z => n5144);
   U7 : CLKBUF_X1 port map( A => n5148, Z => n5145);
   U8 : CLKBUF_X1 port map( A => n5141, Z => n5146);
   U9 : CLKBUF_X1 port map( A => n5142, Z => n5147);
   U10 : CLKBUF_X1 port map( A => n5142, Z => n5148);
   U11 : CLKBUF_X1 port map( A => n5142, Z => n5149);
   U12 : CLKBUF_X1 port map( A => n5142, Z => n5150);
   U13 : CLKBUF_X1 port map( A => n5143, Z => n5151);
   U14 : CLKBUF_X1 port map( A => n5143, Z => n5152);
   U15 : CLKBUF_X1 port map( A => n5143, Z => n5153);
   U16 : CLKBUF_X1 port map( A => n5143, Z => n5154);
   U17 : CLKBUF_X1 port map( A => n5143, Z => n5155);
   U18 : NOR2_X2 port map( A1 => n5412, A2 => n5228, ZN => n6232);
   U19 : CLKBUF_X1 port map( A => n6868, Z => n6858);
   U20 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n5156);
   U21 : INV_X1 port map( A => FUNC(2), ZN => n6773);
   U22 : NAND2_X1 port map( A1 => n5156, A2 => n6773, ZN => n1992);
   U23 : CLKBUF_X1 port map( A => n1992, Z => n7166);
   U24 : CLKBUF_X1 port map( A => DATA1(14), Z => n7169);
   U25 : INV_X1 port map( A => data2_mul_1_port, ZN => n5157);
   U26 : NOR2_X1 port map( A1 => boothmul_pipelined_i_encoder_out_0_0_port, A2 
                           => n5157, ZN => n5166);
   U27 : CLKBUF_X1 port map( A => n5166, Z => n7139);
   U28 : NAND2_X1 port map( A1 => n5157, A2 => 
                           boothmul_pipelined_i_encoder_out_0_0_port, ZN => 
                           n7142);
   U29 : INV_X1 port map( A => n7142, ZN => n5174);
   U30 : INV_X1 port map( A => boothmul_pipelined_i_encoder_out_0_0_port, ZN =>
                           n6870);
   U31 : NOR2_X1 port map( A1 => n5157, A2 => n6870, ZN => n7140);
   U32 : CLKBUF_X1 port map( A => n7140, Z => n5171);
   U33 : AOI222_X1 port map( A1 => data1_mul_0_port, A2 => n7139, B1 => 
                           data1_mul_1_port, B2 => n5174, C1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, C2 => 
                           n5171, ZN => n5158);
   U34 : INV_X1 port map( A => n5158, ZN => n1988);
   U35 : AOI222_X1 port map( A1 => n7139, A2 => 
                           boothmul_pipelined_i_muxes_in_0_115_port, B1 => 
                           data1_mul_3_port, B2 => n5174, C1 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, C2 => 
                           n7140, ZN => n5159);
   U36 : INV_X1 port map( A => n5159, ZN => n1985);
   U37 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, A2
                           => n5166, B1 => data1_mul_4_port, B2 => n5174, C1 =>
                           boothmul_pipelined_i_muxes_in_0_113_port, C2 => 
                           n7140, ZN => n5160);
   U38 : INV_X1 port map( A => n5160, ZN => n1983);
   U39 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, A2
                           => n5166, B1 => data1_mul_5_port, B2 => n5174, C1 =>
                           boothmul_pipelined_i_muxes_in_0_112_port, C2 => 
                           n5171, ZN => n5161);
   U40 : INV_X1 port map( A => n5161, ZN => n1981);
   U41 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, A2
                           => n5166, B1 => data1_mul_6_port, B2 => n5174, C1 =>
                           boothmul_pipelined_i_muxes_in_0_111_port, C2 => 
                           n5171, ZN => n5162);
   U42 : INV_X1 port map( A => n5162, ZN => n1979);
   U43 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, A2
                           => n5166, B1 => data1_mul_7_port, B2 => n5174, C1 =>
                           boothmul_pipelined_i_muxes_in_0_110_port, C2 => 
                           n7140, ZN => n5163);
   U44 : INV_X1 port map( A => n5163, ZN => n1977);
   U45 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, A2
                           => n5166, B1 => data1_mul_8_port, B2 => n5174, C1 =>
                           boothmul_pipelined_i_muxes_in_0_109_port, C2 => 
                           n5171, ZN => n5164);
   U46 : INV_X1 port map( A => n5164, ZN => n1975);
   U47 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, A2
                           => n5166, B1 => data1_mul_9_port, B2 => n5174, C1 =>
                           boothmul_pipelined_i_muxes_in_0_108_port, C2 => 
                           n5171, ZN => n5165);
   U48 : INV_X1 port map( A => n5165, ZN => n1973);
   U49 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, A2
                           => n5166, B1 => data1_mul_10_port, B2 => n5174, C1 
                           => boothmul_pipelined_i_muxes_in_0_107_port, C2 => 
                           n5171, ZN => n5167);
   U50 : INV_X1 port map( A => n5167, ZN => n1971);
   U51 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, A2
                           => n7139, B1 => data1_mul_11_port, B2 => n5174, C1 
                           => boothmul_pipelined_i_muxes_in_0_106_port, C2 => 
                           n7140, ZN => n5168);
   U52 : INV_X1 port map( A => n5168, ZN => n1969);
   U53 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, A2
                           => n7139, B1 => data1_mul_12_port, B2 => n5174, C1 
                           => boothmul_pipelined_i_muxes_in_0_105_port, C2 => 
                           n5171, ZN => n5169);
   U54 : INV_X1 port map( A => n5169, ZN => n1967);
   U55 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, A2
                           => n7139, B1 => data1_mul_13_port, B2 => n5174, C1 
                           => boothmul_pipelined_i_muxes_in_0_104_port, C2 => 
                           n7140, ZN => n5170);
   U56 : INV_X1 port map( A => n5170, ZN => n1965);
   U57 : AOI222_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, A2
                           => n7139, B1 => data1_mul_14_port, B2 => n5174, C1 
                           => boothmul_pipelined_i_muxes_in_0_103_port, C2 => 
                           n5171, ZN => n5172);
   U58 : INV_X1 port map( A => n5172, ZN => n1963);
   U59 : INV_X1 port map( A => data1_mul_0_port, ZN => n1990);
   U60 : CLKBUF_X1 port map( A => DATA1(12), Z => n7168);
   U61 : CLKBUF_X1 port map( A => DATA1(10), Z => n7167);
   U62 : NOR3_X1 port map( A1 => FUNC(0), A2 => FUNC(1), A3 => n6773, ZN => 
                           n5343);
   U63 : INV_X1 port map( A => FUNC(3), ZN => n6832);
   U64 : NAND2_X1 port map( A1 => n5343, A2 => n6832, ZN => n553);
   U65 : INV_X1 port map( A => data1_mul_1_port, ZN => n1989);
   U66 : INV_X1 port map( A => data1_mul_2_port, ZN => n1987);
   U67 : INV_X1 port map( A => data1_mul_3_port, ZN => n1986);
   U68 : INV_X1 port map( A => data1_mul_4_port, ZN => n1984);
   U69 : INV_X1 port map( A => data1_mul_5_port, ZN => n1982);
   U70 : INV_X1 port map( A => data1_mul_6_port, ZN => n1980);
   U71 : INV_X1 port map( A => data1_mul_7_port, ZN => n1978);
   U72 : INV_X1 port map( A => data1_mul_8_port, ZN => n1976);
   U73 : INV_X1 port map( A => data1_mul_9_port, ZN => n1974);
   U74 : INV_X1 port map( A => data1_mul_10_port, ZN => n1972);
   U75 : INV_X1 port map( A => data1_mul_11_port, ZN => n1970);
   U76 : INV_X1 port map( A => data1_mul_12_port, ZN => n1968);
   U77 : INV_X1 port map( A => data1_mul_13_port, ZN => n1966);
   U78 : INV_X1 port map( A => data1_mul_14_port, ZN => n1964);
   U79 : INV_X1 port map( A => data1_mul_15_port, ZN => n1962);
   U80 : XOR2_X1 port map( A => n1962, B => 
                           boothmul_pipelined_i_minusA_0_add_0_root_add_22_ni_carry_16_port, Z 
                           => boothmul_pipelined_i_muxes_in_0_119_port);
   U81 : AOI22_X1 port map( A1 => n7140, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n7139, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n5173);
   U82 : OAI21_X1 port map( B1 => n7142, B2 => n1962, A => n5173, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_18_port);
   U83 : AOI222_X1 port map( A1 => n5174, A2 => data1_mul_2_port, B1 => n7140, 
                           B2 => boothmul_pipelined_i_muxes_in_0_115_port, C1 
                           => n7139, C2 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, ZN => 
                           n5176);
   U84 : NOR2_X1 port map( A1 => data2_mul_1_port, A2 => data2_mul_2_port, ZN 
                           => n6911);
   U85 : AOI21_X1 port map( B1 => data2_mul_2_port, B2 => data2_mul_1_port, A 
                           => n6911, ZN => n6871);
   U86 : NAND2_X1 port map( A1 => data1_mul_0_port, A2 => n6871, ZN => n5175);
   U87 : NOR2_X1 port map( A1 => n5176, A2 => n5175, ZN => n3083);
   U88 : AOI21_X1 port map( B1 => n5176, B2 => n5175, A => n3083, ZN => n3086);
   U89 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n5177);
   U90 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, A
                           => n5177, ZN => n6913);
   U91 : NOR3_X1 port map( A1 => n5130, A2 => n6913, A3 => n1990, ZN => n3085);
   U92 : OR2_X1 port map( A1 => n1990, A2 => n6913, ZN => n5178);
   U93 : AOI21_X1 port map( B1 => n5130, B2 => n5178, A => n3085, ZN => n3091);
   U94 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n5179);
   U95 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, A
                           => n5179, ZN => n6953);
   U96 : NOR3_X1 port map( A1 => n3077, A2 => n5124, A3 => n6953, ZN => n3084);
   U97 : AOI221_X1 port map( B1 => n3077, B2 => n5124, C1 => n6953, C2 => n5124
                           , A => n3084, ZN => n3092);
   U98 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n5180);
   U99 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, A
                           => n5180, ZN => n6989);
   U100 : NOR3_X1 port map( A1 => n5121, A2 => n5131, A3 => n6989, ZN => n3090)
                           ;
   U101 : AOI221_X1 port map( B1 => n5121, B2 => n5131, C1 => n6989, C2 => 
                           n5131, A => n3090, ZN => n3093);
   U102 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n5181);
   U103 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, A
                           => n5181, ZN => n7025);
   U104 : NOR3_X1 port map( A1 => n5122, A2 => n5132, A3 => n7025, ZN => n3089)
                           ;
   U105 : AOI221_X1 port map( B1 => n5122, B2 => n5132, C1 => n7025, C2 => 
                           n5132, A => n3089, ZN => n3094);
   U106 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n5182);
   U107 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           A => n5182, ZN => n7061);
   U108 : NOR3_X1 port map( A1 => n5123, A2 => n5133, A3 => n7061, ZN => n3088)
                           ;
   U109 : AOI221_X1 port map( B1 => n5123, B2 => n5133, C1 => n7061, C2 => 
                           n5133, A => n3088, ZN => n3095);
   U110 : INV_X1 port map( A => DATA2(2), ZN => n6865);
   U111 : INV_X1 port map( A => DATA2(4), ZN => n6863);
   U112 : NOR2_X1 port map( A1 => n6865, A2 => n6863, ZN => n5324);
   U113 : INV_X1 port map( A => DATA2(3), ZN => n6864);
   U114 : INV_X1 port map( A => DATA2(5), ZN => n6862);
   U115 : NAND2_X1 port map( A1 => n6863, A2 => n6862, ZN => n6579);
   U116 : INV_X1 port map( A => n6579, ZN => n5894);
   U117 : NOR2_X1 port map( A1 => n6864, A2 => n5894, ZN => n6605);
   U118 : CLKBUF_X1 port map( A => n6605, Z => n6316);
   U119 : NOR2_X1 port map( A1 => n5324, A2 => n6316, ZN => n6590);
   U120 : NAND2_X1 port map( A1 => DATA2(1), A2 => DATA2(0), ZN => n5504);
   U121 : NAND2_X1 port map( A1 => DATA2(3), A2 => DATA2(2), ZN => n5223);
   U122 : OAI21_X1 port map( B1 => n5504, B2 => n5223, A => n5894, ZN => n5183)
                           ;
   U123 : INV_X1 port map( A => n5183, ZN => n6582);
   U124 : INV_X1 port map( A => n6582, ZN => n6410);
   U125 : NAND2_X1 port map( A1 => n6410, A2 => n5894, ZN => n6409);
   U126 : INV_X1 port map( A => DATA2(1), ZN => n6866);
   U127 : OAI21_X1 port map( B1 => n6866, B2 => n5223, A => n5894, ZN => n6072)
                           ;
   U128 : INV_X1 port map( A => DATA2(0), ZN => n6867);
   U129 : NAND2_X1 port map( A1 => n6866, A2 => n6867, ZN => n5412);
   U130 : NOR2_X1 port map( A1 => n6579, A2 => DATA2(3), ZN => n5189);
   U131 : INV_X1 port map( A => n5189, ZN => n5195);
   U132 : NOR2_X1 port map( A1 => n5195, A2 => DATA2(2), ZN => n5691);
   U133 : CLKBUF_X1 port map( A => n5691, Z => n6055);
   U134 : INV_X1 port map( A => n6055, ZN => n5601);
   U135 : OR2_X1 port map( A1 => n5412, A2 => n5601, ZN => n6326);
   U136 : INV_X1 port map( A => n6326, ZN => n5825);
   U137 : AOI22_X1 port map( A1 => DATA1(23), A2 => n5825, B1 => DATA1(27), B2 
                           => n5601, ZN => n5184);
   U138 : INV_X1 port map( A => n5504, ZN => n5371);
   U139 : NAND2_X1 port map( A1 => n5691, A2 => n5371, ZN => n6113);
   U140 : INV_X1 port map( A => n6113, ZN => n6542);
   U141 : CLKBUF_X1 port map( A => n6542, Z => n6058);
   U142 : NAND2_X1 port map( A1 => n6058, A2 => DATA1(26), ZN => n5753);
   U143 : NAND3_X1 port map( A1 => n6867, A2 => DATA2(1), A3 => n5691, ZN => 
                           n6112);
   U144 : INV_X1 port map( A => n6112, ZN => n6097);
   U145 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(25), ZN => n5704);
   U146 : NOR2_X1 port map( A1 => n6867, A2 => DATA2(1), ZN => n5926);
   U147 : NAND2_X1 port map( A1 => n5691, A2 => n5926, ZN => n6283);
   U148 : INV_X1 port map( A => n6283, ZN => n6044);
   U149 : CLKBUF_X1 port map( A => DATA1(24), Z => n6691);
   U150 : NAND2_X1 port map( A1 => n6044, A2 => n6691, ZN => n5692);
   U151 : NAND4_X1 port map( A1 => n5184, A2 => n5753, A3 => n5704, A4 => n5692
                           , ZN => n5243);
   U152 : OAI21_X1 port map( B1 => n6866, B2 => n6865, A => n5189, ZN => n5672)
                           ;
   U153 : INV_X1 port map( A => n6326, ZN => n5185);
   U154 : AOI22_X1 port map( A1 => n6058, A2 => DATA1(24), B1 => n5185, B2 => 
                           DATA1(21), ZN => n5186);
   U155 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(23), ZN => n5693);
   U156 : CLKBUF_X1 port map( A => DATA1(22), Z => n6753);
   U157 : NAND2_X1 port map( A1 => n6044, A2 => n6753, ZN => n5666);
   U158 : NAND2_X1 port map( A1 => DATA1(25), A2 => n5601, ZN => n5754);
   U159 : NAND4_X1 port map( A1 => n5186, A2 => n5693, A3 => n5666, A4 => n5754
                           , ZN => n5198);
   U160 : INV_X1 port map( A => n5672, ZN => n6061);
   U161 : INV_X1 port map( A => n6061, ZN => n6551);
   U162 : AOI21_X1 port map( B1 => DATA2(0), B2 => DATA2(2), A => n6551, ZN => 
                           n6152);
   U163 : INV_X1 port map( A => n6064, ZN => n6549);
   U164 : AOI22_X1 port map( A1 => n6542, A2 => DATA1(25), B1 => n5185, B2 => 
                           n6753, ZN => n5187);
   U165 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(24), ZN => n5710);
   U166 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(23), ZN => n5681);
   U167 : NAND2_X1 port map( A1 => DATA1(26), A2 => n5601, ZN => n5823);
   U168 : NAND4_X1 port map( A1 => n5187, A2 => n5710, A3 => n5681, A4 => n5823
                           , ZN => n5193);
   U169 : NOR4_X1 port map( A1 => n6865, A2 => n6867, A3 => n5195, A4 => 
                           DATA2(1), ZN => n5253);
   U170 : INV_X1 port map( A => n5253, ZN => n6063);
   U171 : INV_X1 port map( A => n6063, ZN => n6547);
   U172 : AOI222_X1 port map( A1 => n5243, A2 => n5672, B1 => n5198, B2 => 
                           n6549, C1 => n5193, C2 => n6547, ZN => n5313);
   U173 : NOR2_X1 port map( A1 => DATA2(2), A2 => DATA2(1), ZN => n5291);
   U174 : CLKBUF_X1 port map( A => n5894, Z => n5983);
   U175 : OAI21_X1 port map( B1 => n5291, B2 => n6864, A => n5983, ZN => n5188)
                           ;
   U176 : INV_X1 port map( A => n5188, ZN => n6561);
   U177 : INV_X1 port map( A => n6561, ZN => n6067);
   U178 : INV_X1 port map( A => n5412, ZN => n5552);
   U179 : OR3_X1 port map( A1 => n6067, A2 => n5552, A3 => n5189, ZN => n6295);
   U180 : NAND3_X1 port map( A1 => n6865, A2 => DATA2(3), A3 => n5983, ZN => 
                           n5228);
   U181 : INV_X1 port map( A => n6232, ZN => n6554);
   U182 : INV_X1 port map( A => DATA1(23), ZN => n6198);
   U183 : NOR2_X1 port map( A1 => n6113, A2 => n6198, ZN => n5707);
   U184 : INV_X1 port map( A => DATA1(24), ZN => n6680);
   U185 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(21), ZN => n5655);
   U186 : NAND2_X1 port map( A1 => n6097, A2 => n6753, ZN => n5682);
   U187 : OAI211_X1 port map( C1 => n6055, C2 => n6680, A => n5655, B => n5682,
                           ZN => n5190);
   U188 : AOI211_X1 port map( C1 => DATA1(20), C2 => n5825, A => n5707, B => 
                           n5190, ZN => n5201);
   U189 : INV_X1 port map( A => n5201, ZN => n5197);
   U190 : AOI222_X1 port map( A1 => n5193, A2 => n5672, B1 => n5197, B2 => 
                           n6152, C1 => n5198, C2 => n5253, ZN => n5299);
   U191 : INV_X1 port map( A => DATA1(26), ZN => n6763);
   U192 : NOR2_X1 port map( A1 => n6112, A2 => n6763, ZN => n5726);
   U193 : INV_X1 port map( A => DATA1(28), ZN => n6768);
   U194 : NAND2_X1 port map( A1 => n5185, A2 => n6691, ZN => n5680);
   U195 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(25), ZN => n5709);
   U196 : OAI211_X1 port map( C1 => n6055, C2 => n6768, A => n5680, B => n5709,
                           ZN => n5191);
   U197 : AOI211_X1 port map( C1 => DATA1(27), C2 => n6058, A => n5726, B => 
                           n5191, ZN => n5192);
   U198 : INV_X1 port map( A => n5192, ZN => n5298);
   U199 : AOI222_X1 port map( A1 => n6549, A2 => n5193, B1 => n6547, B2 => 
                           n5243, C1 => n6551, C2 => n5298, ZN => n5312);
   U200 : OAI22_X1 port map( A1 => n6554, A2 => n5299, B1 => n6561, B2 => n5312
                           , ZN => n5194);
   U201 : INV_X1 port map( A => n5194, ZN => n5203);
   U202 : OAI21_X1 port map( B1 => n5195, B2 => DATA2(0), A => n5672, ZN => 
                           n6197);
   U203 : NOR2_X1 port map( A1 => n5195, A2 => n6197, ZN => n6298);
   U204 : CLKBUF_X1 port map( A => n6298, Z => n6230);
   U205 : AOI22_X1 port map( A1 => n6542, A2 => DATA1(22), B1 => DATA1(19), B2 
                           => n5185, ZN => n5196);
   U206 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(21), ZN => n5667);
   U207 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(20), ZN => n5642);
   U208 : NAND2_X1 port map( A1 => DATA1(23), A2 => n5601, ZN => n5705);
   U209 : NAND4_X1 port map( A1 => n5196, A2 => n5667, A3 => n5642, A4 => n5705
                           , ZN => n5200);
   U210 : AOI222_X1 port map( A1 => n5198, A2 => n5672, B1 => n5200, B2 => 
                           n6152, C1 => n5197, C2 => n5253, ZN => n5244);
   U211 : INV_X1 port map( A => n5244, ZN => n5210);
   U212 : INV_X1 port map( A => DATA1(21), ZN => n6248);
   U213 : NOR2_X1 port map( A1 => n6113, A2 => n6248, ZN => n5679);
   U214 : INV_X1 port map( A => DATA1(22), ZN => n6677);
   U215 : NAND2_X1 port map( A1 => DATA1(19), A2 => n6044, ZN => n5627);
   U216 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(20), ZN => n5656);
   U217 : OAI211_X1 port map( C1 => n6055, C2 => n6677, A => n5627, B => n5656,
                           ZN => n5199);
   U218 : AOI211_X1 port map( C1 => n5185, C2 => DATA1(18), A => n5679, B => 
                           n5199, ZN => n5206);
   U219 : INV_X1 port map( A => n5200, ZN => n5207);
   U220 : OAI222_X1 port map( A1 => n6064, A2 => n5206, B1 => n6063, B2 => 
                           n5207, C1 => n6061, C2 => n5201, ZN => n5216);
   U221 : AOI22_X1 port map( A1 => n6230, A2 => n5210, B1 => n6197, B2 => n5216
                           , ZN => n5202);
   U222 : OAI211_X1 port map( C1 => n5313, C2 => n6295, A => n5203, B => n5202,
                           ZN => n5247);
   U223 : INV_X1 port map( A => n6295, ZN => n6565);
   U224 : INV_X1 port map( A => n5216, ZN => n5225);
   U225 : OAI22_X1 port map( A1 => n6561, A2 => n5299, B1 => n5225, B2 => n6554
                           , ZN => n5209);
   U226 : INV_X1 port map( A => n6197, ZN => n6292);
   U227 : INV_X1 port map( A => n6152, ZN => n6064);
   U228 : INV_X1 port map( A => DATA1(19), ZN => n6340);
   U229 : NOR2_X1 port map( A1 => n6113, A2 => n6340, ZN => n5654);
   U230 : INV_X1 port map( A => DATA1(20), ZN => n6747);
   U231 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(17), ZN => n5591);
   U232 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(18), ZN => n5628);
   U233 : OAI211_X1 port map( C1 => n6055, C2 => n6747, A => n5591, B => n5628,
                           ZN => n5204);
   U234 : AOI211_X1 port map( C1 => n5185, C2 => DATA1(16), A => n5654, B => 
                           n5204, ZN => n5218);
   U235 : NOR2_X1 port map( A1 => n6113, A2 => n6747, ZN => n5665);
   U236 : NAND2_X1 port map( A1 => DATA1(18), A2 => n6044, ZN => n5616);
   U237 : NAND2_X1 port map( A1 => DATA1(19), A2 => n6097, ZN => n5643);
   U238 : OAI211_X1 port map( C1 => n5691, C2 => n6248, A => n5616, B => n5643,
                           ZN => n5205);
   U239 : AOI211_X1 port map( C1 => DATA1(17), C2 => n5825, A => n5665, B => 
                           n5205, ZN => n5215);
   U240 : OAI222_X1 port map( A1 => n6064, A2 => n5218, B1 => n6063, B2 => 
                           n5215, C1 => n6061, C2 => n5206, ZN => n5258);
   U241 : INV_X1 port map( A => n5258, ZN => n5236);
   U242 : OAI222_X1 port map( A1 => n5207, A2 => n6061, B1 => n5215, B2 => 
                           n6064, C1 => n5206, C2 => n6063, ZN => n5219);
   U243 : INV_X1 port map( A => n5219, ZN => n5235);
   U244 : INV_X1 port map( A => n6298, ZN => n6181);
   U245 : CLKBUF_X1 port map( A => n6181, Z => n6558);
   U246 : OAI22_X1 port map( A1 => n6292, A2 => n5236, B1 => n5235, B2 => n6558
                           , ZN => n5208);
   U247 : AOI211_X1 port map( C1 => n6565, C2 => n5210, A => n5209, B => n5208,
                           ZN => n5302);
   U248 : INV_X1 port map( A => n5223, ZN => n5213);
   U249 : NAND3_X1 port map( A1 => n5983, A2 => n5552, A3 => n5213, ZN => n6568
                           );
   U250 : INV_X1 port map( A => n6568, ZN => n6468);
   U251 : INV_X1 port map( A => n6468, ZN => n6451);
   U252 : OAI22_X1 port map( A1 => n5244, A2 => n6554, B1 => n5299, B2 => n6295
                           , ZN => n5212);
   U253 : OAI22_X1 port map( A1 => n6561, A2 => n5313, B1 => n5225, B2 => n6558
                           , ZN => n5211);
   U254 : AOI211_X1 port map( C1 => n6197, C2 => n5219, A => n5212, B => n5211,
                           ZN => n5316);
   U255 : INV_X1 port map( A => n6072, ZN => n6573);
   U256 : NAND3_X1 port map( A1 => DATA2(0), A2 => n5213, A3 => n6573, ZN => 
                           n6450);
   U257 : OAI22_X1 port map( A1 => n5302, A2 => n6451, B1 => n5316, B2 => n6450
                           , ZN => n5230);
   U258 : INV_X1 port map( A => DATA1(17), ZN => n6375);
   U259 : NOR2_X1 port map( A1 => n6112, A2 => n6375, ZN => n5615);
   U260 : INV_X1 port map( A => DATA1(15), ZN => n6403);
   U261 : NAND2_X1 port map( A1 => DATA1(16), A2 => n6044, ZN => n5594);
   U262 : NAND2_X1 port map( A1 => DATA1(19), A2 => n5601, ZN => n5669);
   U263 : OAI211_X1 port map( C1 => n6403, C2 => n6326, A => n5594, B => n5669,
                           ZN => n5214);
   U264 : AOI211_X1 port map( C1 => DATA1(18), C2 => n6058, A => n5615, B => 
                           n5214, ZN => n5231);
   U265 : OAI222_X1 port map( A1 => n6063, A2 => n5218, B1 => n6064, B2 => 
                           n5231, C1 => n6061, C2 => n5215, ZN => n5269);
   U266 : AOI22_X1 port map( A1 => n6298, A2 => n5269, B1 => n6067, B2 => n5216
                           , ZN => n5221);
   U267 : NOR2_X1 port map( A1 => n6283, A2 => n6403, ZN => n5600);
   U268 : INV_X1 port map( A => n7169, ZN => n6427);
   U269 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(16), ZN => n5590);
   U270 : NAND2_X1 port map( A1 => DATA1(18), A2 => n5601, ZN => n5652);
   U271 : OAI211_X1 port map( C1 => n6326, C2 => n6427, A => n5590, B => n5652,
                           ZN => n5217);
   U272 : AOI211_X1 port map( C1 => DATA1(17), C2 => n6058, A => n5600, B => 
                           n5217, ZN => n5233);
   U273 : OAI222_X1 port map( A1 => n6064, A2 => n5233, B1 => n6063, B2 => 
                           n5231, C1 => n6061, C2 => n5218, ZN => n5265);
   U274 : AOI22_X1 port map( A1 => n6565, A2 => n5219, B1 => n5265, B2 => n6197
                           , ZN => n5220);
   U275 : OAI211_X1 port map( C1 => n5236, C2 => n6554, A => n5221, B => n5220,
                           ZN => n5222);
   U276 : INV_X1 port map( A => n5222, ZN => n5286);
   U277 : OAI211_X1 port map( C1 => n6864, C2 => n5504, A => n5223, B => n5983,
                           ZN => n5224);
   U278 : INV_X1 port map( A => n5224, ZN => n6526);
   U279 : INV_X1 port map( A => n5269, ZN => n5255);
   U280 : OAI22_X1 port map( A1 => n6561, A2 => n5244, B1 => n6292, B2 => n5255
                           , ZN => n5227);
   U281 : OAI22_X1 port map( A1 => n5235, A2 => n6554, B1 => n5225, B2 => n6295
                           , ZN => n5226);
   U282 : AOI211_X1 port map( C1 => n6230, C2 => n5258, A => n5227, B => n5226,
                           ZN => n5287);
   U283 : NOR2_X1 port map( A1 => n5504, A2 => n5228, ZN => n6073);
   U284 : INV_X1 port map( A => n6073, ZN => n6570);
   U285 : OAI22_X1 port map( A1 => n5286, A2 => n5224, B1 => n5287, B2 => n6570
                           , ZN => n5229);
   U286 : AOI211_X1 port map( C1 => n6072, C2 => n5247, A => n5230, B => n5229,
                           ZN => n5306);
   U287 : INV_X1 port map( A => n5287, ZN => n5241);
   U288 : INV_X1 port map( A => n5231, ZN => n5234);
   U289 : AOI22_X1 port map( A1 => DATA1(13), A2 => n5825, B1 => DATA1(17), B2 
                           => n5601, ZN => n5232);
   U290 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(14), ZN => n5608);
   U291 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(15), ZN => n5593);
   U292 : NAND2_X1 port map( A1 => n6058, A2 => DATA1(16), ZN => n5618);
   U293 : NAND4_X1 port map( A1 => n5232, A2 => n5608, A3 => n5593, A4 => n5618
                           , ZN => n5262);
   U294 : INV_X1 port map( A => n5233, ZN => n5254);
   U295 : AOI222_X1 port map( A1 => n5234, A2 => n6551, B1 => n5262, B2 => 
                           n6152, C1 => n5254, C2 => n6547, ZN => n5279);
   U296 : OAI22_X1 port map( A1 => n6561, A2 => n5235, B1 => n6292, B2 => n5279
                           , ZN => n5238);
   U297 : INV_X1 port map( A => n5265, ZN => n5266);
   U298 : OAI22_X1 port map( A1 => n5266, A2 => n6558, B1 => n5236, B2 => n6295
                           , ZN => n5237);
   U299 : AOI211_X1 port map( C1 => n6232, C2 => n5269, A => n5238, B => n5237,
                           ZN => n5285);
   U300 : INV_X1 port map( A => n6526, ZN => n6566);
   U301 : OAI22_X1 port map( A1 => n6573, A2 => n5316, B1 => n5285, B2 => n6566
                           , ZN => n5240);
   U302 : OAI22_X1 port map( A1 => n5286, A2 => n6570, B1 => n5302, B2 => n6450
                           , ZN => n5239);
   U303 : AOI211_X1 port map( C1 => n6468, C2 => n5241, A => n5240, B => n5239,
                           ZN => n5294);
   U304 : INV_X1 port map( A => n5316, ZN => n5250);
   U305 : INV_X1 port map( A => n5312, ZN => n6227);
   U306 : AOI22_X1 port map( A1 => DATA1(25), A2 => n5825, B1 => DATA1(29), B2 
                           => n5601, ZN => n5242);
   U307 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(27), ZN => n5752);
   U308 : NAND2_X1 port map( A1 => n6058, A2 => DATA1(28), ZN => n5933);
   U309 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(26), ZN => n5703);
   U310 : NAND4_X1 port map( A1 => n5242, A2 => n5752, A3 => n5933, A4 => n5703
                           , ZN => n5310);
   U311 : AOI222_X1 port map( A1 => n5310, A2 => n5672, B1 => n5243, B2 => 
                           n6152, C1 => n5298, C2 => n5253, ZN => n5311);
   U312 : OAI22_X1 port map( A1 => n6561, A2 => n5311, B1 => n5313, B2 => n6554
                           , ZN => n5246);
   U313 : CLKBUF_X1 port map( A => n6292, Z => n6557);
   U314 : OAI22_X1 port map( A1 => n6557, A2 => n5244, B1 => n5299, B2 => n6181
                           , ZN => n5245);
   U315 : AOI211_X1 port map( C1 => n6565, C2 => n6227, A => n5246, B => n5245,
                           ZN => n6357);
   U316 : INV_X1 port map( A => n5247, ZN => n6358);
   U317 : OAI22_X1 port map( A1 => n6573, A2 => n6357, B1 => n6358, B2 => n6450
                           , ZN => n5249);
   U318 : OAI22_X1 port map( A1 => n5287, A2 => n5224, B1 => n5302, B2 => n6570
                           , ZN => n5248);
   U319 : AOI211_X1 port map( C1 => n6468, C2 => n5250, A => n5249, B => n5248,
                           ZN => n5320);
   U320 : OAI222_X1 port map( A1 => n6409, A2 => n5306, B1 => n6410, B2 => 
                           n5294, C1 => n5320, C2 => n5983, ZN => n6474);
   U321 : INV_X1 port map( A => n6474, ZN => n5323);
   U322 : NOR2_X1 port map( A1 => DATA2(2), A2 => n5412, ZN => n5251);
   U323 : AOI21_X1 port map( B1 => n5251, B2 => n6864, A => n5894, ZN => n6307)
                           ;
   U324 : CLKBUF_X1 port map( A => n6307, Z => n6588);
   U325 : INV_X1 port map( A => n6588, ZN => n6472);
   U326 : AOI22_X1 port map( A1 => DATA1(12), A2 => n5825, B1 => DATA1(16), B2 
                           => n5601, ZN => n5252);
   U327 : NAND2_X1 port map( A1 => n6058, A2 => DATA1(15), ZN => n5589);
   U328 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(13), ZN => n5612);
   U329 : NAND2_X1 port map( A1 => n6097, A2 => n7169, ZN => n5597);
   U330 : NAND4_X1 port map( A1 => n5252, A2 => n5589, A3 => n5612, A4 => n5597
                           , ZN => n5261);
   U331 : AOI222_X1 port map( A1 => n5254, A2 => n6551, B1 => n5261, B2 => 
                           n6152, C1 => n5262, C2 => n5253, ZN => n5275);
   U332 : OAI22_X1 port map( A1 => n6557, A2 => n5275, B1 => n5266, B2 => n6554
                           , ZN => n5257);
   U333 : OAI22_X1 port map( A1 => n5279, A2 => n6181, B1 => n5255, B2 => n6295
                           , ZN => n5256);
   U334 : AOI211_X1 port map( C1 => n6067, C2 => n5258, A => n5257, B => n5256,
                           ZN => n5381);
   U335 : INV_X1 port map( A => n5381, ZN => n5284);
   U336 : AOI22_X1 port map( A1 => DATA1(10), A2 => n5825, B1 => DATA1(14), B2 
                           => n5601, ZN => n5259);
   U337 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(11), ZN => n5636);
   U338 : NAND2_X1 port map( A1 => n6058, A2 => DATA1(13), ZN => n5598);
   U339 : NAND2_X1 port map( A1 => n6097, A2 => n7168, ZN => n5611);
   U340 : NAND4_X1 port map( A1 => n5259, A2 => n5636, A3 => n5598, A4 => n5611
                           , ZN => n5374);
   U341 : AOI22_X1 port map( A1 => n7169, A2 => n6542, B1 => DATA1(15), B2 => 
                           n5601, ZN => n5260);
   U342 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(12), ZN => n5604);
   U343 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(13), ZN => n5607);
   U344 : CLKBUF_X1 port map( A => DATA1(11), Z => n6000);
   U345 : NAND2_X1 port map( A1 => n5825, A2 => n6000, ZN => n5770);
   U346 : NAND4_X1 port map( A1 => n5260, A2 => n5604, A3 => n5607, A4 => n5770
                           , ZN => n5273);
   U347 : AOI222_X1 port map( A1 => n5261, A2 => n5672, B1 => n5374, B2 => 
                           n6549, C1 => n5273, C2 => n6547, ZN => n5447);
   U348 : OAI22_X1 port map( A1 => n5275, A2 => n6554, B1 => n6557, B2 => n5447
                           , ZN => n5264);
   U349 : AOI222_X1 port map( A1 => n5262, A2 => n6551, B1 => n5273, B2 => 
                           n6549, C1 => n5261, C2 => n6547, ZN => n5276);
   U350 : OAI22_X1 port map( A1 => n5279, A2 => n6295, B1 => n5276, B2 => n6181
                           , ZN => n5263);
   U351 : AOI211_X1 port map( C1 => n6067, C2 => n5265, A => n5264, B => n5263,
                           ZN => n5450);
   U352 : OAI22_X1 port map( A1 => n6566, A2 => n5450, B1 => n6573, B2 => n5286
                           , ZN => n5271);
   U353 : OAI22_X1 port map( A1 => n5279, A2 => n6554, B1 => n5276, B2 => n6292
                           , ZN => n5268);
   U354 : OAI22_X1 port map( A1 => n5266, A2 => n6295, B1 => n5275, B2 => n6181
                           , ZN => n5267);
   U355 : AOI211_X1 port map( C1 => n6067, C2 => n5269, A => n5268, B => n5267,
                           ZN => n5421);
   U356 : OAI22_X1 port map( A1 => n6450, A2 => n5285, B1 => n6570, B2 => n5421
                           , ZN => n5270);
   U357 : AOI211_X1 port map( C1 => n5284, C2 => n6468, A => n5271, B => n5270,
                           ZN => n5384);
   U358 : INV_X1 port map( A => n6450, ZN => n6577);
   U359 : INV_X1 port map( A => n5447, ZN => n5376);
   U360 : INV_X1 port map( A => DATA1(10), ZN => n6662);
   U361 : NOR2_X1 port map( A1 => n6283, A2 => n6662, ZN => n5773);
   U362 : INV_X1 port map( A => DATA1(13), ZN => n6447);
   U363 : NAND2_X1 port map( A1 => n5185, A2 => DATA1(9), ZN => n5344);
   U364 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(11), ZN => n5603);
   U365 : OAI211_X1 port map( C1 => n6055, C2 => n6447, A => n5344, B => n5603,
                           ZN => n5272);
   U366 : AOI211_X1 port map( C1 => n7168, C2 => n6542, A => n5773, B => n5272,
                           ZN => n5417);
   U367 : INV_X1 port map( A => n5417, ZN => n5274);
   U368 : AOI222_X1 port map( A1 => n6549, A2 => n5274, B1 => n6547, B2 => 
                           n5374, C1 => n6551, C2 => n5273, ZN => n5380);
   U369 : INV_X1 port map( A => n5380, ZN => n5485);
   U370 : AOI22_X1 port map( A1 => n6230, A2 => n5376, B1 => n6197, B2 => n5485
                           , ZN => n5278);
   U371 : INV_X1 port map( A => n5275, ZN => n5377);
   U372 : INV_X1 port map( A => n5276, ZN => n5418);
   U373 : AOI22_X1 port map( A1 => n6565, A2 => n5377, B1 => n6232, B2 => n5418
                           , ZN => n5277);
   U374 : OAI211_X1 port map( C1 => n6561, C2 => n5279, A => n5278, B => n5277,
                           ZN => n5488);
   U375 : INV_X1 port map( A => n5488, ZN => n5413);
   U376 : OAI22_X1 port map( A1 => n5413, A2 => n6566, B1 => n5421, B2 => n6451
                           , ZN => n5281);
   U377 : OAI22_X1 port map( A1 => n6573, A2 => n5285, B1 => n5450, B2 => n6570
                           , ZN => n5280);
   U378 : AOI211_X1 port map( C1 => n6577, C2 => n5284, A => n5281, B => n5280,
                           ZN => n5425);
   U379 : CLKBUF_X1 port map( A => n6073, Z => n6495);
   U380 : OAI22_X1 port map( A1 => n5421, A2 => n6566, B1 => n5286, B2 => n6450
                           , ZN => n5283);
   U381 : OAI22_X1 port map( A1 => n6573, A2 => n5287, B1 => n5285, B2 => n6451
                           , ZN => n5282);
   U382 : AOI211_X1 port map( C1 => n6495, C2 => n5284, A => n5283, B => n5282,
                           ZN => n5292);
   U383 : OAI222_X1 port map( A1 => n6409, A2 => n5384, B1 => n6410, B2 => 
                           n5425, C1 => n5292, C2 => n5894, ZN => n5498);
   U384 : INV_X1 port map( A => n6590, ZN => n5985);
   U385 : NOR4_X1 port map( A1 => n5894, A2 => n5291, A3 => n5371, A4 => n5985,
                           ZN => n5908);
   U386 : CLKBUF_X1 port map( A => n5908, Z => n6470);
   U387 : INV_X1 port map( A => n5285, ZN => n5290);
   U388 : OAI22_X1 port map( A1 => n5381, A2 => n6566, B1 => n5286, B2 => n6451
                           , ZN => n5289);
   U389 : OAI22_X1 port map( A1 => n6573, A2 => n5302, B1 => n5287, B2 => n6450
                           , ZN => n5288);
   U390 : AOI211_X1 port map( C1 => n6073, C2 => n5290, A => n5289, B => n5288,
                           ZN => n5293);
   U391 : OAI222_X1 port map( A1 => n6409, A2 => n5293, B1 => n6410, B2 => 
                           n5292, C1 => n5294, C2 => n5894, ZN => n5426);
   U392 : AOI22_X1 port map( A1 => n6472, A2 => n5498, B1 => n6470, B2 => n5426
                           , ZN => n5296);
   U393 : INV_X1 port map( A => n6605, ZN => n6081);
   U394 : NAND3_X1 port map( A1 => n5291, A2 => n6081, A3 => n6588, ZN => n6592
                           );
   U395 : INV_X1 port map( A => n6592, ZN => n6475);
   U396 : OAI222_X1 port map( A1 => n6409, A2 => n5292, B1 => n6410, B2 => 
                           n5384, C1 => n5293, C2 => n5894, ZN => n5455);
   U397 : NAND3_X1 port map( A1 => DATA2(4), A2 => n6590, A3 => n5371, ZN => 
                           n6310);
   U398 : INV_X1 port map( A => n6310, ZN => n6595);
   U399 : OAI222_X1 port map( A1 => n6409, A2 => n5294, B1 => n6410, B2 => 
                           n5293, C1 => n5306, C2 => n5894, ZN => n6471);
   U400 : AOI22_X1 port map( A1 => n6475, A2 => n5455, B1 => n6595, B2 => n6471
                           , ZN => n5295);
   U401 : OAI211_X1 port map( C1 => n6590, C2 => n5323, A => n5296, B => n5295,
                           ZN => n5478);
   U402 : OAI21_X1 port map( B1 => n5412, B2 => n6316, A => n5985, ZN => n6509)
                           ;
   U403 : INV_X1 port map( A => n6357, ZN => n5305);
   U404 : INV_X1 port map( A => n5311, ZN => n6229);
   U405 : INV_X1 port map( A => DATA1(29), ZN => n6095);
   U406 : INV_X1 port map( A => n5691, ZN => n5785);
   U407 : NOR2_X1 port map( A1 => n6326, A2 => n6763, ZN => n5708);
   U408 : INV_X1 port map( A => DATA1(27), ZN => n6136);
   U409 : NOR2_X1 port map( A1 => n6283, A2 => n6136, ZN => n5725);
   U410 : AOI211_X1 port map( C1 => DATA1(30), C2 => n5785, A => n5708, B => 
                           n5725, ZN => n5297);
   U411 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(28), ZN => n5822);
   U412 : OAI211_X1 port map( C1 => n6095, C2 => n6113, A => n5297, B => n5822,
                           ZN => n6151);
   U413 : AOI222_X1 port map( A1 => n6151, A2 => n6551, B1 => n5298, B2 => 
                           n6549, C1 => n5310, C2 => n6547, ZN => n6182);
   U414 : OAI22_X1 port map( A1 => n6561, A2 => n6182, B1 => n5312, B2 => n6554
                           , ZN => n5301);
   U415 : OAI22_X1 port map( A1 => n6557, A2 => n5299, B1 => n5313, B2 => n6181
                           , ZN => n5300);
   U416 : AOI211_X1 port map( C1 => n6565, C2 => n6229, A => n5301, B => n5300,
                           ZN => n6360);
   U417 : OAI22_X1 port map( A1 => n6573, A2 => n6360, B1 => n5316, B2 => n6570
                           , ZN => n5304);
   U418 : OAI22_X1 port map( A1 => n5302, A2 => n6566, B1 => n6358, B2 => n6451
                           , ZN => n5303);
   U419 : AOI211_X1 port map( C1 => n6577, C2 => n5305, A => n5304, B => n5303,
                           ZN => n6392);
   U420 : OAI222_X1 port map( A1 => n6409, A2 => n5320, B1 => n6410, B2 => 
                           n5306, C1 => n6392, C2 => n5894, ZN => n6469);
   U421 : AOI22_X1 port map( A1 => n6595, A2 => n6474, B1 => n5985, B2 => n6469
                           , ZN => n5308);
   U422 : AOI22_X1 port map( A1 => n6475, A2 => n5426, B1 => n6470, B2 => n6471
                           , ZN => n5307);
   U423 : NAND2_X1 port map( A1 => n5308, A2 => n5307, ZN => n5456);
   U424 : AOI21_X1 port map( B1 => n6472, B2 => n5455, A => n5456, ZN => n5431)
                           ;
   U425 : INV_X1 port map( A => n5431, ZN => n6515);
   U426 : NAND3_X1 port map( A1 => n6864, A2 => n5324, A3 => n5926, ZN => n6608
                           );
   U427 : INV_X1 port map( A => n6608, ZN => n6518);
   U428 : INV_X1 port map( A => n5908, ZN => n6586);
   U429 : INV_X1 port map( A => n6360, ZN => n5319);
   U430 : INV_X1 port map( A => n6182, ZN => n6231);
   U431 : INV_X1 port map( A => DATA1(31), ZN => n6689);
   U432 : NOR2_X1 port map( A1 => n6112, A2 => n6095, ZN => n5932);
   U433 : NOR2_X1 port map( A1 => n6283, A2 => n6768, ZN => n5756);
   U434 : AOI211_X1 port map( C1 => DATA1(30), C2 => n6542, A => n5932, B => 
                           n5756, ZN => n5309);
   U435 : NAND2_X1 port map( A1 => n5825, A2 => DATA1(27), ZN => n5702);
   U436 : OAI211_X1 port map( C1 => n6055, C2 => n6689, A => n5309, B => n5702,
                           ZN => n6150);
   U437 : AOI222_X1 port map( A1 => n6150, A2 => n5672, B1 => n5310, B2 => 
                           n6549, C1 => n6151, C2 => n6547, ZN => n6196);
   U438 : OAI22_X1 port map( A1 => n6561, A2 => n6196, B1 => n5311, B2 => n6554
                           , ZN => n5315);
   U439 : OAI22_X1 port map( A1 => n6557, A2 => n5313, B1 => n5312, B2 => n6181
                           , ZN => n5314);
   U440 : AOI211_X1 port map( C1 => n6565, C2 => n6231, A => n5315, B => n5314,
                           ZN => n6359);
   U441 : OAI22_X1 port map( A1 => n6573, A2 => n6359, B1 => n6357, B2 => n6568
                           , ZN => n5318);
   U442 : OAI22_X1 port map( A1 => n5316, A2 => n5224, B1 => n6358, B2 => n6570
                           , ZN => n5317);
   U443 : AOI211_X1 port map( C1 => n6577, C2 => n5319, A => n5318, B => n5317,
                           ZN => n6391);
   U444 : OAI222_X1 port map( A1 => n6409, A2 => n6392, B1 => n6410, B2 => 
                           n5320, C1 => n6391, C2 => n5894, ZN => n6473);
   U445 : AOI22_X1 port map( A1 => n6472, A2 => n5426, B1 => n5985, B2 => n6473
                           , ZN => n5322);
   U446 : AOI22_X1 port map( A1 => n6475, A2 => n6471, B1 => n6595, B2 => n6469
                           , ZN => n5321);
   U447 : OAI211_X1 port map( C1 => n5323, C2 => n6586, A => n5322, B => n5321,
                           ZN => n6517);
   U448 : INV_X1 port map( A => n5324, ZN => n5369);
   U449 : NOR4_X1 port map( A1 => n6866, A2 => n5369, A3 => n6316, A4 => 
                           DATA2(0), ZN => n6315);
   U450 : CLKBUF_X1 port map( A => n6315, Z => n6236);
   U451 : AOI222_X1 port map( A1 => n5478, A2 => n6509, B1 => n6515, B2 => 
                           n6518, C1 => n6517, C2 => n6236, ZN => n5368);
   U452 : NOR2_X1 port map( A1 => n6864, A2 => n5369, ZN => n5927);
   U453 : NAND2_X1 port map( A1 => n5927, A2 => DATA2(1), ZN => n6622);
   U454 : INV_X1 port map( A => n6622, ZN => n5326);
   U455 : NOR2_X1 port map( A1 => DATA2(5), A2 => FUNC(0), ZN => n5325);
   U456 : NAND3_X1 port map( A1 => n5325, A2 => FUNC(2), A3 => FUNC(1), ZN => 
                           n5999);
   U457 : AOI21_X1 port map( B1 => DATA2(0), B2 => n5326, A => n5999, ZN => 
                           n5357);
   U458 : NAND2_X1 port map( A1 => FUNC(3), A2 => n5357, ZN => n6830);
   U459 : NOR4_X1 port map( A1 => DATA2(9), A2 => DATA2(8), A3 => DATA2(6), A4 
                           => DATA2(7), ZN => n5334);
   U460 : INV_X1 port map( A => DATA2(12), ZN => n6853);
   U461 : INV_X1 port map( A => DATA2(10), ZN => n6855);
   U462 : INV_X1 port map( A => DATA2(11), ZN => n6854);
   U463 : INV_X1 port map( A => DATA2(13), ZN => n6852);
   U464 : NAND4_X1 port map( A1 => n6853, A2 => n6855, A3 => n6854, A4 => n6852
                           , ZN => n5327);
   U465 : NOR4_X1 port map( A1 => DATA2(14), A2 => DATA2(15), A3 => n6326, A4 
                           => n5327, ZN => n5333);
   U466 : NOR4_X1 port map( A1 => DATA1(15), A2 => DATA1(14), A3 => DATA1(13), 
                           A4 => DATA1(12), ZN => n5331);
   U467 : CLKBUF_X1 port map( A => DATA1(8), Z => n5774);
   U468 : NOR4_X1 port map( A1 => n6000, A2 => DATA1(10), A3 => DATA1(9), A4 =>
                           n5774, ZN => n5330);
   U469 : CLKBUF_X1 port map( A => DATA1(5), Z => n6059);
   U470 : NOR4_X1 port map( A1 => DATA1(7), A2 => DATA1(6), A3 => n6059, A4 => 
                           DATA1(4), ZN => n5329);
   U471 : NOR4_X1 port map( A1 => DATA1(3), A2 => DATA1(2), A3 => DATA1(1), A4 
                           => DATA1(0), ZN => n5328);
   U472 : AND4_X1 port map( A1 => n5331, A2 => n5330, A3 => n5329, A4 => n5328,
                           ZN => n5332);
   U473 : AOI211_X1 port map( C1 => n5334, C2 => n5333, A => n5332, B => n553, 
                           ZN => n6183);
   U474 : CLKBUF_X1 port map( A => n6183, Z => n6641);
   U475 : NOR2_X1 port map( A1 => DATA1(8), A2 => DATA2_I_8_port, ZN => n5389);
   U476 : XOR2_X1 port map( A => DATA2_I_9_port, B => DATA1(9), Z => n5365);
   U477 : INV_X1 port map( A => n5365, ZN => n6002);
   U478 : NOR2_X1 port map( A1 => n5389, A2 => n6002, ZN => n6537);
   U479 : INV_X1 port map( A => n1992, ZN => n6833);
   U480 : NAND2_X1 port map( A1 => DATA1(7), A2 => DATA2_I_7_port, ZN => n5340)
                           ;
   U481 : OAI21_X1 port map( B1 => DATA1(7), B2 => DATA2_I_7_port, A => n5340, 
                           ZN => n5434);
   U482 : NAND2_X1 port map( A1 => DATA1(6), A2 => DATA2_I_6_port, ZN => n5407)
                           ;
   U483 : NAND2_X1 port map( A1 => DATA1(5), A2 => DATA2_I_5_port, ZN => n5337)
                           ;
   U484 : INV_X1 port map( A => n5337, ZN => n5406);
   U485 : XOR2_X1 port map( A => DATA2_I_3_port, B => DATA1(3), Z => n5587);
   U486 : NAND2_X1 port map( A1 => DATA1(2), A2 => DATA2_I_2_port, ZN => n5403)
                           ;
   U487 : OAI21_X1 port map( B1 => DATA1(2), B2 => DATA2_I_2_port, A => n5403, 
                           ZN => n6048);
   U488 : NAND2_X1 port map( A1 => DATA1(1), A2 => DATA2_I_1_port, ZN => n5401)
                           ;
   U489 : NAND2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n6630)
                           ;
   U490 : INV_X1 port map( A => n6630, ZN => n6280);
   U491 : NOR2_X1 port map( A1 => DATA1(0), A2 => DATA2_I_0_port, ZN => n6277);
   U492 : OAI21_X1 port map( B1 => DATA1(1), B2 => DATA2_I_1_port, A => n5401, 
                           ZN => n6278);
   U493 : NOR2_X1 port map( A1 => n6277, A2 => n6278, ZN => n6276);
   U494 : OAI21_X1 port map( B1 => n6280, B2 => cin, A => n6276, ZN => n5335);
   U495 : OAI221_X1 port map( B1 => n6048, B2 => n5401, C1 => n6048, C2 => 
                           n5335, A => n5403, ZN => n5336);
   U496 : AND2_X1 port map( A1 => DATA1(3), A2 => DATA2_I_3_port, ZN => n5404);
   U497 : AOI21_X1 port map( B1 => n5587, B2 => n5336, A => n5404, ZN => n5338)
                           ;
   U498 : NAND2_X1 port map( A1 => DATA1(4), A2 => DATA2_I_4_port, ZN => n5405)
                           ;
   U499 : OAI21_X1 port map( B1 => DATA1(4), B2 => DATA2_I_4_port, A => n5405, 
                           ZN => n5547);
   U500 : OAI21_X1 port map( B1 => n6059, B2 => DATA2_I_5_port, A => n5337, ZN 
                           => n5508);
   U501 : AOI221_X1 port map( B1 => n5338, B2 => n5405, C1 => n5547, C2 => 
                           n5405, A => n5508, ZN => n5339);
   U502 : XOR2_X1 port map( A => DATA2_I_6_port, B => DATA1(6), Z => n5468);
   U503 : OAI21_X1 port map( B1 => n5406, B2 => n5339, A => n5468, ZN => n5341)
                           ;
   U504 : OAI221_X1 port map( B1 => n5434, B2 => n5407, C1 => n5434, C2 => 
                           n5341, A => n5340, ZN => n6457);
   U505 : NAND2_X1 port map( A1 => n6833, A2 => n6457, ZN => n5390);
   U506 : AOI211_X1 port map( C1 => n5389, C2 => n6002, A => n6537, B => n5390,
                           ZN => n5363);
   U507 : INV_X1 port map( A => DATA1(9), ZN => n5481);
   U508 : NOR2_X1 port map( A1 => n5481, A2 => DATA2(9), ZN => n6717);
   U509 : INV_X1 port map( A => n6717, ZN => n6661);
   U510 : NAND2_X1 port map( A1 => DATA2(9), A2 => n5481, ZN => n6718);
   U511 : AND2_X1 port map( A1 => n6661, A2 => n6718, ZN => n6787);
   U512 : INV_X1 port map( A => FUNC(0), ZN => n5342);
   U513 : NAND3_X1 port map( A1 => n5342, A2 => n6773, A3 => FUNC(1), ZN => 
                           n6492);
   U514 : INV_X1 port map( A => n6492, ZN => n6631);
   U515 : INV_X1 port map( A => n6631, ZN => n6531);
   U516 : NAND2_X1 port map( A1 => FUNC(3), A2 => n5343, ZN => n6389);
   U517 : NOR2_X1 port map( A1 => n6492, A2 => FUNC(3), ZN => n6493);
   U518 : INV_X1 port map( A => n6493, ZN => n6388);
   U519 : NAND2_X1 port map( A1 => n6389, A2 => n6388, ZN => n6528);
   U520 : NAND3_X1 port map( A1 => DATA2(9), A2 => DATA1(9), A3 => n6528, ZN =>
                           n5361);
   U521 : INV_X1 port map( A => DATA1(8), ZN => n6715);
   U522 : NOR2_X1 port map( A1 => n6283, A2 => n6715, ZN => n5416);
   U523 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(7), ZN => n5480);
   U524 : NAND2_X1 port map( A1 => n6058, A2 => DATA1(6), ZN => n5555);
   U525 : NAND2_X1 port map( A1 => n6059, A2 => n5601, ZN => n6285);
   U526 : NAND4_X1 port map( A1 => n5344, A2 => n5480, A3 => n5555, A4 => n6285
                           , ZN => n5345);
   U527 : NOR2_X1 port map( A1 => n5416, A2 => n5345, ZN => n5849);
   U528 : INV_X1 port map( A => DATA1(7), ZN => n5782);
   U529 : NOR2_X1 port map( A1 => n6283, A2 => n5782, ZN => n5443);
   U530 : INV_X1 port map( A => DATA1(6), ZN => n6695);
   U531 : NOR2_X1 port map( A1 => n6112, A2 => n6695, ZN => n5522);
   U532 : AOI211_X1 port map( C1 => n6058, C2 => DATA1(5), A => n5443, B => 
                           n5522, ZN => n5346);
   U533 : NAND2_X1 port map( A1 => n5185, A2 => n5774, ZN => n5372);
   U534 : NAND2_X1 port map( A1 => DATA1(4), A2 => n5785, ZN => n6543);
   U535 : AND3_X1 port map( A1 => n5346, A2 => n5372, A3 => n6543, ZN => n5851)
                           ;
   U536 : NOR2_X1 port map( A1 => n6283, A2 => n6695, ZN => n5483);
   U537 : INV_X1 port map( A => DATA1(3), ZN => n5577);
   U538 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(5), ZN => n5553);
   U539 : NAND2_X1 port map( A1 => n5825, A2 => DATA1(7), ZN => n5414);
   U540 : OAI211_X1 port map( C1 => n6055, C2 => n5577, A => n5553, B => n5414,
                           ZN => n5347);
   U541 : AOI211_X1 port map( C1 => n6058, C2 => DATA1(4), A => n5483, B => 
                           n5347, ZN => n5351);
   U542 : OAI222_X1 port map( A1 => n6064, A2 => n5849, B1 => n6063, B2 => 
                           n5851, C1 => n6061, C2 => n5351, ZN => n5885);
   U543 : INV_X1 port map( A => n5885, ZN => n5975);
   U544 : INV_X1 port map( A => DATA1(4), ZN => n5514);
   U545 : NOR2_X1 port map( A1 => n6112, A2 => n5514, ZN => n6057);
   U546 : INV_X1 port map( A => DATA1(2), ZN => n6648);
   U547 : NAND2_X1 port map( A1 => n6044, A2 => n6059, ZN => n5520);
   U548 : NAND2_X1 port map( A1 => n5185, A2 => DATA1(6), ZN => n5441);
   U549 : OAI211_X1 port map( C1 => n5691, C2 => n6648, A => n5520, B => n5441,
                           ZN => n5348);
   U550 : AOI211_X1 port map( C1 => DATA1(3), C2 => n6542, A => n6057, B => 
                           n5348, ZN => n5352);
   U551 : OAI222_X1 port map( A1 => n6064, A2 => n5851, B1 => n6063, B2 => 
                           n5351, C1 => n6061, C2 => n5352, ZN => n5903);
   U552 : INV_X1 port map( A => n5903, ZN => n5973);
   U553 : OAI22_X1 port map( A1 => n6557, A2 => n5975, B1 => n5973, B2 => n6558
                           , ZN => n5359);
   U554 : NOR2_X1 port map( A1 => n6112, A2 => n5577, ZN => n6288);
   U555 : NAND2_X1 port map( A1 => n5185, A2 => DATA1(5), ZN => n5479);
   U556 : INV_X1 port map( A => n5479, ZN => n5349);
   U557 : AOI211_X1 port map( C1 => DATA1(1), C2 => n5785, A => n6288, B => 
                           n5349, ZN => n5350);
   U558 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(4), ZN => n5554);
   U559 : OAI211_X1 port map( C1 => n6113, C2 => n6648, A => n5350, B => n5554,
                           ZN => n5472);
   U560 : INV_X1 port map( A => n5351, ZN => n5353);
   U561 : INV_X1 port map( A => n5352, ZN => n5356);
   U562 : AOI222_X1 port map( A1 => n5472, A2 => n5672, B1 => n5353, B2 => 
                           n6549, C1 => n5356, C2 => n6547, ZN => n5899);
   U563 : INV_X1 port map( A => DATA1(1), ZN => n6327);
   U564 : NAND2_X1 port map( A1 => n5185, A2 => DATA1(4), ZN => n5519);
   U565 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(2), ZN => n6545);
   U566 : NAND2_X1 port map( A1 => n5519, A2 => n6545, ZN => n5354);
   U567 : AOI21_X1 port map( B1 => DATA1(0), B2 => n5785, A => n5354, ZN => 
                           n5355);
   U568 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(3), ZN => n6053);
   U569 : OAI211_X1 port map( C1 => n6113, C2 => n6327, A => n5355, B => n6053,
                           ZN => n5515);
   U570 : AOI222_X1 port map( A1 => n5515, A2 => n5672, B1 => n5356, B2 => 
                           n6549, C1 => n5472, C2 => n6547, ZN => n5976);
   U571 : OAI22_X1 port map( A1 => n5899, A2 => n6554, B1 => n5976, B2 => n6295
                           , ZN => n5358);
   U572 : NAND2_X1 port map( A1 => n5357, A2 => n6832, ZN => n6496);
   U573 : INV_X1 port map( A => n6496, ZN => n6527);
   U574 : OAI21_X1 port map( B1 => n5359, B2 => n5358, A => n6527, ZN => n5360)
                           ;
   U575 : OAI211_X1 port map( C1 => n6787, C2 => n6531, A => n5361, B => n5360,
                           ZN => n5362);
   U576 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_9_port, A => n5363
                           , B => n5362, ZN => n5367);
   U577 : AND2_X1 port map( A1 => n5774, A2 => DATA2_I_8_port, ZN => n5364);
   U578 : NOR2_X1 port map( A1 => n7166, A2 => n6457, ZN => n6504);
   U579 : NAND3_X1 port map( A1 => n5774, A2 => n5365, A3 => DATA2_I_8_port, ZN
                           => n6523);
   U580 : OAI211_X1 port map( C1 => n5365, C2 => n5364, A => n6504, B => n6523,
                           ZN => n5366);
   U581 : OAI211_X1 port map( C1 => n5368, C2 => n6830, A => n5367, B => n5366,
                           ZN => OUTALU(9));
   U582 : AOI22_X1 port map( A1 => n6236, A2 => n6515, B1 => n6518, B2 => n5478
                           , ZN => n5399);
   U583 : NOR2_X1 port map( A1 => DATA2(3), A2 => n5369, ZN => n5370);
   U584 : NAND2_X1 port map( A1 => n5371, A2 => n5370, ZN => n6083);
   U585 : INV_X1 port map( A => n6083, ZN => n6603);
   U586 : NOR2_X1 port map( A1 => n6112, A2 => n6662, ZN => n5638);
   U587 : INV_X1 port map( A => DATA1(12), ZN => n6693);
   U588 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(9), ZN => n5781);
   U589 : OAI211_X1 port map( C1 => n6055, C2 => n6693, A => n5781, B => n5372,
                           ZN => n5373);
   U590 : AOI211_X1 port map( C1 => DATA1(11), C2 => n6542, A => n5638, B => 
                           n5373, ZN => n5444);
   U591 : INV_X1 port map( A => n5374, ZN => n5375);
   U592 : OAI222_X1 port map( A1 => n6064, A2 => n5444, B1 => n6063, B2 => 
                           n5417, C1 => n6061, C2 => n5375, ZN => n5524);
   U593 : AOI22_X1 port map( A1 => n6232, A2 => n5376, B1 => n6197, B2 => n5524
                           , ZN => n5379);
   U594 : AOI22_X1 port map( A1 => n6565, A2 => n5418, B1 => n6067, B2 => n5377
                           , ZN => n5378);
   U595 : OAI211_X1 port map( C1 => n5380, C2 => n6558, A => n5379, B => n5378,
                           ZN => n5527);
   U596 : INV_X1 port map( A => n5527, ZN => n5492);
   U597 : OAI22_X1 port map( A1 => n5492, A2 => n5224, B1 => n5450, B2 => n6568
                           , ZN => n5383);
   U598 : OAI22_X1 port map( A1 => n6573, A2 => n5381, B1 => n5421, B2 => n6450
                           , ZN => n5382);
   U599 : AOI211_X1 port map( C1 => n6495, C2 => n5488, A => n5383, B => n5382,
                           ZN => n5451);
   U600 : OAI222_X1 port map( A1 => n5384, A2 => n5983, B1 => n5425, B2 => 
                           n6409, C1 => n5451, C2 => n6410, ZN => n5385);
   U601 : INV_X1 port map( A => n5385, ZN => n5532);
   U602 : INV_X1 port map( A => n5498, ZN => n5452);
   U603 : OAI22_X1 port map( A1 => n5532, A2 => n6588, B1 => n5452, B2 => n6592
                           , ZN => n5388);
   U604 : AOI22_X1 port map( A1 => n5455, A2 => n6470, B1 => n5426, B2 => n6595
                           , ZN => n5386);
   U605 : INV_X1 port map( A => n5386, ZN => n5387);
   U606 : AOI211_X1 port map( C1 => n5985, C2 => n6471, A => n5388, B => n5387,
                           ZN => n5539);
   U607 : INV_X1 port map( A => n5539, ZN => n5499);
   U608 : AOI22_X1 port map( A1 => n6603, A2 => n6517, B1 => n6509, B2 => n5499
                           , ZN => n5398);
   U609 : AOI21_X1 port map( B1 => DATA2_I_8_port, B2 => DATA1(8), A => n5389, 
                           ZN => n6004);
   U610 : INV_X1 port map( A => n5390, ZN => n6535);
   U611 : INV_X1 port map( A => n6004, ZN => n5396);
   U612 : INV_X1 port map( A => n5976, ZN => n5391);
   U613 : INV_X1 port map( A => n5899, ZN => n5979);
   U614 : AOI222_X1 port map( A1 => n5903, A2 => n6197, B1 => n5391, B2 => 
                           n6232, C1 => n5979, C2 => n6298, ZN => n5394);
   U615 : CLKBUF_X1 port map( A => n6183, Z => n6501);
   U616 : INV_X1 port map( A => DATA2(8), ZN => n6857);
   U617 : AOI22_X1 port map( A1 => DATA1(8), A2 => DATA2(8), B1 => n6857, B2 =>
                           n6715, ZN => n6813);
   U618 : AOI22_X1 port map( A1 => dataout_mul_8_port, A2 => n6501, B1 => n6631
                           , B2 => n6813, ZN => n5393);
   U619 : NAND3_X1 port map( A1 => DATA2(8), A2 => DATA1(8), A3 => n6528, ZN =>
                           n5392);
   U620 : OAI211_X1 port map( C1 => n5394, C2 => n6496, A => n5393, B => n5392,
                           ZN => n5395);
   U621 : AOI221_X1 port map( B1 => n6504, B2 => n6004, C1 => n6535, C2 => 
                           n5396, A => n5395, ZN => n5397);
   U622 : OAI221_X1 port map( B1 => n6830, B2 => n5399, C1 => n6830, C2 => 
                           n5398, A => n5397, ZN => OUTALU(8));
   U623 : OAI22_X1 port map( A1 => n6557, A2 => n5899, B1 => n5976, B2 => n6181
                           , ZN => n5400);
   U624 : AOI22_X1 port map( A1 => n6527, A2 => n5400, B1 => n6183, B2 => 
                           dataout_mul_7_port, ZN => n5440);
   U625 : INV_X1 port map( A => n5434, ZN => n5436);
   U626 : NOR2_X1 port map( A1 => n7166, A2 => cin, ZN => n6047);
   U627 : INV_X1 port map( A => n6047, ZN => n6637);
   U628 : INV_X1 port map( A => n6278, ZN => n6279);
   U629 : INV_X1 port map( A => n5401, ZN => n5402);
   U630 : AOI21_X1 port map( B1 => n6280, B2 => n6279, A => n5402, ZN => n6046)
                           ;
   U631 : OAI21_X1 port map( B1 => n6046, B2 => n6048, A => n5403, ZN => n5550)
                           ;
   U632 : AOI21_X1 port map( B1 => n5587, B2 => n5550, A => n5404, ZN => n5542)
                           ;
   U633 : OAI21_X1 port map( B1 => n5542, B2 => n5547, A => n5405, ZN => n5476)
                           ;
   U634 : INV_X1 port map( A => n5508, ZN => n5510);
   U635 : AOI21_X1 port map( B1 => n5476, B2 => n5510, A => n5406, ZN => n5464)
                           ;
   U636 : INV_X1 port map( A => n5468, ZN => n5465);
   U637 : OAI21_X1 port map( B1 => n5464, B2 => n5465, A => n5407, ZN => n5409)
                           ;
   U638 : NAND2_X1 port map( A1 => n6833, A2 => cin, ZN => n6042);
   U639 : NOR2_X1 port map( A1 => n5402, A2 => n6276, ZN => n6045);
   U640 : OAI21_X1 port map( B1 => n6045, B2 => n6048, A => n5403, ZN => n5549)
                           ;
   U641 : AOI21_X1 port map( B1 => n5587, B2 => n5549, A => n5404, ZN => n5541)
                           ;
   U642 : OAI21_X1 port map( B1 => n5541, B2 => n5547, A => n5405, ZN => n5475)
                           ;
   U643 : AOI21_X1 port map( B1 => n5475, B2 => n5510, A => n5406, ZN => n5463)
                           ;
   U644 : OAI21_X1 port map( B1 => n5463, B2 => n5465, A => n5407, ZN => n5408)
                           ;
   U645 : OAI22_X1 port map( A1 => n6637, A2 => n5409, B1 => n6042, B2 => n5408
                           , ZN => n5435);
   U646 : INV_X1 port map( A => n6042, ZN => n6632);
   U647 : AOI22_X1 port map( A1 => n5409, A2 => n6047, B1 => n5408, B2 => n6632
                           , ZN => n5410);
   U648 : INV_X1 port map( A => n5410, ZN => n5433);
   U649 : NOR2_X1 port map( A1 => n6864, A2 => n6863, ZN => n5411);
   U650 : OAI21_X1 port map( B1 => n5412, B2 => DATA2(2), A => n5411, ZN => 
                           n6610);
   U651 : CLKBUF_X1 port map( A => n6509, Z => n6516);
   U652 : INV_X1 port map( A => n5450, ZN => n5424);
   U653 : OAI22_X1 port map( A1 => n5492, A2 => n6570, B1 => n5413, B2 => n6568
                           , ZN => n5423);
   U654 : CLKBUF_X1 port map( A => n6197, Z => n6228);
   U655 : INV_X1 port map( A => n6000, ZN => n6491);
   U656 : NAND2_X1 port map( A1 => n6097, A2 => DATA1(9), ZN => n5771);
   U657 : OAI211_X1 port map( C1 => n6055, C2 => n6491, A => n5771, B => n5414,
                           ZN => n5415);
   U658 : AOI211_X1 port map( C1 => DATA1(10), C2 => n6542, A => n5416, B => 
                           n5415, ZN => n5484);
   U659 : OAI222_X1 port map( A1 => n6064, A2 => n5484, B1 => n6063, B2 => 
                           n5444, C1 => n6061, C2 => n5417, ZN => n5561);
   U660 : AOI22_X1 port map( A1 => n6298, A2 => n5524, B1 => n6228, B2 => n5561
                           , ZN => n5420);
   U661 : AOI22_X1 port map( A1 => n6232, A2 => n5485, B1 => n6067, B2 => n5418
                           , ZN => n5419);
   U662 : OAI211_X1 port map( C1 => n5447, C2 => n6295, A => n5420, B => n5419,
                           ZN => n5489);
   U663 : INV_X1 port map( A => n5489, ZN => n5564);
   U664 : OAI22_X1 port map( A1 => n5564, A2 => n5224, B1 => n6573, B2 => n5421
                           , ZN => n5422);
   U665 : AOI211_X1 port map( C1 => n6577, C2 => n5424, A => n5423, B => n5422,
                           ZN => n5493);
   U666 : OAI222_X1 port map( A1 => n6409, A2 => n5451, B1 => n6410, B2 => 
                           n5493, C1 => n5425, C2 => n5894, ZN => n5567);
   U667 : AOI22_X1 port map( A1 => n6595, A2 => n5455, B1 => n5985, B2 => n5426
                           , ZN => n5427);
   U668 : OAI21_X1 port map( B1 => n5452, B2 => n6586, A => n5427, ZN => n5428)
                           ;
   U669 : AOI21_X1 port map( B1 => n6472, B2 => n5567, A => n5428, ZN => n5571)
                           ;
   U670 : OAI21_X1 port map( B1 => n5532, B2 => n6592, A => n5571, ZN => n5535)
                           ;
   U671 : AOI22_X1 port map( A1 => n6518, A2 => n5499, B1 => n6516, B2 => n5535
                           , ZN => n5430);
   U672 : AOI22_X1 port map( A1 => n6605, A2 => n6517, B1 => n6236, B2 => n5478
                           , ZN => n5429);
   U673 : OAI211_X1 port map( C1 => n5431, C2 => n6083, A => n5430, B => n5429,
                           ZN => n5503);
   U674 : INV_X1 port map( A => n6830, ZN => n6510);
   U675 : AND3_X1 port map( A1 => n6610, A2 => n5503, A3 => n6510, ZN => n5432)
                           ;
   U676 : AOI221_X1 port map( B1 => n5436, B2 => n5435, C1 => n5434, C2 => 
                           n5433, A => n5432, ZN => n5439);
   U677 : INV_X1 port map( A => n6389, ZN => n6633);
   U678 : OAI211_X1 port map( C1 => n6493, C2 => n6633, A => DATA1(7), B => 
                           DATA2(7), ZN => n5438);
   U679 : NOR2_X1 port map( A1 => DATA2(7), A2 => n5782, ZN => n6712);
   U680 : INV_X1 port map( A => DATA2(7), ZN => n6860);
   U681 : NOR2_X1 port map( A1 => DATA1(7), A2 => n6860, ZN => n6694);
   U682 : OAI21_X1 port map( B1 => n6712, B2 => n6694, A => n6631, ZN => n5437)
                           ;
   U683 : NAND4_X1 port map( A1 => n5440, A2 => n5439, A3 => n5438, A4 => n5437
                           , ZN => OUTALU(7));
   U684 : AOI211_X1 port map( C1 => n6865, C2 => n6866, A => n6864, B => n6863,
                           ZN => n5923);
   U685 : CLKBUF_X1 port map( A => n6610, Z => n6321);
   U686 : NOR2_X1 port map( A1 => n5923, A2 => n6321, ZN => n6089);
   U687 : INV_X1 port map( A => n6315, ZN => n6600);
   U688 : NAND2_X1 port map( A1 => n6097, A2 => n5774, ZN => n5780);
   U689 : OAI211_X1 port map( C1 => n5691, C2 => n6662, A => n5780, B => n5441,
                           ZN => n5442);
   U690 : AOI211_X1 port map( C1 => DATA1(9), C2 => n6542, A => n5443, B => 
                           n5442, ZN => n5523);
   U691 : OAI222_X1 port map( A1 => n6064, A2 => n5523, B1 => n6063, B2 => 
                           n5484, C1 => n6061, C2 => n5444, ZN => n6066);
   U692 : AOI22_X1 port map( A1 => n6230, A2 => n5561, B1 => n6228, B2 => n6066
                           , ZN => n5446);
   U693 : AOI22_X1 port map( A1 => n6565, A2 => n5485, B1 => n6232, B2 => n5524
                           , ZN => n5445);
   U694 : OAI211_X1 port map( C1 => n6561, C2 => n5447, A => n5446, B => n5445,
                           ZN => n6071);
   U695 : AOI22_X1 port map( A1 => n6495, A2 => n5489, B1 => n6526, B2 => n6071
                           , ZN => n5449);
   U696 : AOI22_X1 port map( A1 => n6468, A2 => n5527, B1 => n6577, B2 => n5488
                           , ZN => n5448);
   U697 : OAI211_X1 port map( C1 => n5450, C2 => n6573, A => n5449, B => n5448,
                           ZN => n5530);
   U698 : INV_X1 port map( A => n5530, ZN => n5495);
   U699 : OAI222_X1 port map( A1 => n6410, A2 => n5495, B1 => n6409, B2 => 
                           n5493, C1 => n5451, C2 => n5894, ZN => n5568);
   U700 : INV_X1 port map( A => n5568, ZN => n6077);
   U701 : OAI22_X1 port map( A1 => n6077, A2 => n6588, B1 => n5532, B2 => n6586
                           , ZN => n5454);
   U702 : INV_X1 port map( A => n5567, ZN => n5531);
   U703 : OAI22_X1 port map( A1 => n5531, A2 => n6592, B1 => n5452, B2 => n6310
                           , ZN => n5453);
   U704 : AOI211_X1 port map( C1 => n5985, C2 => n5455, A => n5454, B => n5453,
                           ZN => n6082);
   U705 : INV_X1 port map( A => n6082, ZN => n5536);
   U706 : AOI22_X1 port map( A1 => n6605, A2 => n5456, B1 => n6516, B2 => n5536
                           , ZN => n5458);
   U707 : AOI22_X1 port map( A1 => n6603, A2 => n5478, B1 => n6518, B2 => n5535
                           , ZN => n5457);
   U708 : OAI211_X1 port map( C1 => n5539, C2 => n6600, A => n5458, B => n5457,
                           ZN => n5540);
   U709 : AOI22_X1 port map( A1 => n6089, A2 => n5503, B1 => n6321, B2 => n5540
                           , ZN => n5471);
   U710 : NOR3_X1 port map( A1 => n6292, A2 => n5976, A3 => n6496, ZN => n5461)
                           ;
   U711 : INV_X1 port map( A => DATA2(6), ZN => n6861);
   U712 : AOI22_X1 port map( A1 => DATA1(6), A2 => n6861, B1 => DATA2(6), B2 =>
                           n6695, ZN => n6711);
   U713 : AOI21_X1 port map( B1 => n6633, B2 => DATA1(6), A => n6493, ZN => 
                           n5459);
   U714 : OAI22_X1 port map( A1 => n6711, A2 => n6531, B1 => n5459, B2 => n6861
                           , ZN => n5460);
   U715 : AOI211_X1 port map( C1 => dataout_mul_6_port, C2 => n6501, A => n5461
                           , B => n5460, ZN => n5470);
   U716 : AOI22_X1 port map( A1 => n6047, A2 => n5464, B1 => n6632, B2 => n5463
                           , ZN => n5462);
   U717 : INV_X1 port map( A => n5462, ZN => n5467);
   U718 : OAI22_X1 port map( A1 => n5464, A2 => n6637, B1 => n5463, B2 => n6042
                           , ZN => n5466);
   U719 : AOI22_X1 port map( A1 => n5468, A2 => n5467, B1 => n5466, B2 => n5465
                           , ZN => n5469);
   U720 : OAI211_X1 port map( C1 => n5471, C2 => n6830, A => n5470, B => n5469,
                           ZN => OUTALU(6));
   U721 : AOI21_X1 port map( B1 => n6633, B2 => DATA1(5), A => n6493, ZN => 
                           n5513);
   U722 : NAND2_X1 port map( A1 => n6059, A2 => n6862, ZN => n6710);
   U723 : OR2_X1 port map( A1 => n6862, A2 => n6059, ZN => n6706);
   U724 : AND2_X1 port map( A1 => n6710, A2 => n6706, ZN => n6789);
   U725 : AOI22_X1 port map( A1 => n6152, A2 => n5472, B1 => n6547, B2 => n5515
                           , ZN => n5473);
   U726 : OAI22_X1 port map( A1 => n6789, A2 => n6531, B1 => n5473, B2 => n6496
                           , ZN => n5474);
   U727 : AOI21_X1 port map( B1 => n6641, B2 => dataout_mul_5_port, A => n5474,
                           ZN => n5512);
   U728 : OAI22_X1 port map( A1 => n6637, A2 => n5476, B1 => n6042, B2 => n5475
                           , ZN => n5509);
   U729 : AOI22_X1 port map( A1 => n5476, A2 => n6047, B1 => n5475, B2 => n6632
                           , ZN => n5477);
   U730 : INV_X1 port map( A => n5477, ZN => n5507);
   U731 : CLKBUF_X1 port map( A => n5923, Z => n6615);
   U732 : INV_X1 port map( A => n5478, ZN => n5502);
   U733 : INV_X1 port map( A => n6066, ZN => n5558);
   U734 : OAI211_X1 port map( C1 => n6055, C2 => n5481, A => n5480, B => n5479,
                           ZN => n5482);
   U735 : AOI211_X1 port map( C1 => n5774, C2 => n6542, A => n5483, B => n5482,
                           ZN => n5557);
   U736 : OAI222_X1 port map( A1 => n6064, A2 => n5557, B1 => n6063, B2 => 
                           n5523, C1 => n6061, C2 => n5484, ZN => n6068);
   U737 : AOI22_X1 port map( A1 => n6232, A2 => n5561, B1 => n6228, B2 => n6068
                           , ZN => n5487);
   U738 : AOI22_X1 port map( A1 => n6565, A2 => n5524, B1 => n6067, B2 => n5485
                           , ZN => n5486);
   U739 : OAI211_X1 port map( C1 => n5558, C2 => n6181, A => n5487, B => n5486,
                           ZN => n6301);
   U740 : AOI22_X1 port map( A1 => n6495, A2 => n6071, B1 => n6526, B2 => n6301
                           , ZN => n5491);
   U741 : CLKBUF_X1 port map( A => n6072, Z => n6302);
   U742 : AOI22_X1 port map( A1 => n6468, A2 => n5489, B1 => n6302, B2 => n5488
                           , ZN => n5490);
   U743 : OAI211_X1 port map( C1 => n5492, C2 => n6450, A => n5491, B => n5490,
                           ZN => n5565);
   U744 : INV_X1 port map( A => n5565, ZN => n5494);
   U745 : OAI222_X1 port map( A1 => n6409, A2 => n5495, B1 => n6410, B2 => 
                           n5494, C1 => n5493, C2 => n5983, ZN => n5566);
   U746 : INV_X1 port map( A => n5566, ZN => n6309);
   U747 : OAI22_X1 port map( A1 => n5531, A2 => n6586, B1 => n6309, B2 => n6588
                           , ZN => n5497);
   U748 : OAI22_X1 port map( A1 => n6077, A2 => n6592, B1 => n5532, B2 => n6310
                           , ZN => n5496);
   U749 : AOI211_X1 port map( C1 => n5985, C2 => n5498, A => n5497, B => n5496,
                           ZN => n6084);
   U750 : INV_X1 port map( A => n6084, ZN => n6317);
   U751 : AOI22_X1 port map( A1 => n6236, A2 => n5535, B1 => n6516, B2 => n6317
                           , ZN => n5501);
   U752 : AOI22_X1 port map( A1 => n6603, A2 => n5499, B1 => n6518, B2 => n5536
                           , ZN => n5500);
   U753 : OAI211_X1 port map( C1 => n5502, C2 => n6081, A => n5501, B => n5500,
                           ZN => n5575);
   U754 : AOI222_X1 port map( A1 => n6615, A2 => n5503, B1 => n5540, B2 => 
                           n6089, C1 => n5575, C2 => n6321, ZN => n6322);
   U755 : AOI211_X1 port map( C1 => n6865, C2 => n5504, A => n6864, B => n6863,
                           ZN => n5505);
   U756 : CLKBUF_X1 port map( A => n5505, Z => n6616);
   U757 : NOR3_X1 port map( A1 => n6322, A2 => n6830, A3 => n6616, ZN => n5506)
                           ;
   U758 : AOI221_X1 port map( B1 => n5510, B2 => n5509, C1 => n5508, C2 => 
                           n5507, A => n5506, ZN => n5511);
   U759 : OAI211_X1 port map( C1 => n5513, C2 => n6862, A => n5512, B => n5511,
                           ZN => OUTALU(5));
   U760 : AOI22_X1 port map( A1 => n6047, A2 => n5542, B1 => n6632, B2 => n5541
                           , ZN => n5548);
   U761 : AOI211_X1 port map( C1 => n6388, C2 => n6389, A => n6863, B => n5514,
                           ZN => n5518);
   U762 : NAND2_X1 port map( A1 => DATA2(4), A2 => n5514, ZN => n6707);
   U763 : NAND2_X1 port map( A1 => n6863, A2 => DATA1(4), ZN => n6704);
   U764 : NAND3_X1 port map( A1 => n6527, A2 => n6152, A3 => n5515, ZN => n5516
                           );
   U765 : OAI221_X1 port map( B1 => n6492, B2 => n6707, C1 => n6531, C2 => 
                           n6704, A => n5516, ZN => n5517);
   U766 : AOI211_X1 port map( C1 => dataout_mul_4_port, C2 => n6501, A => n5518
                           , B => n5517, ZN => n5546);
   U767 : CLKBUF_X1 port map( A => n6089, Z => n6612);
   U768 : OAI211_X1 port map( C1 => n6055, C2 => n6715, A => n5520, B => n5519,
                           ZN => n5521);
   U769 : AOI211_X1 port map( C1 => DATA1(7), C2 => n6542, A => n5522, B => 
                           n5521, ZN => n6060);
   U770 : OAI222_X1 port map( A1 => n6064, A2 => n6060, B1 => n6063, B2 => 
                           n5557, C1 => n6061, C2 => n5523, ZN => n6065);
   U771 : AOI22_X1 port map( A1 => n6565, A2 => n5561, B1 => n6228, B2 => n6065
                           , ZN => n5526);
   U772 : AOI22_X1 port map( A1 => n6298, A2 => n6068, B1 => n6067, B2 => n5524
                           , ZN => n5525);
   U773 : OAI211_X1 port map( C1 => n5558, C2 => n6554, A => n5526, B => n5525,
                           ZN => n6303);
   U774 : AOI22_X1 port map( A1 => n6468, A2 => n6071, B1 => n6526, B2 => n6303
                           , ZN => n5529);
   U775 : AOI22_X1 port map( A1 => n6073, A2 => n6301, B1 => n6302, B2 => n5527
                           , ZN => n5528);
   U776 : OAI211_X1 port map( C1 => n5564, C2 => n6450, A => n5529, B => n5528,
                           ZN => n6076);
   U777 : INV_X1 port map( A => n6409, ZN => n6584);
   U778 : AOI222_X1 port map( A1 => n5530, A2 => n6579, B1 => n6076, B2 => 
                           n6582, C1 => n5565, C2 => n6584, ZN => n6589);
   U779 : OAI22_X1 port map( A1 => n6589, A2 => n6307, B1 => n6077, B2 => n6586
                           , ZN => n5534);
   U780 : OAI22_X1 port map( A1 => n6590, A2 => n5532, B1 => n5531, B2 => n6310
                           , ZN => n5533);
   U781 : AOI211_X1 port map( C1 => n6475, C2 => n5566, A => n5534, B => n5533,
                           ZN => n6080);
   U782 : INV_X1 port map( A => n6080, ZN => n6604);
   U783 : AOI22_X1 port map( A1 => n6603, A2 => n5535, B1 => n6516, B2 => n6604
                           , ZN => n5538);
   U784 : AOI22_X1 port map( A1 => n6236, A2 => n5536, B1 => n6518, B2 => n6317
                           , ZN => n5537);
   U785 : OAI211_X1 port map( C1 => n5539, C2 => n6081, A => n5538, B => n5537,
                           ZN => n6088);
   U786 : AOI222_X1 port map( A1 => n5923, A2 => n5540, B1 => n5575, B2 => 
                           n6612, C1 => n6088, C2 => n6321, ZN => n6623);
   U787 : INV_X1 port map( A => n6616, ZN => n5998);
   U788 : NOR2_X1 port map( A1 => n5927, A2 => n5998, ZN => n6627);
   U789 : INV_X1 port map( A => n6627, ZN => n6139);
   U790 : OAI22_X1 port map( A1 => n6623, A2 => n6616, B1 => n6322, B2 => n6139
                           , ZN => n5544);
   U791 : OAI22_X1 port map( A1 => n5542, A2 => n6637, B1 => n5541, B2 => n6042
                           , ZN => n5543);
   U792 : AOI22_X1 port map( A1 => n6510, A2 => n5544, B1 => n5547, B2 => n5543
                           , ZN => n5545);
   U793 : OAI211_X1 port map( C1 => n5548, C2 => n5547, A => n5546, B => n5545,
                           ZN => OUTALU(4));
   U794 : AOI22_X1 port map( A1 => n6047, A2 => n5550, B1 => n6632, B2 => n5549
                           , ZN => n5586);
   U795 : INV_X1 port map( A => n5587, ZN => n5585);
   U796 : OAI22_X1 port map( A1 => n6637, A2 => n5550, B1 => n6042, B2 => n5549
                           , ZN => n5551);
   U797 : INV_X1 port map( A => n5551, ZN => n5584);
   U798 : NAND2_X1 port map( A1 => n5927, A2 => n5552, ZN => n6618);
   U799 : AOI22_X1 port map( A1 => DATA1(3), A2 => n5825, B1 => DATA1(7), B2 =>
                           n5601, ZN => n5556);
   U800 : NAND4_X1 port map( A1 => n5556, A2 => n5555, A3 => n5554, A4 => n5553
                           , ZN => n6291);
   U801 : INV_X1 port map( A => n6291, ZN => n6062);
   U802 : OAI222_X1 port map( A1 => n5557, A2 => n6061, B1 => n6062, B2 => 
                           n6064, C1 => n6060, C2 => n6063, ZN => n6564);
   U803 : INV_X1 port map( A => n6564, ZN => n6293);
   U804 : OAI22_X1 port map( A1 => n6292, A2 => n6293, B1 => n5558, B2 => n6295
                           , ZN => n5560);
   U805 : INV_X1 port map( A => n6068, ZN => n6294);
   U806 : INV_X1 port map( A => n6065, ZN => n6560);
   U807 : OAI22_X1 port map( A1 => n6294, A2 => n6554, B1 => n6560, B2 => n6181
                           , ZN => n5559);
   U808 : AOI211_X1 port map( C1 => n6067, C2 => n5561, A => n5560, B => n5559,
                           ZN => n6299);
   U809 : INV_X1 port map( A => n6299, ZN => n6576);
   U810 : AOI22_X1 port map( A1 => n6071, A2 => n6577, B1 => n6576, B2 => n6526
                           , ZN => n5563);
   U811 : AOI22_X1 port map( A1 => n6301, A2 => n6468, B1 => n6303, B2 => n6495
                           , ZN => n5562);
   U812 : OAI211_X1 port map( C1 => n6573, C2 => n5564, A => n5563, B => n5562,
                           ZN => n6306);
   U813 : AOI222_X1 port map( A1 => n6584, A2 => n6076, B1 => n6582, B2 => 
                           n6306, C1 => n5565, C2 => n6579, ZN => n6308);
   U814 : INV_X1 port map( A => n6308, ZN => n6596);
   U815 : AOI22_X1 port map( A1 => n6472, A2 => n6596, B1 => n6470, B2 => n5566
                           , ZN => n5570);
   U816 : AOI22_X1 port map( A1 => n6595, A2 => n5568, B1 => n5985, B2 => n5567
                           , ZN => n5569);
   U817 : OAI211_X1 port map( C1 => n6589, C2 => n6592, A => n5570, B => n5569,
                           ZN => n6602);
   U818 : OAI22_X1 port map( A1 => n6080, A2 => n6608, B1 => n5571, B2 => n6081
                           , ZN => n5573);
   U819 : OAI22_X1 port map( A1 => n6084, A2 => n6600, B1 => n6082, B2 => n6083
                           , ZN => n5572);
   U820 : AOI211_X1 port map( C1 => n6509, C2 => n6602, A => n5573, B => n5572,
                           ZN => n5574);
   U821 : INV_X1 port map( A => n5574, ZN => n6320);
   U822 : AOI222_X1 port map( A1 => n5923, A2 => n5575, B1 => n6088, B2 => 
                           n6089, C1 => n6321, C2 => n6320, ZN => n6621);
   U823 : OAI222_X1 port map( A1 => n6139, A2 => n6623, B1 => n6618, B2 => 
                           n6322, C1 => n6616, C2 => n6621, ZN => n5582);
   U824 : INV_X1 port map( A => n6528, ZN => n6149);
   U825 : NOR3_X1 port map( A1 => n6149, A2 => n5577, A3 => n6864, ZN => n5581)
                           ;
   U826 : NOR2_X1 port map( A1 => n6864, A2 => DATA1(3), ZN => n6701);
   U827 : INV_X1 port map( A => n6701, ZN => n6652);
   U828 : NAND2_X1 port map( A1 => n6864, A2 => DATA1(3), ZN => n6705);
   U829 : AOI22_X1 port map( A1 => n6542, A2 => DATA1(0), B1 => n6097, B2 => 
                           DATA1(1), ZN => n5576);
   U830 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(2), ZN => n6286);
   U831 : OAI211_X1 port map( C1 => n5577, C2 => n6326, A => n5576, B => n6286,
                           ZN => n5578);
   U832 : AOI22_X1 port map( A1 => n6527, A2 => n5578, B1 => n6183, B2 => 
                           dataout_mul_3_port, ZN => n5579);
   U833 : OAI221_X1 port map( B1 => n6531, B2 => n6652, C1 => n6531, C2 => 
                           n6705, A => n5579, ZN => n5580);
   U834 : AOI211_X1 port map( C1 => n6510, C2 => n5582, A => n5581, B => n5580,
                           ZN => n5583);
   U835 : OAI221_X1 port map( B1 => n5587, B2 => n5586, C1 => n5585, C2 => 
                           n5584, A => n5583, ZN => OUTALU(3));
   U836 : NAND2_X1 port map( A1 => n7169, A2 => n5785, ZN => n5588);
   U837 : NAND4_X1 port map( A1 => n5591, A2 => n5590, A3 => n5589, A4 => n5588
                           , ZN => n5592);
   U838 : AOI21_X1 port map( B1 => DATA1(18), B2 => n5825, A => n5592, ZN => 
                           n5631);
   U839 : NOR2_X1 port map( A1 => n5691, A2 => n6447, ZN => n5596);
   U840 : OAI211_X1 port map( C1 => n6375, C2 => n6326, A => n5594, B => n5593,
                           ZN => n5595);
   U841 : AOI211_X1 port map( C1 => DATA1(14), C2 => n6542, A => n5596, B => 
                           n5595, ZN => n5620);
   U842 : OAI211_X1 port map( C1 => n6055, C2 => n6693, A => n5598, B => n5597,
                           ZN => n5599);
   U843 : AOI211_X1 port map( C1 => DATA1(16), C2 => n5825, A => n5600, B => 
                           n5599, ZN => n5623);
   U844 : OAI222_X1 port map( A1 => n6064, A2 => n5631, B1 => n6063, B2 => 
                           n5620, C1 => n6061, C2 => n5623, ZN => n5660);
   U845 : AOI22_X1 port map( A1 => n6058, A2 => DATA1(10), B1 => n5825, B2 => 
                           DATA1(13), ZN => n5605);
   U846 : NAND2_X1 port map( A1 => DATA1(9), A2 => n5601, ZN => n5602);
   U847 : NAND4_X1 port map( A1 => n5605, A2 => n5604, A3 => n5603, A4 => n5602
                           , ZN => n5634);
   U848 : AOI22_X1 port map( A1 => n6058, A2 => DATA1(12), B1 => n5185, B2 => 
                           DATA1(15), ZN => n5609);
   U849 : NAND2_X1 port map( A1 => n6000, A2 => n5785, ZN => n5606);
   U850 : NAND4_X1 port map( A1 => n5609, A2 => n5608, A3 => n5607, A4 => n5606
                           , ZN => n5614);
   U851 : AOI22_X1 port map( A1 => n6542, A2 => n6000, B1 => n5825, B2 => 
                           DATA1(14), ZN => n5613);
   U852 : NAND2_X1 port map( A1 => n7167, A2 => n5785, ZN => n5610);
   U853 : NAND4_X1 port map( A1 => n5613, A2 => n5612, A3 => n5611, A4 => n5610
                           , ZN => n5621);
   U854 : AOI222_X1 port map( A1 => n5634, A2 => n6551, B1 => n5614, B2 => 
                           n6549, C1 => n5621, C2 => n6547, ZN => n5807);
   U855 : INV_X1 port map( A => n5614, ZN => n5622);
   U856 : OAI222_X1 port map( A1 => n5622, A2 => n6061, B1 => n5620, B2 => 
                           n6064, C1 => n5623, C2 => n6063, ZN => n5647);
   U857 : INV_X1 port map( A => n5647, ZN => n5776);
   U858 : OAI22_X1 port map( A1 => n6561, A2 => n5807, B1 => n5776, B2 => n6554
                           , ZN => n5626);
   U859 : AOI21_X1 port map( B1 => n5185, B2 => DATA1(19), A => n5615, ZN => 
                           n5619);
   U860 : NAND2_X1 port map( A1 => DATA1(15), A2 => n5785, ZN => n5617);
   U861 : AND4_X1 port map( A1 => n5619, A2 => n5618, A3 => n5617, A4 => n5616,
                           ZN => n5646);
   U862 : OAI222_X1 port map( A1 => n5620, A2 => n6061, B1 => n5646, B2 => 
                           n6064, C1 => n5631, C2 => n6063, ZN => n5673);
   U863 : INV_X1 port map( A => n5621, ZN => n5639);
   U864 : OAI222_X1 port map( A1 => n5639, A2 => n6061, B1 => n5623, B2 => 
                           n6064, C1 => n5622, C2 => n6063, ZN => n5787);
   U865 : AOI22_X1 port map( A1 => n6197, A2 => n5673, B1 => n5787, B2 => n6565
                           , ZN => n5624);
   U866 : INV_X1 port map( A => n5624, ZN => n5625);
   U867 : AOI211_X1 port map( C1 => n6298, C2 => n5660, A => n5626, B => n5625,
                           ZN => n5811);
   U868 : INV_X1 port map( A => DATA1(16), ZN => n6735);
   U869 : NOR2_X1 port map( A1 => n6055, A2 => n6735, ZN => n5630);
   U870 : OAI211_X1 port map( C1 => n6326, C2 => n6747, A => n5628, B => n5627,
                           ZN => n5629);
   U871 : AOI211_X1 port map( C1 => DATA1(17), C2 => n6542, A => n5630, B => 
                           n5629, ZN => n5651);
   U872 : OAI222_X1 port map( A1 => n6064, A2 => n5651, B1 => n6063, B2 => 
                           n5646, C1 => n6061, C2 => n5631, ZN => n5688);
   U873 : AOI22_X1 port map( A1 => n6067, A2 => n5787, B1 => n6228, B2 => n5688
                           , ZN => n5633);
   U874 : AOI22_X1 port map( A1 => n6230, A2 => n5673, B1 => n6232, B2 => n5660
                           , ZN => n5632);
   U875 : OAI211_X1 port map( C1 => n5776, C2 => n6295, A => n5633, B => n5632,
                           ZN => n5794);
   U876 : INV_X1 port map( A => n5634, ZN => n5775);
   U877 : NAND2_X1 port map( A1 => n5185, A2 => n7168, ZN => n5635);
   U878 : OAI211_X1 port map( C1 => n6055, C2 => n6715, A => n5636, B => n5635,
                           ZN => n5637);
   U879 : AOI211_X1 port map( C1 => DATA1(9), C2 => n6058, A => n5638, B => 
                           n5637, ZN => n5786);
   U880 : OAI222_X1 port map( A1 => n6064, A2 => n5639, B1 => n6063, B2 => 
                           n5775, C1 => n6061, C2 => n5786, ZN => n5853);
   U881 : AOI22_X1 port map( A1 => n6232, A2 => n5787, B1 => n6067, B2 => n5853
                           , ZN => n5641);
   U882 : AOI22_X1 port map( A1 => n6298, A2 => n5647, B1 => n6228, B2 => n5660
                           , ZN => n5640);
   U883 : OAI211_X1 port map( C1 => n5807, C2 => n6295, A => n5641, B => n5640,
                           ZN => n5858);
   U884 : AOI22_X1 port map( A1 => n6468, A2 => n5794, B1 => n6302, B2 => n5858
                           , ZN => n5664);
   U885 : INV_X1 port map( A => n5688, ZN => n5650);
   U886 : NOR2_X1 port map( A1 => n5691, A2 => n6375, ZN => n5645);
   U887 : OAI211_X1 port map( C1 => n6248, C2 => n6326, A => n5643, B => n5642,
                           ZN => n5644);
   U888 : AOI211_X1 port map( C1 => DATA1(18), C2 => n6542, A => n5645, B => 
                           n5644, ZN => n5658);
   U889 : OAI222_X1 port map( A1 => n6064, A2 => n5658, B1 => n6063, B2 => 
                           n5651, C1 => n6061, C2 => n5646, ZN => n5699);
   U890 : AOI22_X1 port map( A1 => n6067, A2 => n5647, B1 => n6228, B2 => n5699
                           , ZN => n5649);
   U891 : AOI22_X1 port map( A1 => n6565, A2 => n5660, B1 => n6232, B2 => n5673
                           , ZN => n5648);
   U892 : OAI211_X1 port map( C1 => n5650, C2 => n6558, A => n5649, B => n5648,
                           ZN => n5793);
   U893 : INV_X1 port map( A => n5651, ZN => n5659);
   U894 : INV_X1 port map( A => n5652, ZN => n5653);
   U895 : AOI211_X1 port map( C1 => n5185, C2 => DATA1(22), A => n5654, B => 
                           n5653, ZN => n5657);
   U896 : NAND3_X1 port map( A1 => n5657, A2 => n5656, A3 => n5655, ZN => n5684
                           );
   U897 : INV_X1 port map( A => n5658, ZN => n5671);
   U898 : AOI222_X1 port map( A1 => n5659, A2 => n6551, B1 => n5684, B2 => 
                           n6549, C1 => n5671, C2 => n6547, ZN => n5719);
   U899 : AOI22_X1 port map( A1 => n6230, A2 => n5699, B1 => n6067, B2 => n5660
                           , ZN => n5662);
   U900 : AOI22_X1 port map( A1 => n6565, A2 => n5673, B1 => n6232, B2 => n5688
                           , ZN => n5661);
   U901 : OAI211_X1 port map( C1 => n6292, C2 => n5719, A => n5662, B => n5661,
                           ZN => n5744);
   U902 : AOI22_X1 port map( A1 => n6073, A2 => n5793, B1 => n6526, B2 => n5744
                           , ZN => n5663);
   U903 : OAI211_X1 port map( C1 => n5811, C2 => n6450, A => n5664, B => n5663,
                           ZN => n5799);
   U904 : INV_X1 port map( A => n5794, ZN => n5678);
   U905 : INV_X1 port map( A => n5665, ZN => n5668);
   U906 : AND4_X1 port map( A1 => n5669, A2 => n5668, A3 => n5667, A4 => n5666,
                           ZN => n5670);
   U907 : OAI21_X1 port map( B1 => n6326, B2 => n6198, A => n5670, ZN => n5697)
                           ;
   U908 : AOI222_X1 port map( A1 => n6549, A2 => n5697, B1 => n6547, B2 => 
                           n5684, C1 => n5672, C2 => n5671, ZN => n5718);
   U909 : INV_X1 port map( A => n5718, ZN => n5698);
   U910 : AOI22_X1 port map( A1 => n6067, A2 => n5673, B1 => n6228, B2 => n5698
                           , ZN => n5675);
   U911 : AOI22_X1 port map( A1 => n6565, A2 => n5688, B1 => n6232, B2 => n5699
                           , ZN => n5674);
   U912 : OAI211_X1 port map( C1 => n5719, C2 => n6558, A => n5675, B => n5674,
                           ZN => n5740);
   U913 : INV_X1 port map( A => n5811, ZN => n5792);
   U914 : AOI22_X1 port map( A1 => n6526, A2 => n5740, B1 => n6072, B2 => n5792
                           , ZN => n5677);
   U915 : AOI22_X1 port map( A1 => n6468, A2 => n5793, B1 => n6073, B2 => n5744
                           , ZN => n5676);
   U916 : OAI211_X1 port map( C1 => n5678, C2 => n6450, A => n5677, B => n5676,
                           ZN => n5798);
   U917 : AOI21_X1 port map( B1 => DATA1(20), B2 => n5785, A => n5679, ZN => 
                           n5683);
   U918 : NAND4_X1 port map( A1 => n5683, A2 => n5682, A3 => n5681, A4 => n5680
                           , ZN => n5713);
   U919 : AOI222_X1 port map( A1 => n5684, A2 => n6551, B1 => n5713, B2 => 
                           n6549, C1 => n5697, C2 => n6547, ZN => n5714);
   U920 : OAI22_X1 port map( A1 => n6557, A2 => n5714, B1 => n5718, B2 => n6558
                           , ZN => n5687);
   U921 : INV_X1 port map( A => n5699, ZN => n5685);
   U922 : OAI22_X1 port map( A1 => n5685, A2 => n6295, B1 => n5719, B2 => n6554
                           , ZN => n5686);
   U923 : AOI211_X1 port map( C1 => n6067, C2 => n5688, A => n5687, B => n5686,
                           ZN => n5739);
   U924 : INV_X1 port map( A => n5740, ZN => n5736);
   U925 : AOI22_X1 port map( A1 => n6468, A2 => n5744, B1 => n6577, B2 => n5793
                           , ZN => n5689);
   U926 : OAI21_X1 port map( B1 => n5736, B2 => n6570, A => n5689, ZN => n5690)
                           ;
   U927 : AOI21_X1 port map( B1 => n6302, B2 => n5794, A => n5690, ZN => n5747)
                           ;
   U928 : OAI21_X1 port map( B1 => n5739, B2 => n6566, A => n5747, ZN => n5746)
                           ;
   U929 : AOI222_X1 port map( A1 => n5799, A2 => n6579, B1 => n5798, B2 => 
                           n6584, C1 => n5746, C2 => n6582, ZN => n5816);
   U930 : NOR2_X1 port map( A1 => n5691, A2 => n6248, ZN => n5695);
   U931 : INV_X1 port map( A => DATA1(25), ZN => n6166);
   U932 : OAI211_X1 port map( C1 => n6326, C2 => n6166, A => n5693, B => n5692,
                           ZN => n5694);
   U933 : AOI211_X1 port map( C1 => DATA1(22), C2 => n6058, A => n5695, B => 
                           n5694, ZN => n5696);
   U934 : INV_X1 port map( A => n5696, ZN => n5712);
   U935 : AOI222_X1 port map( A1 => n6549, A2 => n5712, B1 => n6547, B2 => 
                           n5713, C1 => n6551, C2 => n5697, ZN => n5759);
   U936 : INV_X1 port map( A => n5759, ZN => n5717);
   U937 : AOI22_X1 port map( A1 => n6232, A2 => n5698, B1 => n6228, B2 => n5717
                           , ZN => n5701);
   U938 : INV_X1 port map( A => n5714, ZN => n5732);
   U939 : AOI22_X1 port map( A1 => n6298, A2 => n5732, B1 => n6067, B2 => n5699
                           , ZN => n5700);
   U940 : OAI211_X1 port map( C1 => n5719, C2 => n6295, A => n5701, B => n5700,
                           ZN => n5724);
   U941 : AND3_X1 port map( A1 => n5704, A2 => n5703, A3 => n5702, ZN => n5706)
                           ;
   U942 : OAI211_X1 port map( C1 => n6113, C2 => n6680, A => n5706, B => n5705,
                           ZN => n5758);
   U943 : AOI211_X1 port map( C1 => n6753, C2 => n5785, A => n5708, B => n5707,
                           ZN => n5711);
   U944 : NAND3_X1 port map( A1 => n5711, A2 => n5710, A3 => n5709, ZN => n5729
                           );
   U945 : AOI222_X1 port map( A1 => n5712, A2 => n6551, B1 => n5758, B2 => 
                           n6549, C1 => n5729, C2 => n6547, ZN => n5931);
   U946 : AOI222_X1 port map( A1 => n5713, A2 => n6551, B1 => n5729, B2 => 
                           n6549, C1 => n5712, C2 => n6547, ZN => n5828);
   U947 : OAI22_X1 port map( A1 => n6292, A2 => n5931, B1 => n5828, B2 => n6181
                           , ZN => n5716);
   U948 : OAI22_X1 port map( A1 => n6561, A2 => n5718, B1 => n5714, B2 => n6295
                           , ZN => n5715);
   U949 : AOI211_X1 port map( C1 => n6232, C2 => n5717, A => n5716, B => n5715,
                           ZN => n5928);
   U950 : OAI22_X1 port map( A1 => n6573, A2 => n5736, B1 => n5928, B2 => n6566
                           , ZN => n5723);
   U951 : OAI22_X1 port map( A1 => n5718, A2 => n6295, B1 => n5759, B2 => n6558
                           , ZN => n5721);
   U952 : OAI22_X1 port map( A1 => n6561, A2 => n5719, B1 => n6557, B2 => n5828
                           , ZN => n5720);
   U953 : AOI211_X1 port map( C1 => n6232, C2 => n5732, A => n5721, B => n5720,
                           ZN => n5832);
   U954 : OAI22_X1 port map( A1 => n5739, A2 => n6450, B1 => n5832, B2 => n6570
                           , ZN => n5722);
   U955 : AOI211_X1 port map( C1 => n6468, C2 => n5724, A => n5723, B => n5722,
                           ZN => n5767);
   U956 : INV_X1 port map( A => n5739, ZN => n5735);
   U957 : INV_X1 port map( A => n5724, ZN => n5763);
   U958 : AOI211_X1 port map( C1 => n5185, C2 => DATA1(28), A => n5726, B => 
                           n5725, ZN => n5728);
   U959 : NAND2_X1 port map( A1 => n6691, A2 => n5785, ZN => n5727);
   U960 : OAI211_X1 port map( C1 => n6113, C2 => n6166, A => n5728, B => n5727,
                           ZN => n5827);
   U961 : AOI222_X1 port map( A1 => n5729, A2 => n6551, B1 => n5827, B2 => 
                           n6549, C1 => n5758, C2 => n6547, ZN => n5941);
   U962 : OAI22_X1 port map( A1 => n6557, A2 => n5941, B1 => n5759, B2 => n6295
                           , ZN => n5731);
   U963 : OAI22_X1 port map( A1 => n5828, A2 => n6554, B1 => n5931, B2 => n6181
                           , ZN => n5730);
   U964 : AOI211_X1 port map( C1 => n6067, C2 => n5732, A => n5731, B => n5730,
                           ZN => n5946);
   U965 : OAI22_X1 port map( A1 => n5763, A2 => n6450, B1 => n5946, B2 => n6566
                           , ZN => n5734);
   U966 : OAI22_X1 port map( A1 => n5832, A2 => n6568, B1 => n5928, B2 => n6570
                           , ZN => n5733);
   U967 : AOI211_X1 port map( C1 => n6072, C2 => n5735, A => n5734, B => n5733,
                           ZN => n5836);
   U968 : OAI22_X1 port map( A1 => n5763, A2 => n6570, B1 => n5832, B2 => n6566
                           , ZN => n5738);
   U969 : OAI22_X1 port map( A1 => n5739, A2 => n6451, B1 => n5736, B2 => n6450
                           , ZN => n5737);
   U970 : AOI211_X1 port map( C1 => n6072, C2 => n5744, A => n5738, B => n5737,
                           ZN => n5748);
   U971 : OAI222_X1 port map( A1 => n6409, A2 => n5767, B1 => n6410, B2 => 
                           n5836, C1 => n5748, C2 => n5983, ZN => n5837);
   U972 : OAI22_X1 port map( A1 => n5739, A2 => n6570, B1 => n5763, B2 => n5224
                           , ZN => n5743);
   U973 : AOI22_X1 port map( A1 => n6072, A2 => n5793, B1 => n5740, B2 => n6468
                           , ZN => n5741);
   U974 : INV_X1 port map( A => n5741, ZN => n5742);
   U975 : AOI211_X1 port map( C1 => n6577, C2 => n5744, A => n5743, B => n5742,
                           ZN => n5749);
   U976 : OAI222_X1 port map( A1 => n6409, A2 => n5748, B1 => n6410, B2 => 
                           n5767, C1 => n5749, C2 => n5983, ZN => n5955);
   U977 : AOI22_X1 port map( A1 => n6472, A2 => n5837, B1 => n6475, B2 => n5955
                           , ZN => n5751);
   U978 : INV_X1 port map( A => n5749, ZN => n5745);
   U979 : AOI222_X1 port map( A1 => n6584, A2 => n5746, B1 => n6582, B2 => 
                           n5745, C1 => n5798, C2 => n6579, ZN => n5813);
   U980 : INV_X1 port map( A => n5813, ZN => n5819);
   U981 : OAI222_X1 port map( A1 => n6409, A2 => n5749, B1 => n6410, B2 => 
                           n5748, C1 => n5747, C2 => n5983, ZN => n5800);
   U982 : AOI22_X1 port map( A1 => n6595, A2 => n5819, B1 => n6470, B2 => n5800
                           , ZN => n5750);
   U983 : OAI211_X1 port map( C1 => n6590, C2 => n5816, A => n5751, B => n5750,
                           ZN => n5962);
   U984 : INV_X1 port map( A => n5962, ZN => n5865);
   U985 : INV_X1 port map( A => n5837, ZN => n5959);
   U986 : INV_X1 port map( A => n5946, ZN => n5766);
   U987 : INV_X1 port map( A => n5941, ZN => n5762);
   U988 : NAND3_X1 port map( A1 => n5754, A2 => n5753, A3 => n5752, ZN => n5755
                           );
   U989 : AOI211_X1 port map( C1 => DATA1(29), C2 => n5825, A => n5756, B => 
                           n5755, ZN => n5757);
   U990 : INV_X1 port map( A => n5757, ZN => n5937);
   U991 : AOI222_X1 port map( A1 => n6549, A2 => n5937, B1 => n6547, B2 => 
                           n5827, C1 => n6551, C2 => n5758, ZN => n5938);
   U992 : OAI22_X1 port map( A1 => n6554, A2 => n5931, B1 => n6557, B2 => n5938
                           , ZN => n5761);
   U993 : OAI22_X1 port map( A1 => n6295, A2 => n5828, B1 => n6561, B2 => n5759
                           , ZN => n5760);
   U994 : AOI211_X1 port map( C1 => n5762, C2 => n6298, A => n5761, B => n5760,
                           ZN => n5930);
   U995 : OAI22_X1 port map( A1 => n6568, A2 => n5928, B1 => n6566, B2 => n5930
                           , ZN => n5765);
   U996 : OAI22_X1 port map( A1 => n6450, A2 => n5832, B1 => n6573, B2 => n5763
                           , ZN => n5764);
   U997 : AOI211_X1 port map( C1 => n5766, C2 => n6073, A => n5765, B => n5764,
                           ZN => n5950);
   U998 : OAI222_X1 port map( A1 => n5767, A2 => n5983, B1 => n5836, B2 => 
                           n6409, C1 => n5950, C2 => n6410, ZN => n5953);
   U999 : AOI22_X1 port map( A1 => n5955, A2 => n5908, B1 => n5953, B2 => n6472
                           , ZN => n5769);
   U1000 : AOI22_X1 port map( A1 => n5985, A2 => n5819, B1 => n5800, B2 => 
                           n6595, ZN => n5768);
   U1001 : OAI211_X1 port map( C1 => n6592, C2 => n5959, A => n5769, B => n5768
                           , ZN => n5961);
   U1002 : INV_X1 port map( A => n5816, ZN => n5861);
   U1003 : INV_X1 port map( A => n5858, ZN => n5797);
   U1004 : OAI211_X1 port map( C1 => n6055, C2 => n5782, A => n5771, B => n5770
                           , ZN => n5772);
   U1005 : AOI211_X1 port map( C1 => n6058, C2 => n5774, A => n5773, B => n5772
                           , ZN => n5804);
   U1006 : OAI222_X1 port map( A1 => n6064, A2 => n5775, B1 => n6063, B2 => 
                           n5786, C1 => n6061, C2 => n5804, ZN => n5852);
   U1007 : INV_X1 port map( A => n5852, ZN => n5871);
   U1008 : OAI22_X1 port map( A1 => n6554, A2 => n5807, B1 => n6561, B2 => 
                           n5871, ZN => n5779);
   U1009 : INV_X1 port map( A => n5787, ZN => n5777);
   U1010 : OAI22_X1 port map( A1 => n6181, A2 => n5777, B1 => n6557, B2 => 
                           n5776, ZN => n5778);
   U1011 : AOI211_X1 port map( C1 => n5853, C2 => n6565, A => n5779, B => n5778
                           , ZN => n5875);
   U1012 : INV_X1 port map( A => n5875, ZN => n5808);
   U1013 : AOI22_X1 port map( A1 => n6565, A2 => n5852, B1 => n6232, B2 => 
                           n5853, ZN => n5789);
   U1014 : NOR2_X1 port map( A1 => n6326, A2 => n6662, ZN => n5784);
   U1015 : OAI211_X1 port map( C1 => n6113, C2 => n5782, A => n5781, B => n5780
                           , ZN => n5783);
   U1016 : AOI211_X1 port map( C1 => DATA1(6), C2 => n5785, A => n5784, B => 
                           n5783, ZN => n5850);
   U1017 : OAI222_X1 port map( A1 => n6064, A2 => n5786, B1 => n6063, B2 => 
                           n5804, C1 => n6061, C2 => n5850, ZN => n5870);
   U1018 : AOI22_X1 port map( A1 => n6067, A2 => n5870, B1 => n6228, B2 => 
                           n5787, ZN => n5788);
   U1019 : OAI211_X1 port map( C1 => n5807, C2 => n6558, A => n5789, B => n5788
                           , ZN => n5892);
   U1020 : AOI22_X1 port map( A1 => n6577, A2 => n5808, B1 => n6302, B2 => 
                           n5892, ZN => n5791);
   U1021 : AOI22_X1 port map( A1 => n6495, A2 => n5792, B1 => n6526, B2 => 
                           n5794, ZN => n5790);
   U1022 : OAI211_X1 port map( C1 => n5797, C2 => n6451, A => n5791, B => n5790
                           , ZN => n5847);
   U1023 : AOI22_X1 port map( A1 => n6468, A2 => n5792, B1 => n6302, B2 => 
                           n5808, ZN => n5796);
   U1024 : AOI22_X1 port map( A1 => n6073, A2 => n5794, B1 => n6526, B2 => 
                           n5793, ZN => n5795);
   U1025 : OAI211_X1 port map( C1 => n5797, C2 => n6450, A => n5796, B => n5795
                           , ZN => n5812);
   U1026 : AOI222_X1 port map( A1 => n5847, A2 => n6579, B1 => n5812, B2 => 
                           n6584, C1 => n5799, C2 => n6582, ZN => n5803);
   U1027 : AOI222_X1 port map( A1 => n5812, A2 => n6579, B1 => n5799, B2 => 
                           n6584, C1 => n5798, C2 => n6582, ZN => n5882);
   U1028 : OAI22_X1 port map( A1 => n6590, A2 => n5803, B1 => n5882, B2 => 
                           n6310, ZN => n5802);
   U1029 : INV_X1 port map( A => n5800, ZN => n5840);
   U1030 : OAI22_X1 port map( A1 => n5813, A2 => n6592, B1 => n5840, B2 => 
                           n6307, ZN => n5801);
   U1031 : AOI211_X1 port map( C1 => n6470, C2 => n5861, A => n5802, B => n5801
                           , ZN => n5864);
   U1032 : INV_X1 port map( A => n5864, ZN => n5919);
   U1033 : AOI22_X1 port map( A1 => n6509, A2 => n5961, B1 => n5919, B2 => 
                           n6603, ZN => n5821);
   U1034 : INV_X1 port map( A => n5803, ZN => n5897);
   U1035 : AOI22_X1 port map( A1 => n6565, A2 => n5870, B1 => n6232, B2 => 
                           n5852, ZN => n5806);
   U1036 : OAI222_X1 port map( A1 => n6064, A2 => n5804, B1 => n6063, B2 => 
                           n5850, C1 => n6061, C2 => n5849, ZN => n5886);
   U1037 : AOI22_X1 port map( A1 => n6230, A2 => n5853, B1 => n6067, B2 => 
                           n5886, ZN => n5805);
   U1038 : OAI211_X1 port map( C1 => n6292, C2 => n5807, A => n5806, B => n5805
                           , ZN => n5848);
   U1039 : AOI22_X1 port map( A1 => n6468, A2 => n5808, B1 => n6302, B2 => 
                           n5848, ZN => n5810);
   U1040 : AOI22_X1 port map( A1 => n6577, A2 => n5892, B1 => n6495, B2 => 
                           n5858, ZN => n5809);
   U1041 : OAI211_X1 port map( C1 => n5811, C2 => n6566, A => n5810, B => n5809
                           , ZN => n5846);
   U1042 : AOI222_X1 port map( A1 => n5846, A2 => n6579, B1 => n5847, B2 => 
                           n6584, C1 => n5812, C2 => n6582, ZN => n5911);
   U1043 : OAI22_X1 port map( A1 => n6590, A2 => n5911, B1 => n5816, B2 => 
                           n6592, ZN => n5815);
   U1044 : OAI22_X1 port map( A1 => n5882, A2 => n6586, B1 => n5813, B2 => 
                           n6307, ZN => n5814);
   U1045 : AOI211_X1 port map( C1 => n6595, C2 => n5897, A => n5815, B => n5814
                           , ZN => n5914);
   U1046 : INV_X1 port map( A => n5914, ZN => n5918);
   U1047 : INV_X1 port map( A => n5955, ZN => n5839);
   U1048 : OAI22_X1 port map( A1 => n5816, A2 => n6310, B1 => n5839, B2 => 
                           n6588, ZN => n5818);
   U1049 : OAI22_X1 port map( A1 => n6590, A2 => n5882, B1 => n5840, B2 => 
                           n6592, ZN => n5817);
   U1050 : AOI211_X1 port map( C1 => n6470, C2 => n5819, A => n5818, B => n5817
                           , ZN => n5922);
   U1051 : INV_X1 port map( A => n5922, ZN => n5963);
   U1052 : AOI22_X1 port map( A1 => n5918, A2 => n6605, B1 => n5963, B2 => 
                           n6236, ZN => n5820);
   U1053 : OAI211_X1 port map( C1 => n6608, C2 => n5865, A => n5821, B => n5820
                           , ZN => n5969);
   U1054 : INV_X1 port map( A => n6509, ZN => n6598);
   U1055 : INV_X1 port map( A => n5930, ZN => n5835);
   U1056 : INV_X1 port map( A => n5938, ZN => n5831);
   U1057 : NOR2_X1 port map( A1 => n6283, A2 => n6095, ZN => n6117);
   U1058 : OAI211_X1 port map( C1 => n6113, C2 => n6136, A => n5823, B => n5822
                           , ZN => n5824);
   U1059 : AOI211_X1 port map( C1 => DATA1(30), C2 => n5825, A => n6117, B => 
                           n5824, ZN => n5826);
   U1060 : INV_X1 port map( A => n5826, ZN => n5935);
   U1061 : AOI222_X1 port map( A1 => n6549, A2 => n5935, B1 => n6547, B2 => 
                           n5937, C1 => n6551, C2 => n5827, ZN => n5940);
   U1062 : OAI22_X1 port map( A1 => n6554, A2 => n5941, B1 => n6557, B2 => 
                           n5940, ZN => n5830);
   U1063 : OAI22_X1 port map( A1 => n6295, A2 => n5931, B1 => n6561, B2 => 
                           n5828, ZN => n5829);
   U1064 : AOI211_X1 port map( C1 => n5831, C2 => n6230, A => n5830, B => n5829
                           , ZN => n5929);
   U1065 : OAI22_X1 port map( A1 => n6568, A2 => n5946, B1 => n6566, B2 => 
                           n5929, ZN => n5834);
   U1066 : OAI22_X1 port map( A1 => n6450, A2 => n5928, B1 => n6573, B2 => 
                           n5832, ZN => n5833);
   U1067 : AOI211_X1 port map( C1 => n5835, C2 => n6073, A => n5834, B => n5833
                           , ZN => n5952);
   U1068 : OAI222_X1 port map( A1 => n5836, A2 => n5983, B1 => n5950, B2 => 
                           n6409, C1 => n5952, C2 => n6410, ZN => n5956);
   U1069 : AOI22_X1 port map( A1 => n5837, A2 => n6470, B1 => n5956, B2 => 
                           n6472, ZN => n5838);
   U1070 : INV_X1 port map( A => n5838, ZN => n5842);
   U1071 : OAI22_X1 port map( A1 => n6590, A2 => n5840, B1 => n5839, B2 => 
                           n6310, ZN => n5841);
   U1072 : AOI211_X1 port map( C1 => n6475, C2 => n5953, A => n5842, B => n5841
                           , ZN => n5966);
   U1073 : OAI22_X1 port map( A1 => n6598, A2 => n5966, B1 => n5865, B2 => 
                           n6600, ZN => n5844);
   U1074 : OAI22_X1 port map( A1 => n5922, A2 => n6083, B1 => n5864, B2 => 
                           n6081, ZN => n5843);
   U1075 : AOI211_X1 port map( C1 => n6518, C2 => n5961, A => n5844, B => n5843
                           , ZN => n5845);
   U1076 : INV_X1 port map( A => n5845, ZN => n5968);
   U1077 : INV_X1 port map( A => n5846, ZN => n5879);
   U1078 : INV_X1 port map( A => n5847, ZN => n5859);
   U1079 : INV_X1 port map( A => n5892, ZN => n5874);
   U1080 : INV_X1 port map( A => n5848, ZN => n5904);
   U1081 : OAI22_X1 port map( A1 => n5874, A2 => n6451, B1 => n5904, B2 => 
                           n6450, ZN => n5857);
   U1082 : INV_X1 port map( A => n5886, ZN => n5900);
   U1083 : OAI222_X1 port map( A1 => n5851, A2 => n6061, B1 => n5850, B2 => 
                           n6064, C1 => n5849, C2 => n6063, ZN => n5884);
   U1084 : AOI22_X1 port map( A1 => n6067, A2 => n5884, B1 => n5870, B2 => 
                           n6232, ZN => n5855);
   U1085 : AOI22_X1 port map( A1 => n6197, A2 => n5853, B1 => n5852, B2 => 
                           n6230, ZN => n5854);
   U1086 : OAI211_X1 port map( C1 => n6295, C2 => n5900, A => n5855, B => n5854
                           , ZN => n5878);
   U1087 : INV_X1 port map( A => n5878, ZN => n5980);
   U1088 : OAI22_X1 port map( A1 => n6573, A2 => n5980, B1 => n5875, B2 => 
                           n6570, ZN => n5856);
   U1089 : AOI211_X1 port map( C1 => n6526, C2 => n5858, A => n5857, B => n5856
                           , ZN => n5893);
   U1090 : OAI222_X1 port map( A1 => n6409, A2 => n5879, B1 => n6410, B2 => 
                           n5859, C1 => n5893, C2 => n5983, ZN => n5986);
   U1091 : AOI22_X1 port map( A1 => n5908, A2 => n5897, B1 => n5985, B2 => 
                           n5986, ZN => n5863);
   U1092 : INV_X1 port map( A => n5882, ZN => n5860);
   U1093 : AOI22_X1 port map( A1 => n6472, A2 => n5861, B1 => n6475, B2 => 
                           n5860, ZN => n5862);
   U1094 : OAI211_X1 port map( C1 => n5911, C2 => n6310, A => n5863, B => n5862
                           , ZN => n5990);
   U1095 : OAI22_X1 port map( A1 => n6598, A2 => n5865, B1 => n5864, B2 => 
                           n6600, ZN => n5867);
   U1096 : OAI22_X1 port map( A1 => n5914, A2 => n6083, B1 => n5922, B2 => 
                           n6608, ZN => n5866);
   U1097 : AOI211_X1 port map( C1 => n6316, C2 => n5990, A => n5867, B => n5866
                           , ZN => n5868);
   U1098 : INV_X1 port map( A => n5868, ZN => n5924);
   U1099 : AOI222_X1 port map( A1 => n6089, A2 => n5969, B1 => n6610, B2 => 
                           n5968, C1 => n5924, C2 => n6615, ZN => n5869);
   U1100 : INV_X1 port map( A => n5869, ZN => n5997);
   U1101 : INV_X1 port map( A => n5911, ZN => n5883);
   U1102 : INV_X1 port map( A => n5870, ZN => n5889);
   U1103 : INV_X1 port map( A => n5884, ZN => n5974);
   U1104 : OAI22_X1 port map( A1 => n5889, A2 => n6558, B1 => n5974, B2 => 
                           n6295, ZN => n5873);
   U1105 : OAI22_X1 port map( A1 => n6292, A2 => n5871, B1 => n5900, B2 => 
                           n6554, ZN => n5872);
   U1106 : AOI211_X1 port map( C1 => n6067, C2 => n5885, A => n5873, B => n5872
                           , ZN => n6449);
   U1107 : OAI22_X1 port map( A1 => n6573, A2 => n6449, B1 => n5904, B2 => 
                           n6451, ZN => n5877);
   U1108 : OAI22_X1 port map( A1 => n5875, A2 => n5224, B1 => n5874, B2 => 
                           n6570, ZN => n5876);
   U1109 : AOI211_X1 port map( C1 => n6577, C2 => n5878, A => n5877, B => n5876
                           , ZN => n5907);
   U1110 : OAI222_X1 port map( A1 => n6409, A2 => n5893, B1 => n6410, B2 => 
                           n5879, C1 => n5907, C2 => n5983, ZN => n6333);
   U1111 : AOI22_X1 port map( A1 => n6470, A2 => n5883, B1 => n5985, B2 => 
                           n6333, ZN => n5881);
   U1112 : AOI22_X1 port map( A1 => n6475, A2 => n5897, B1 => n6595, B2 => 
                           n5986, ZN => n5880);
   U1113 : OAI211_X1 port map( C1 => n5882, C2 => n6307, A => n5881, B => n5880
                           , ZN => n6218);
   U1114 : AOI22_X1 port map( A1 => n5883, A2 => n6475, B1 => n5986, B2 => 
                           n6470, ZN => n5896);
   U1115 : AOI22_X1 port map( A1 => n6565, A2 => n5885, B1 => n6232, B2 => 
                           n5884, ZN => n5888);
   U1116 : AOI22_X1 port map( A1 => n6298, A2 => n5886, B1 => n6067, B2 => 
                           n5903, ZN => n5887);
   U1117 : OAI211_X1 port map( C1 => n6292, C2 => n5889, A => n5888, B => n5887
                           , ZN => n6467);
   U1118 : INV_X1 port map( A => n6467, ZN => n6448);
   U1119 : OAI22_X1 port map( A1 => n6451, A2 => n5980, B1 => n6573, B2 => 
                           n6448, ZN => n5891);
   U1120 : OAI22_X1 port map( A1 => n6450, A2 => n6449, B1 => n6570, B2 => 
                           n5904, ZN => n5890);
   U1121 : AOI211_X1 port map( C1 => n5892, C2 => n6526, A => n5891, B => n5890
                           , ZN => n5984);
   U1122 : OAI222_X1 port map( A1 => n5984, A2 => n5894, B1 => n5907, B2 => 
                           n6409, C1 => n5893, C2 => n6410, ZN => n6350);
   U1123 : AOI22_X1 port map( A1 => n5985, A2 => n6350, B1 => n6333, B2 => 
                           n6595, ZN => n5895);
   U1124 : NAND2_X1 port map( A1 => n5896, A2 => n5895, ZN => n5915);
   U1125 : AOI21_X1 port map( B1 => n5897, B2 => n6472, A => n5915, ZN => n5898
                           );
   U1126 : INV_X1 port map( A => n5898, ZN => n6237);
   U1127 : AOI22_X1 port map( A1 => n6236, A2 => n6218, B1 => n6603, B2 => 
                           n6237, ZN => n5913);
   U1128 : OAI22_X1 port map( A1 => n6561, A2 => n5899, B1 => n5974, B2 => 
                           n6558, ZN => n5902);
   U1129 : OAI22_X1 port map( A1 => n6557, A2 => n5900, B1 => n5975, B2 => 
                           n6554, ZN => n5901);
   U1130 : AOI211_X1 port map( C1 => n6565, C2 => n5903, A => n5902, B => n5901
                           , ZN => n6452);
   U1131 : OAI22_X1 port map( A1 => n6573, A2 => n6452, B1 => n6449, B2 => 
                           n6568, ZN => n5906);
   U1132 : OAI22_X1 port map( A1 => n5904, A2 => n5224, B1 => n5980, B2 => 
                           n6570, ZN => n5905);
   U1133 : AOI211_X1 port map( C1 => n6577, C2 => n6467, A => n5906, B => n5905
                           , ZN => n6411);
   U1134 : OAI222_X1 port map( A1 => n6409, A2 => n5984, B1 => n6410, B2 => 
                           n5907, C1 => n6411, C2 => n5983, ZN => n6372);
   U1135 : AOI22_X1 port map( A1 => n5908, A2 => n6333, B1 => n5985, B2 => 
                           n6372, ZN => n5910);
   U1136 : AOI22_X1 port map( A1 => n6475, A2 => n5986, B1 => n6595, B2 => 
                           n6350, ZN => n5909);
   U1137 : OAI211_X1 port map( C1 => n5911, C2 => n6307, A => n5910, B => n5909
                           , ZN => n6247);
   U1138 : AOI22_X1 port map( A1 => n6316, A2 => n6247, B1 => n6518, B2 => 
                           n5990, ZN => n5912);
   U1139 : OAI211_X1 port map( C1 => n6598, C2 => n5914, A => n5913, B => n5912
                           , ZN => n6165);
   U1140 : INV_X1 port map( A => n6218, ZN => n5993);
   U1141 : AOI22_X1 port map( A1 => n6605, A2 => n5915, B1 => n6516, B2 => 
                           n5919, ZN => n5917);
   U1142 : AOI22_X1 port map( A1 => n6315, A2 => n5990, B1 => n6518, B2 => 
                           n5918, ZN => n5916);
   U1143 : OAI211_X1 port map( C1 => n5993, C2 => n6083, A => n5917, B => n5916
                           , ZN => n5994);
   U1144 : AOI22_X1 port map( A1 => n6316, A2 => n6218, B1 => n6236, B2 => 
                           n5918, ZN => n5921);
   U1145 : AOI22_X1 port map( A1 => n6603, A2 => n5990, B1 => n6518, B2 => 
                           n5919, ZN => n5920);
   U1146 : OAI211_X1 port map( C1 => n6598, C2 => n5922, A => n5921, B => n5920
                           , ZN => n5925);
   U1147 : AOI222_X1 port map( A1 => n5923, A2 => n6165, B1 => n5994, B2 => 
                           n6612, C1 => n5925, C2 => n6610, ZN => n6140);
   U1148 : AOI222_X1 port map( A1 => n5923, A2 => n5925, B1 => n5924, B2 => 
                           n6089, C1 => n5969, C2 => n6610, ZN => n6101);
   U1149 : OAI22_X1 port map( A1 => n6140, A2 => n6622, B1 => n6101, B2 => 
                           n6618, ZN => n5972);
   U1150 : AOI222_X1 port map( A1 => n6615, A2 => n5994, B1 => n5925, B2 => 
                           n6612, C1 => n5924, C2 => n6321, ZN => n6118);
   U1151 : NAND2_X1 port map( A1 => n5927, A2 => n5926, ZN => n6620);
   U1152 : INV_X1 port map( A => n5928, ZN => n5949);
   U1153 : OAI22_X1 port map( A1 => n5930, A2 => n6568, B1 => n5929, B2 => 
                           n6570, ZN => n5948);
   U1154 : INV_X1 port map( A => n5931, ZN => n5944);
   U1155 : INV_X1 port map( A => DATA1(30), ZN => n6686);
   U1156 : NOR2_X1 port map( A1 => n6283, A2 => n6686, ZN => n6096);
   U1157 : AOI211_X1 port map( C1 => n5185, C2 => DATA1(31), A => n5932, B => 
                           n6096, ZN => n5934);
   U1158 : OAI211_X1 port map( C1 => n6055, C2 => n6136, A => n5934, B => n5933
                           , ZN => n5936);
   U1159 : AOI222_X1 port map( A1 => n5937, A2 => n6551, B1 => n5936, B2 => 
                           n6549, C1 => n5935, C2 => n6547, ZN => n5939);
   U1160 : OAI22_X1 port map( A1 => n6292, A2 => n5939, B1 => n5938, B2 => 
                           n6554, ZN => n5943);
   U1161 : OAI22_X1 port map( A1 => n5941, A2 => n6295, B1 => n5940, B2 => 
                           n6181, ZN => n5942);
   U1162 : AOI211_X1 port map( C1 => n6067, C2 => n5944, A => n5943, B => n5942
                           , ZN => n5945);
   U1163 : OAI22_X1 port map( A1 => n5946, A2 => n6450, B1 => n5945, B2 => 
                           n6566, ZN => n5947);
   U1164 : AOI211_X1 port map( C1 => n6302, C2 => n5949, A => n5948, B => n5947
                           , ZN => n5951);
   U1165 : OAI222_X1 port map( A1 => n6409, A2 => n5952, B1 => n6410, B2 => 
                           n5951, C1 => n5950, C2 => n5983, ZN => n5954);
   U1166 : AOI22_X1 port map( A1 => n6472, A2 => n5954, B1 => n6470, B2 => 
                           n5953, ZN => n5958);
   U1167 : AOI22_X1 port map( A1 => n6475, A2 => n5956, B1 => n5985, B2 => 
                           n5955, ZN => n5957);
   U1168 : OAI211_X1 port map( C1 => n5959, C2 => n6310, A => n5958, B => n5957
                           , ZN => n5960);
   U1169 : AOI22_X1 port map( A1 => n6236, A2 => n5961, B1 => n6516, B2 => 
                           n5960, ZN => n5965);
   U1170 : AOI22_X1 port map( A1 => n6316, A2 => n5963, B1 => n6603, B2 => 
                           n5962, ZN => n5964);
   U1171 : OAI211_X1 port map( C1 => n5966, C2 => n6608, A => n5965, B => n5964
                           , ZN => n5967);
   U1172 : AOI222_X1 port map( A1 => n6615, A2 => n5969, B1 => n5968, B2 => 
                           n6089, C1 => n5967, C2 => n6610, ZN => n5970);
   U1173 : OAI22_X1 port map( A1 => n6118, A2 => n6620, B1 => n5970, B2 => 
                           n6616, ZN => n5971);
   U1174 : AOI211_X1 port map( C1 => n6627, C2 => n5997, A => n5972, B => n5971
                           , ZN => n6029);
   U1175 : OAI22_X1 port map( A1 => n6140, A2 => n6620, B1 => n6101, B2 => 
                           n6139, ZN => n5996);
   U1176 : INV_X1 port map( A => n6333, ZN => n5989);
   U1177 : INV_X1 port map( A => n6452, ZN => n6494);
   U1178 : OAI22_X1 port map( A1 => n6557, A2 => n5974, B1 => n5973, B2 => 
                           n6554, ZN => n5978);
   U1179 : OAI22_X1 port map( A1 => n6561, A2 => n5976, B1 => n5975, B2 => 
                           n6558, ZN => n5977);
   U1180 : AOI211_X1 port map( C1 => n6565, C2 => n5979, A => n5978, B => n5977
                           , ZN => n6466);
   U1181 : OAI22_X1 port map( A1 => n6573, A2 => n6466, B1 => n6448, B2 => 
                           n6451, ZN => n5982);
   U1182 : OAI22_X1 port map( A1 => n5980, A2 => n5224, B1 => n6449, B2 => 
                           n6570, ZN => n5981);
   U1183 : AOI211_X1 port map( C1 => n6577, C2 => n6494, A => n5982, B => n5981
                           , ZN => n6431);
   U1184 : OAI222_X1 port map( A1 => n6409, A2 => n6411, B1 => n6410, B2 => 
                           n5984, C1 => n6431, C2 => n5983, ZN => n6390);
   U1185 : AOI22_X1 port map( A1 => n6595, A2 => n6372, B1 => n5985, B2 => 
                           n6390, ZN => n5988);
   U1186 : AOI22_X1 port map( A1 => n6472, A2 => n5986, B1 => n6470, B2 => 
                           n6350, ZN => n5987);
   U1187 : OAI211_X1 port map( C1 => n5989, C2 => n6592, A => n5988, B => n5987
                           , ZN => n6271);
   U1188 : AOI22_X1 port map( A1 => n6605, A2 => n6271, B1 => n6603, B2 => 
                           n6247, ZN => n5992);
   U1189 : AOI22_X1 port map( A1 => n6236, A2 => n6237, B1 => n6516, B2 => 
                           n5990, ZN => n5991);
   U1190 : OAI211_X1 port map( C1 => n5993, C2 => n6608, A => n5992, B => n5991
                           , ZN => n6191);
   U1191 : AOI222_X1 port map( A1 => n6615, A2 => n6191, B1 => n6165, B2 => 
                           n6612, C1 => n5994, C2 => n6610, ZN => n6158);
   U1192 : OAI22_X1 port map( A1 => n6118, A2 => n6618, B1 => n6158, B2 => 
                           n6622, ZN => n5995);
   U1193 : AOI211_X1 port map( C1 => n5998, C2 => n5997, A => n5996, B => n5995
                           , ZN => n6041);
   U1194 : OR3_X1 port map( A1 => n6867, A2 => n6622, A3 => n5999, ZN => n6628)
                           ;
   U1195 : NOR3_X1 port map( A1 => FUNC(3), A2 => n6041, A3 => n6628, ZN => 
                           n6023);
   U1196 : INV_X1 port map( A => DATA2_I_31_port, ZN => n6012);
   U1197 : NAND2_X1 port map( A1 => n6689, A2 => n6012, ZN => n6019);
   U1198 : INV_X1 port map( A => n6019, ZN => n6021);
   U1199 : NAND2_X1 port map( A1 => DATA1(30), A2 => DATA2_I_30_port, ZN => 
                           n6013);
   U1200 : NAND2_X1 port map( A1 => DATA1(29), A2 => DATA2_I_29_port, ZN => 
                           n6014);
   U1201 : INV_X1 port map( A => n6014, ZN => n6038);
   U1202 : XOR2_X1 port map( A => DATA2_I_23_port, B => DATA1(23), Z => n6217);
   U1203 : NAND2_X1 port map( A1 => DATA1(22), A2 => DATA2_I_22_port, ZN => 
                           n6213);
   U1204 : OAI21_X1 port map( B1 => n6753, B2 => DATA2_I_22_port, A => n6213, 
                           ZN => n6234);
   U1205 : XOR2_X1 port map( A => DATA2_I_21_port, B => DATA1(21), Z => n6258);
   U1206 : NAND2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n6387);
   U1207 : INV_X1 port map( A => n6387, ZN => n6373);
   U1208 : XOR2_X1 port map( A => DATA2_I_17_port, B => DATA1(17), Z => n6383);
   U1209 : AOI22_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, B1 => 
                           n6373, B2 => n6383, ZN => n6355);
   U1210 : NAND2_X1 port map( A1 => DATA1(18), A2 => DATA2_I_18_port, ZN => 
                           n6203);
   U1211 : OAI21_X1 port map( B1 => DATA1(18), B2 => DATA2_I_18_port, A => 
                           n6203, ZN => n6367);
   U1212 : OAI21_X1 port map( B1 => n6355, B2 => n6367, A => n6203, ZN => n6335
                           );
   U1213 : OR2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => n6206
                           );
   U1214 : AOI22_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, B1 => 
                           n6335, B2 => n6206, ZN => n6266);
   U1215 : NAND2_X1 port map( A1 => DATA1(20), A2 => DATA2_I_20_port, ZN => 
                           n6207);
   U1216 : OAI21_X1 port map( B1 => DATA1(20), B2 => DATA2_I_20_port, A => 
                           n6207, ZN => n6267);
   U1217 : OAI21_X1 port map( B1 => n6266, B2 => n6267, A => n6207, ZN => n6253
                           );
   U1218 : AOI22_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, B1 => 
                           n6258, B2 => n6253, ZN => n6214);
   U1219 : NOR2_X1 port map( A1 => DATA1(16), A2 => DATA2_I_16_port, ZN => 
                           n6374);
   U1220 : INV_X1 port map( A => n6383, ZN => n6381);
   U1221 : NOR2_X1 port map( A1 => n6374, A2 => n6381, ZN => n6201);
   U1222 : INV_X1 port map( A => n6258, ZN => n6255);
   U1223 : NAND2_X1 port map( A1 => DATA1(19), A2 => DATA2_I_19_port, ZN => 
                           n6204);
   U1224 : OAI21_X1 port map( B1 => DATA1(19), B2 => DATA2_I_19_port, A => 
                           n6204, ZN => n6344);
   U1225 : NOR4_X1 port map( A1 => n6367, A2 => n6267, A3 => n6255, A4 => n6344
                           , ZN => n6007);
   U1226 : NAND2_X1 port map( A1 => DATA1(15), A2 => DATA2_I_15_port, ZN => 
                           n6005);
   U1227 : OAI21_X1 port map( B1 => DATA1(15), B2 => DATA2_I_15_port, A => 
                           n6005, ZN => n6405);
   U1228 : XOR2_X1 port map( A => DATA2_I_14_port, B => n7169, Z => n6439);
   U1229 : NAND2_X1 port map( A1 => DATA1(13), A2 => DATA2_I_13_port, ZN => 
                           n6435);
   U1230 : OAI21_X1 port map( B1 => DATA1(13), B2 => DATA2_I_13_port, A => 
                           n6435, ZN => n6463);
   U1231 : NAND2_X1 port map( A1 => n7168, A2 => DATA2_I_12_port, ZN => n6464);
   U1232 : OAI21_X1 port map( B1 => DATA1(12), B2 => DATA2_I_12_port, A => 
                           n6464, ZN => n6479);
   U1233 : NOR2_X1 port map( A1 => n6463, A2 => n6479, ZN => n6418);
   U1234 : NOR2_X1 port map( A1 => n6000, A2 => DATA2_I_11_port, ZN => n6416);
   U1235 : NAND2_X1 port map( A1 => DATA1(9), A2 => DATA2_I_9_port, ZN => n6519
                           );
   U1236 : NAND2_X1 port map( A1 => DATA1(10), A2 => DATA2_I_10_port, ZN => 
                           n6414);
   U1237 : OAI21_X1 port map( B1 => n7167, B2 => DATA2_I_10_port, A => n6414, 
                           ZN => n6520);
   U1238 : AOI21_X1 port map( B1 => n6519, B2 => n6523, A => n6520, ZN => n6522
                           );
   U1239 : AOI21_X1 port map( B1 => DATA2_I_10_port, B2 => n7167, A => n6522, 
                           ZN => n6508);
   U1240 : NAND2_X1 port map( A1 => n6000, A2 => DATA2_I_11_port, ZN => n6415);
   U1241 : OAI21_X1 port map( B1 => n6416, B2 => n6508, A => n6415, ZN => n6478
                           );
   U1242 : NOR2_X1 port map( A1 => n6464, A2 => n6463, ZN => n6417);
   U1243 : AOI21_X1 port map( B1 => n6418, B2 => n6478, A => n6417, ZN => n6437
                           );
   U1244 : NAND2_X1 port map( A1 => n6437, A2 => n6435, ZN => n6432);
   U1245 : AOI22_X1 port map( A1 => n7169, A2 => DATA2_I_14_port, B1 => n6439, 
                           B2 => n6432, ZN => n6404);
   U1246 : INV_X1 port map( A => n6439, ZN => n6001);
   U1247 : OAI21_X1 port map( B1 => DATA1(11), B2 => DATA2_I_11_port, A => 
                           n6415, ZN => n6507);
   U1248 : NOR4_X1 port map( A1 => n6520, A2 => n6002, A3 => n6001, A4 => n6507
                           , ZN => n6003);
   U1249 : NAND4_X1 port map( A1 => n6418, A2 => n6004, A3 => n6003, A4 => 
                           n6457, ZN => n6006);
   U1250 : OAI221_X1 port map( B1 => n6405, B2 => n6404, C1 => n6405, C2 => 
                           n6006, A => n6005, ZN => n6210);
   U1251 : NAND3_X1 port map( A1 => n6201, A2 => n6007, A3 => n6210, ZN => 
                           n6008);
   U1252 : OAI221_X1 port map( B1 => n6234, B2 => n6214, C1 => n6234, C2 => 
                           n6008, A => n6213, ZN => n6009);
   U1253 : AOI22_X1 port map( A1 => DATA1(23), A2 => DATA2_I_23_port, B1 => 
                           n6217, B2 => n6009, ZN => n6010);
   U1254 : NOR2_X1 port map( A1 => n6010, A2 => n7166, ZN => n6173);
   U1255 : NAND2_X1 port map( A1 => DATA1(28), A2 => DATA2_I_28_port, ZN => 
                           n6104);
   U1256 : INV_X1 port map( A => n6104, ZN => n6011);
   U1257 : XOR2_X1 port map( A => DATA2_I_26_port, B => DATA1(26), Z => n6164);
   U1258 : NAND2_X1 port map( A1 => DATA1(25), A2 => DATA2_I_25_port, ZN => 
                           n6157);
   U1259 : XOR2_X1 port map( A => DATA2_I_25_port, B => DATA1(25), Z => n6176);
   U1260 : INV_X1 port map( A => DATA2_I_24_port, ZN => n6180);
   U1261 : NAND2_X1 port map( A1 => n6680, A2 => n6180, ZN => n6195);
   U1262 : NAND2_X1 port map( A1 => n6176, A2 => n6195, ZN => n6172);
   U1263 : NAND2_X1 port map( A1 => n6157, A2 => n6172, ZN => n6148);
   U1264 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, B1 => 
                           n6164, B2 => n6148, ZN => n6133);
   U1265 : NAND2_X1 port map( A1 => DATA1(27), A2 => DATA2_I_27_port, ZN => 
                           n6121);
   U1266 : OAI21_X1 port map( B1 => DATA1(27), B2 => DATA2_I_27_port, A => 
                           n6121, ZN => n6145);
   U1267 : OAI21_X1 port map( B1 => DATA1(28), B2 => DATA2_I_28_port, A => 
                           n6104, ZN => n6126);
   U1268 : AOI221_X1 port map( B1 => n6133, B2 => n6121, C1 => n6145, C2 => 
                           n6121, A => n6126, ZN => n6120);
   U1269 : XOR2_X1 port map( A => DATA2_I_29_port, B => DATA1(29), Z => n6111);
   U1270 : OAI21_X1 port map( B1 => n6011, B2 => n6120, A => n6111, ZN => n6016
                           );
   U1271 : NAND2_X1 port map( A1 => n6833, A2 => n6010, ZN => n6125);
   U1272 : INV_X1 port map( A => n6125, ZN => n6186);
   U1273 : NAND3_X1 port map( A1 => n6691, A2 => DATA2_I_24_port, A3 => n6176, 
                           ZN => n6167);
   U1274 : NAND2_X1 port map( A1 => n6157, A2 => n6167, ZN => n6147);
   U1275 : AOI22_X1 port map( A1 => DATA1(26), A2 => DATA2_I_26_port, B1 => 
                           n6164, B2 => n6147, ZN => n6132);
   U1276 : AOI221_X1 port map( B1 => n6132, B2 => n6121, C1 => n6145, C2 => 
                           n6121, A => n6126, ZN => n6119);
   U1277 : OAI21_X1 port map( B1 => n6011, B2 => n6119, A => n6111, ZN => n6015
                           );
   U1278 : AOI22_X1 port map( A1 => n6173, A2 => n6016, B1 => n6186, B2 => 
                           n6015, ZN => n6102);
   U1279 : XOR2_X1 port map( A => DATA2_I_30_port, B => DATA1(30), Z => n6037);
   U1280 : OAI22_X1 port map( A1 => n6038, A2 => n6102, B1 => n6037, B2 => 
                           n7166, ZN => n6036);
   U1281 : OAI211_X1 port map( C1 => n6012, C2 => n6689, A => n6013, B => n6036
                           , ZN => n6020);
   U1282 : INV_X1 port map( A => n6037, ZN => n6035);
   U1283 : OAI21_X1 port map( B1 => n6014, B2 => n6035, A => n6013, ZN => n6017
                           );
   U1284 : INV_X1 port map( A => n6173, ZN => n6194);
   U1285 : OAI22_X1 port map( A1 => n6194, A2 => n6016, B1 => n6125, B2 => 
                           n6015, ZN => n6034);
   U1286 : AOI22_X1 port map( A1 => n6833, A2 => n6017, B1 => n6037, B2 => 
                           n6034, ZN => n6024);
   U1287 : OAI211_X1 port map( C1 => n6689, C2 => n6832, A => DATA2(31), B => 
                           n6631, ZN => n6018);
   U1288 : OAI221_X1 port map( B1 => n6021, B2 => n6020, C1 => n6019, C2 => 
                           n6024, A => n6018, ZN => n6022);
   U1289 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_31_port, A => 
                           n6023, B => n6022, ZN => n6028);
   U1290 : INV_X1 port map( A => DATA2(31), ZN => n6834);
   U1291 : NAND2_X1 port map( A1 => n5185, A2 => n6510, ZN => n6114);
   U1292 : OAI221_X1 port map( B1 => DATA2(31), B2 => n6531, C1 => n6834, C2 =>
                           n6389, A => n6114, ZN => n6026);
   U1293 : INV_X1 port map( A => n6024, ZN => n6025);
   U1294 : OAI221_X1 port map( B1 => n6026, B2 => DATA2_I_31_port, C1 => n6026,
                           C2 => n6025, A => DATA1(31), ZN => n6027);
   U1295 : OAI211_X1 port map( C1 => n6029, C2 => n6496, A => n6028, B => n6027
                           , ZN => OUTALU(31));
   U1296 : INV_X1 port map( A => DATA2(30), ZN => n6835);
   U1297 : OAI22_X1 port map( A1 => n6686, A2 => n6835, B1 => DATA2(30), B2 => 
                           DATA1(30), ZN => n6684);
   U1298 : OAI21_X1 port map( B1 => n6149, B2 => n6835, A => n6114, ZN => n6030
                           );
   U1299 : AOI22_X1 port map( A1 => DATA1(30), A2 => n6030, B1 => n6183, B2 => 
                           dataout_mul_30_port, ZN => n6032);
   U1300 : NAND3_X1 port map( A1 => n6044, A2 => n6510, A3 => DATA1(31), ZN => 
                           n6031);
   U1301 : OAI211_X1 port map( C1 => n6684, C2 => n6531, A => n6032, B => n6031
                           , ZN => n6033);
   U1302 : AOI21_X1 port map( B1 => n6035, B2 => n6034, A => n6033, ZN => n6040
                           );
   U1303 : OAI21_X1 port map( B1 => n6038, B2 => n6037, A => n6036, ZN => n6039
                           );
   U1304 : OAI211_X1 port map( C1 => n6041, C2 => n6496, A => n6040, B => n6039
                           , ZN => OUTALU(30));
   U1305 : OAI22_X1 port map( A1 => n6046, A2 => n6637, B1 => n6045, B2 => 
                           n6042, ZN => n6043);
   U1306 : AOI22_X1 port map( A1 => n6501, A2 => dataout_mul_2_port, B1 => 
                           n6048, B2 => n6043, ZN => n6094);
   U1307 : INV_X1 port map( A => DATA1(0), ZN => n6696);
   U1308 : NAND2_X1 port map( A1 => n5825, A2 => DATA1(2), ZN => n6054);
   U1309 : NAND2_X1 port map( A1 => n6044, A2 => DATA1(1), ZN => n6544);
   U1310 : OAI211_X1 port map( C1 => n6112, C2 => n6696, A => n6054, B => n6544
                           , ZN => n6052);
   U1311 : AOI211_X1 port map( C1 => n6388, C2 => n6389, A => n6865, B => n6648
                           , ZN => n6051);
   U1312 : OAI22_X1 port map( A1 => n6865, A2 => DATA1(2), B1 => n6648, B2 => 
                           DATA2(2), ZN => n6814);
   U1313 : INV_X1 port map( A => n6814, ZN => n6703);
   U1314 : AOI22_X1 port map( A1 => n6047, A2 => n6046, B1 => n6632, B2 => 
                           n6045, ZN => n6049);
   U1315 : OAI22_X1 port map( A1 => n6703, A2 => n6492, B1 => n6049, B2 => 
                           n6048, ZN => n6050);
   U1316 : AOI211_X1 port map( C1 => n6527, C2 => n6052, A => n6051, B => n6050
                           , ZN => n6093);
   U1317 : OAI22_X1 port map( A1 => n6621, A2 => n6139, B1 => n6623, B2 => 
                           n6618, ZN => n6091);
   U1318 : INV_X1 port map( A => n6303, ZN => n6572);
   U1319 : OAI211_X1 port map( C1 => n6055, C2 => n6695, A => n6054, B => n6053
                           , ZN => n6056);
   U1320 : AOI211_X1 port map( C1 => n6059, C2 => n6058, A => n6057, B => n6056
                           , ZN => n6290);
   U1321 : OAI222_X1 port map( A1 => n6064, A2 => n6290, B1 => n6063, B2 => 
                           n6062, C1 => n6061, C2 => n6060, ZN => n6553);
   U1322 : AOI22_X1 port map( A1 => n6232, A2 => n6065, B1 => n6228, B2 => 
                           n6553, ZN => n6070);
   U1323 : AOI22_X1 port map( A1 => n6565, A2 => n6068, B1 => n6067, B2 => 
                           n6066, ZN => n6069);
   U1324 : OAI211_X1 port map( C1 => n6293, C2 => n6558, A => n6070, B => n6069
                           , ZN => n6284);
   U1325 : AOI22_X1 port map( A1 => n6577, A2 => n6301, B1 => n6526, B2 => 
                           n6284, ZN => n6075);
   U1326 : AOI22_X1 port map( A1 => n6073, A2 => n6576, B1 => n6072, B2 => 
                           n6071, ZN => n6074);
   U1327 : OAI211_X1 port map( C1 => n6572, C2 => n6451, A => n6075, B => n6074
                           , ZN => n6580);
   U1328 : AOI222_X1 port map( A1 => n6076, A2 => n6579, B1 => n6306, B2 => 
                           n6584, C1 => n6580, C2 => n6582, ZN => n6585);
   U1329 : OAI22_X1 port map( A1 => n6589, A2 => n6586, B1 => n6585, B2 => 
                           n6307, ZN => n6079);
   U1330 : OAI22_X1 port map( A1 => n6590, A2 => n6077, B1 => n6309, B2 => 
                           n6310, ZN => n6078);
   U1331 : AOI211_X1 port map( C1 => n6475, C2 => n6596, A => n6079, B => n6078
                           , ZN => n6599);
   U1332 : OAI22_X1 port map( A1 => n6598, A2 => n6599, B1 => n6080, B2 => 
                           n6600, ZN => n6086);
   U1333 : OAI22_X1 port map( A1 => n6084, A2 => n6083, B1 => n6082, B2 => 
                           n6081, ZN => n6085);
   U1334 : AOI211_X1 port map( C1 => n6518, C2 => n6602, A => n6086, B => n6085
                           , ZN => n6087);
   U1335 : INV_X1 port map( A => n6087, ZN => n6614);
   U1336 : AOI222_X1 port map( A1 => n6321, A2 => n6614, B1 => n6320, B2 => 
                           n6089, C1 => n6088, C2 => n6615, ZN => n6619);
   U1337 : OAI22_X1 port map( A1 => n6619, A2 => n6616, B1 => n6322, B2 => 
                           n6620, ZN => n6090);
   U1338 : OAI21_X1 port map( B1 => n6091, B2 => n6090, A => n6510, ZN => n6092
                           );
   U1339 : NAND3_X1 port map( A1 => n6094, A2 => n6093, A3 => n6092, ZN => 
                           OUTALU(2));
   U1340 : AOI22_X1 port map( A1 => n6173, A2 => n6120, B1 => n6186, B2 => 
                           n6119, ZN => n6110);
   U1341 : INV_X1 port map( A => DATA2(29), ZN => n6836);
   U1342 : AOI221_X1 port map( B1 => n6149, B2 => n6114, C1 => n6836, C2 => 
                           n6114, A => n6095, ZN => n6100);
   U1343 : NOR2_X1 port map( A1 => DATA2(29), A2 => n6095, ZN => n6770);
   U1344 : NOR2_X1 port map( A1 => DATA1(29), A2 => n6836, ZN => n6766);
   U1345 : NOR2_X1 port map( A1 => n6770, A2 => n6766, ZN => n6788);
   U1346 : AOI21_X1 port map( B1 => DATA1(31), B2 => n6097, A => n6096, ZN => 
                           n6098);
   U1347 : OAI22_X1 port map( A1 => n6788, A2 => n6492, B1 => n6098, B2 => 
                           n6830, ZN => n6099);
   U1348 : AOI211_X1 port map( C1 => dataout_mul_29_port, C2 => n6501, A => 
                           n6100, B => n6099, ZN => n6109);
   U1349 : OAI22_X1 port map( A1 => n6140, A2 => n6618, B1 => n6101, B2 => 
                           n6616, ZN => n6107);
   U1350 : OAI22_X1 port map( A1 => n6118, A2 => n6139, B1 => n6158, B2 => 
                           n6620, ZN => n6106);
   U1351 : INV_X1 port map( A => n6111, ZN => n6103);
   U1352 : AOI21_X1 port map( B1 => n6104, B2 => n6103, A => n6102, ZN => n6105
                           );
   U1353 : AOI221_X1 port map( B1 => n6107, B2 => n6527, C1 => n6106, C2 => 
                           n6527, A => n6105, ZN => n6108);
   U1354 : OAI211_X1 port map( C1 => n6111, C2 => n6110, A => n6109, B => n6108
                           , ZN => OUTALU(29));
   U1355 : INV_X1 port map( A => DATA2(28), ZN => n6837);
   U1356 : AOI22_X1 port map( A1 => DATA1(28), A2 => DATA2(28), B1 => n6837, B2
                           => n6768, ZN => n6810);
   U1357 : AOI22_X1 port map( A1 => dataout_mul_28_port, A2 => n6501, B1 => 
                           n6631, B2 => n6810, ZN => n6131);
   U1358 : OAI22_X1 port map( A1 => n6113, A2 => n6689, B1 => n6112, B2 => 
                           n6686, ZN => n6116);
   U1359 : AOI221_X1 port map( B1 => n6149, B2 => n6114, C1 => n6837, C2 => 
                           n6114, A => n6768, ZN => n6115);
   U1360 : AOI221_X1 port map( B1 => n6117, B2 => n6510, C1 => n6116, C2 => 
                           n6510, A => n6115, ZN => n6130);
   U1361 : OAI222_X1 port map( A1 => n6139, A2 => n6140, B1 => n6618, B2 => 
                           n6158, C1 => n6616, C2 => n6118, ZN => n6124);
   U1362 : OAI22_X1 port map( A1 => n6120, A2 => n6194, B1 => n6119, B2 => 
                           n6125, ZN => n6123);
   U1363 : NAND2_X1 port map( A1 => n6121, A2 => n6126, ZN => n6122);
   U1364 : AOI22_X1 port map( A1 => n6527, A2 => n6124, B1 => n6123, B2 => 
                           n6122, ZN => n6129);
   U1365 : INV_X1 port map( A => n6145, ZN => n6127);
   U1366 : OAI22_X1 port map( A1 => n6133, A2 => n6194, B1 => n6132, B2 => 
                           n6125, ZN => n6141);
   U1367 : NAND3_X1 port map( A1 => n6127, A2 => n6126, A3 => n6141, ZN => 
                           n6128);
   U1368 : NAND4_X1 port map( A1 => n6131, A2 => n6130, A3 => n6129, A4 => 
                           n6128, ZN => OUTALU(28));
   U1369 : AOI22_X1 port map( A1 => n6173, A2 => n6133, B1 => n6186, B2 => 
                           n6132, ZN => n6146);
   U1370 : AOI21_X1 port map( B1 => n6633, B2 => DATA2(27), A => n6493, ZN => 
                           n6137);
   U1371 : NOR2_X1 port map( A1 => DATA2(27), A2 => n6136, ZN => n6764);
   U1372 : INV_X1 port map( A => DATA2(27), ZN => n6838);
   U1373 : NOR2_X1 port map( A1 => DATA1(27), A2 => n6838, ZN => n6762);
   U1374 : OAI21_X1 port map( B1 => n6764, B2 => n6762, A => n6631, ZN => n6135
                           );
   U1375 : NAND3_X1 port map( A1 => n6510, A2 => n6152, A3 => n6150, ZN => 
                           n6134);
   U1376 : OAI211_X1 port map( C1 => n6137, C2 => n6136, A => n6135, B => n6134
                           , ZN => n6138);
   U1377 : AOI21_X1 port map( B1 => n6641, B2 => dataout_mul_27_port, A => 
                           n6138, ZN => n6144);
   U1378 : OAI22_X1 port map( A1 => n6140, A2 => n6616, B1 => n6158, B2 => 
                           n6139, ZN => n6142);
   U1379 : AOI22_X1 port map( A1 => n6527, A2 => n6142, B1 => n6145, B2 => 
                           n6141, ZN => n6143);
   U1380 : OAI211_X1 port map( C1 => n6146, C2 => n6145, A => n6144, B => n6143
                           , ZN => OUTALU(27));
   U1381 : AOI22_X1 port map( A1 => n6173, A2 => n6148, B1 => n6186, B2 => 
                           n6147, ZN => n6163);
   U1382 : INV_X1 port map( A => DATA2(26), ZN => n6839);
   U1383 : NOR3_X1 port map( A1 => n6149, A2 => n6839, A3 => n6763, ZN => n6155
                           );
   U1384 : AOI22_X1 port map( A1 => DATA1(26), A2 => n6839, B1 => DATA2(26), B2
                           => n6763, ZN => n6758);
   U1385 : AOI22_X1 port map( A1 => n6152, A2 => n6151, B1 => n6547, B2 => 
                           n6150, ZN => n6153);
   U1386 : OAI22_X1 port map( A1 => n6758, A2 => n6531, B1 => n6153, B2 => 
                           n6830, ZN => n6154);
   U1387 : AOI211_X1 port map( C1 => dataout_mul_26_port, C2 => n6501, A => 
                           n6155, B => n6154, ZN => n6162);
   U1388 : AOI22_X1 port map( A1 => n6173, A2 => n6172, B1 => n6186, B2 => 
                           n6167, ZN => n6156);
   U1389 : INV_X1 port map( A => n6156, ZN => n6175);
   U1390 : AND2_X1 port map( A1 => n6157, A2 => n6175, ZN => n6160);
   U1391 : NOR3_X1 port map( A1 => n6158, A2 => n6496, A3 => n6616, ZN => n6159
                           );
   U1392 : AOI21_X1 port map( B1 => n6160, B2 => n6164, A => n6159, ZN => n6161
                           );
   U1393 : OAI211_X1 port map( C1 => n6164, C2 => n6163, A => n6162, B => n6161
                           , ZN => OUTALU(26));
   U1394 : AOI22_X1 port map( A1 => n6612, A2 => n6191, B1 => n6610, B2 => 
                           n6165, ZN => n6179);
   U1395 : NOR3_X1 port map( A1 => n6292, A2 => n6196, A3 => n6830, ZN => n6171
                           );
   U1396 : INV_X1 port map( A => DATA2(25), ZN => n6840);
   U1397 : NAND2_X1 port map( A1 => DATA1(25), A2 => n6840, ZN => n6759);
   U1398 : NAND2_X1 port map( A1 => DATA2(25), A2 => n6166, ZN => n6690);
   U1399 : AND2_X1 port map( A1 => n6759, A2 => n6690, ZN => n6778);
   U1400 : NAND3_X1 port map( A1 => DATA2(25), A2 => DATA1(25), A3 => n6528, ZN
                           => n6169);
   U1401 : NAND4_X1 port map( A1 => DATA2_I_24_port, A2 => DATA1(24), A3 => 
                           n6186, A4 => n6167, ZN => n6168);
   U1402 : OAI211_X1 port map( C1 => n6778, C2 => n6531, A => n6169, B => n6168
                           , ZN => n6170);
   U1403 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_25_port, A => 
                           n6171, B => n6170, ZN => n6178);
   U1404 : AND2_X1 port map( A1 => n6173, A2 => n6172, ZN => n6174);
   U1405 : AOI22_X1 port map( A1 => n6176, A2 => n6175, B1 => n6174, B2 => 
                           n6195, ZN => n6177);
   U1406 : OAI211_X1 port map( C1 => n6179, C2 => n6496, A => n6178, B => n6177
                           , ZN => OUTALU(25));
   U1407 : INV_X1 port map( A => DATA2(24), ZN => n6841);
   U1408 : OAI22_X1 port map( A1 => n6841, A2 => n6389, B1 => n6194, B2 => 
                           n6180, ZN => n6190);
   U1409 : OAI22_X1 port map( A1 => n6680, A2 => DATA2(24), B1 => n6841, B2 => 
                           n6691, ZN => n6811);
   U1410 : INV_X1 port map( A => n6811, ZN => n6755);
   U1411 : OAI22_X1 port map( A1 => n6292, A2 => n6182, B1 => n6196, B2 => 
                           n6181, ZN => n6184);
   U1412 : AOI22_X1 port map( A1 => n6510, A2 => n6184, B1 => n6183, B2 => 
                           dataout_mul_24_port, ZN => n6188);
   U1413 : NAND2_X1 port map( A1 => n6691, A2 => DATA2_I_24_port, ZN => n6185);
   U1414 : NAND3_X1 port map( A1 => n6186, A2 => n6195, A3 => n6185, ZN => 
                           n6187);
   U1415 : OAI211_X1 port map( C1 => n6755, C2 => n6492, A => n6188, B => n6187
                           , ZN => n6189);
   U1416 : AOI221_X1 port map( B1 => n6493, B2 => DATA1(24), C1 => n6190, C2 =>
                           DATA1(24), A => n6189, ZN => n6193);
   U1417 : NAND3_X1 port map( A1 => n6527, A2 => n6321, A3 => n6191, ZN => 
                           n6192);
   U1418 : OAI211_X1 port map( C1 => n6195, C2 => n6194, A => n6193, B => n6192
                           , ZN => OUTALU(24));
   U1419 : INV_X1 port map( A => n6196, ZN => n6233);
   U1420 : AOI222_X1 port map( A1 => n6229, A2 => n6197, B1 => n6233, B2 => 
                           n6232, C1 => n6231, C2 => n6230, ZN => n6226);
   U1421 : INV_X1 port map( A => DATA2(23), ZN => n6842);
   U1422 : NAND2_X1 port map( A1 => DATA1(23), A2 => n6842, ZN => n6754);
   U1423 : NAND2_X1 port map( A1 => DATA2(23), A2 => n6198, ZN => n6752);
   U1424 : AOI21_X1 port map( B1 => n6754, B2 => n6752, A => n6531, ZN => n6200
                           );
   U1425 : AOI211_X1 port map( C1 => n6388, C2 => n6389, A => n6198, B => n6842
                           , ZN => n6199);
   U1426 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_23_port, A => 
                           n6200, B => n6199, ZN => n6225);
   U1427 : NAND2_X1 port map( A1 => n6833, A2 => n6210, ZN => n6401);
   U1428 : AND2_X1 port map( A1 => DATA1(17), A2 => DATA2_I_17_port, ZN => 
                           n6202);
   U1429 : NOR2_X1 port map( A1 => n6202, A2 => n6201, ZN => n6354);
   U1430 : OAI21_X1 port map( B1 => n6367, B2 => n6354, A => n6203, ZN => n6334
                           );
   U1431 : INV_X1 port map( A => n6204, ZN => n6205);
   U1432 : AOI21_X1 port map( B1 => n6206, B2 => n6334, A => n6205, ZN => n6265
                           );
   U1433 : OAI21_X1 port map( B1 => n6267, B2 => n6265, A => n6207, ZN => n6252
                           );
   U1434 : INV_X1 port map( A => n6252, ZN => n6209);
   U1435 : NAND2_X1 port map( A1 => DATA1(21), A2 => DATA2_I_21_port, ZN => 
                           n6208);
   U1436 : OAI21_X1 port map( B1 => n6209, B2 => n6255, A => n6208, ZN => n6216
                           );
   U1437 : NOR2_X1 port map( A1 => n7166, A2 => n6210, ZN => n6352);
   U1438 : AOI21_X1 port map( B1 => n6214, B2 => n6352, A => n6234, ZN => n6211
                           );
   U1439 : OAI21_X1 port map( B1 => n6401, B2 => n6216, A => n6211, ZN => n6243
                           );
   U1440 : NAND3_X1 port map( A1 => n6243, A2 => n6217, A3 => n6213, ZN => 
                           n6212);
   U1441 : OAI21_X1 port map( B1 => n6217, B2 => n6213, A => n6212, ZN => n6223
                           );
   U1442 : INV_X1 port map( A => n6401, ZN => n6351);
   U1443 : INV_X1 port map( A => n6214, ZN => n6215);
   U1444 : AOI22_X1 port map( A1 => n6351, A2 => n6216, B1 => n6352, B2 => 
                           n6215, ZN => n6235);
   U1445 : NOR3_X1 port map( A1 => n6217, A2 => n6235, A3 => n6234, ZN => n6222
                           );
   U1446 : AOI22_X1 port map( A1 => n6315, A2 => n6247, B1 => n6516, B2 => 
                           n6218, ZN => n6220);
   U1447 : AOI22_X1 port map( A1 => n6603, A2 => n6271, B1 => n6518, B2 => 
                           n6237, ZN => n6219);
   U1448 : AOI21_X1 port map( B1 => n6220, B2 => n6219, A => n6496, ZN => n6221
                           );
   U1449 : AOI211_X1 port map( C1 => n6833, C2 => n6223, A => n6222, B => n6221
                           , ZN => n6224);
   U1450 : OAI211_X1 port map( C1 => n6226, C2 => n6830, A => n6225, B => n6224
                           , ZN => OUTALU(23));
   U1451 : AOI22_X1 port map( A1 => n6230, A2 => n6229, B1 => n6228, B2 => 
                           n6227, ZN => n6246);
   U1452 : AOI22_X1 port map( A1 => n6565, A2 => n6233, B1 => n6232, B2 => 
                           n6231, ZN => n6245);
   U1453 : NAND2_X1 port map( A1 => n6235, A2 => n6234, ZN => n6242);
   U1454 : AOI222_X1 port map( A1 => n6237, A2 => n6509, B1 => n6247, B2 => 
                           n6518, C1 => n6271, C2 => n6236, ZN => n6240);
   U1455 : INV_X1 port map( A => DATA2(22), ZN => n6843);
   U1456 : AOI22_X1 port map( A1 => DATA1(22), A2 => DATA2(22), B1 => n6843, B2
                           => n6677, ZN => n6748);
   U1457 : AOI22_X1 port map( A1 => dataout_mul_22_port, A2 => n6501, B1 => 
                           n6631, B2 => n6748, ZN => n6239);
   U1458 : NAND3_X1 port map( A1 => DATA2(22), A2 => n6753, A3 => n6528, ZN => 
                           n6238);
   U1459 : OAI211_X1 port map( C1 => n6240, C2 => n6496, A => n6239, B => n6238
                           , ZN => n6241);
   U1460 : AOI21_X1 port map( B1 => n6243, B2 => n6242, A => n6241, ZN => n6244
                           );
   U1461 : OAI221_X1 port map( B1 => n6830, B2 => n6246, C1 => n6830, C2 => 
                           n6245, A => n6244, ZN => OUTALU(22));
   U1462 : AOI22_X1 port map( A1 => n6518, A2 => n6271, B1 => n6516, B2 => 
                           n6247, ZN => n6261);
   U1463 : NOR3_X1 port map( A1 => n6359, A2 => n6830, A3 => n6566, ZN => n6251
                           );
   U1464 : NOR2_X1 port map( A1 => DATA2(21), A2 => n6248, ZN => n6749);
   U1465 : NAND2_X1 port map( A1 => n6248, A2 => DATA2(21), ZN => n6750);
   U1466 : INV_X1 port map( A => n6750, ZN => n6675);
   U1467 : NOR2_X1 port map( A1 => n6749, A2 => n6675, ZN => n6786);
   U1468 : AOI21_X1 port map( B1 => n6633, B2 => DATA2(21), A => n6493, ZN => 
                           n6249);
   U1469 : OAI22_X1 port map( A1 => n6786, A2 => n6492, B1 => n6249, B2 => 
                           n6248, ZN => n6250);
   U1470 : AOI211_X1 port map( C1 => dataout_mul_21_port, C2 => n6501, A => 
                           n6251, B => n6250, ZN => n6260);
   U1471 : INV_X1 port map( A => n6352, ZN => n6399);
   U1472 : OAI22_X1 port map( A1 => n6253, A2 => n6399, B1 => n6401, B2 => 
                           n6252, ZN => n6257);
   U1473 : AOI22_X1 port map( A1 => n6253, A2 => n6352, B1 => n6252, B2 => 
                           n6351, ZN => n6254);
   U1474 : INV_X1 port map( A => n6254, ZN => n6256);
   U1475 : AOI22_X1 port map( A1 => n6258, A2 => n6257, B1 => n6256, B2 => 
                           n6255, ZN => n6259);
   U1476 : OAI211_X1 port map( C1 => n6261, C2 => n6496, A => n6260, B => n6259
                           , ZN => OUTALU(21));
   U1477 : OAI22_X1 port map( A1 => n6360, A2 => n5224, B1 => n6359, B2 => 
                           n6570, ZN => n6262);
   U1478 : AOI22_X1 port map( A1 => n6510, A2 => n6262, B1 => n6641, B2 => 
                           dataout_mul_20_port, ZN => n6275);
   U1479 : INV_X1 port map( A => DATA2(20), ZN => n6845);
   U1480 : OAI21_X1 port map( B1 => n6389, B2 => n6845, A => n6388, ZN => n6263
                           );
   U1481 : NAND2_X1 port map( A1 => DATA1(20), A2 => n6845, ZN => n6673);
   U1482 : OAI21_X1 port map( B1 => DATA1(20), B2 => n6845, A => n6673, ZN => 
                           n6642);
   U1483 : AOI22_X1 port map( A1 => DATA1(20), A2 => n6263, B1 => n6631, B2 => 
                           n6642, ZN => n6274);
   U1484 : INV_X1 port map( A => n6267, ZN => n6270);
   U1485 : AOI22_X1 port map( A1 => n6266, A2 => n6352, B1 => n6351, B2 => 
                           n6265, ZN => n6264);
   U1486 : INV_X1 port map( A => n6264, ZN => n6269);
   U1487 : OAI22_X1 port map( A1 => n6266, A2 => n6399, B1 => n6265, B2 => 
                           n6401, ZN => n6268);
   U1488 : AOI22_X1 port map( A1 => n6270, A2 => n6269, B1 => n6268, B2 => 
                           n6267, ZN => n6273);
   U1489 : NAND3_X1 port map( A1 => n6527, A2 => n6509, A3 => n6271, ZN => 
                           n6272);
   U1490 : NAND4_X1 port map( A1 => n6275, A2 => n6274, A3 => n6273, A4 => 
                           n6272, ZN => OUTALU(20));
   U1491 : NOR2_X1 port map( A1 => n6327, A2 => DATA2(1), ZN => n6699);
   U1492 : NAND2_X1 port map( A1 => n6327, A2 => DATA2(1), ZN => n6697);
   U1493 : INV_X1 port map( A => n6697, ZN => n6647);
   U1494 : NOR2_X1 port map( A1 => n6699, A2 => n6647, ZN => n6779);
   U1495 : AOI21_X1 port map( B1 => n6277, B2 => n6278, A => n6276, ZN => n6282
                           );
   U1496 : AOI221_X1 port map( B1 => n6280, B2 => n6279, C1 => n6630, C2 => 
                           n6278, A => n6637, ZN => n6281);
   U1497 : AOI21_X1 port map( B1 => n6282, B2 => n6632, A => n6281, ZN => n6332
                           );
   U1498 : NOR3_X1 port map( A1 => n6283, A2 => n6696, A3 => n6496, ZN => n6330
                           );
   U1499 : INV_X1 port map( A => n6619, ZN => n6325);
   U1500 : INV_X1 port map( A => n6585, ZN => n6313);
   U1501 : INV_X1 port map( A => n6284, ZN => n6569);
   U1502 : OAI211_X1 port map( C1 => n6326, C2 => n6327, A => n6286, B => n6285
                           , ZN => n6287);
   U1503 : AOI211_X1 port map( C1 => DATA1(4), C2 => n6542, A => n6288, B => 
                           n6287, ZN => n6289);
   U1504 : INV_X1 port map( A => n6289, ZN => n6548);
   U1505 : INV_X1 port map( A => n6290, ZN => n6552);
   U1506 : AOI222_X1 port map( A1 => n6549, A2 => n6548, B1 => n6547, B2 => 
                           n6552, C1 => n6551, C2 => n6291, ZN => n6559);
   U1507 : OAI22_X1 port map( A1 => n6554, A2 => n6293, B1 => n6292, B2 => 
                           n6559, ZN => n6297);
   U1508 : OAI22_X1 port map( A1 => n6295, A2 => n6560, B1 => n6561, B2 => 
                           n6294, ZN => n6296);
   U1509 : AOI211_X1 port map( C1 => n6553, C2 => n6298, A => n6297, B => n6296
                           , ZN => n6571);
   U1510 : OAI22_X1 port map( A1 => n6451, A2 => n6299, B1 => n6566, B2 => 
                           n6571, ZN => n6300);
   U1511 : INV_X1 port map( A => n6300, ZN => n6305);
   U1512 : AOI22_X1 port map( A1 => n6577, A2 => n6303, B1 => n6302, B2 => 
                           n6301, ZN => n6304);
   U1513 : OAI211_X1 port map( C1 => n6569, C2 => n6570, A => n6305, B => n6304
                           , ZN => n6583);
   U1514 : AOI222_X1 port map( A1 => n6306, A2 => n6579, B1 => n6580, B2 => 
                           n6584, C1 => n6583, C2 => n6582, ZN => n6591);
   U1515 : OAI22_X1 port map( A1 => n6308, A2 => n6586, B1 => n6591, B2 => 
                           n6307, ZN => n6312);
   U1516 : OAI22_X1 port map( A1 => n6589, A2 => n6310, B1 => n6590, B2 => 
                           n6309, ZN => n6311);
   U1517 : AOI211_X1 port map( C1 => n6475, C2 => n6313, A => n6312, B => n6311
                           , ZN => n6609);
   U1518 : INV_X1 port map( A => n6609, ZN => n6314);
   U1519 : AOI22_X1 port map( A1 => n6602, A2 => n6315, B1 => n6516, B2 => 
                           n6314, ZN => n6319);
   U1520 : AOI22_X1 port map( A1 => n6317, A2 => n6316, B1 => n6604, B2 => 
                           n6603, ZN => n6318);
   U1521 : OAI211_X1 port map( C1 => n6608, C2 => n6599, A => n6319, B => n6318
                           , ZN => n6613);
   U1522 : AOI222_X1 port map( A1 => n6612, A2 => n6614, B1 => n6321, B2 => 
                           n6613, C1 => n6320, C2 => n6615, ZN => n6541);
   U1523 : OAI22_X1 port map( A1 => n6541, A2 => n6616, B1 => n6623, B2 => 
                           n6620, ZN => n6324);
   U1524 : OAI22_X1 port map( A1 => n6621, A2 => n6618, B1 => n6322, B2 => 
                           n6622, ZN => n6323);
   U1525 : AOI211_X1 port map( C1 => n6627, C2 => n6325, A => n6324, B => n6323
                           , ZN => n6629);
   U1526 : OAI21_X1 port map( B1 => n6496, B2 => n6326, A => n6388, ZN => n6634
                           );
   U1527 : AOI21_X1 port map( B1 => DATA2(1), B2 => n6633, A => n6634, ZN => 
                           n6328);
   U1528 : OAI22_X1 port map( A1 => n6629, A2 => n6830, B1 => n6328, B2 => 
                           n6327, ZN => n6329);
   U1529 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_1_port, A => 
                           n6330, B => n6329, ZN => n6331);
   U1530 : OAI211_X1 port map( C1 => n6779, C2 => n6492, A => n6332, B => n6331
                           , ZN => OUTALU(1));
   U1531 : AOI22_X1 port map( A1 => n6472, A2 => n6333, B1 => n6475, B2 => 
                           n6350, ZN => n6349);
   U1532 : AOI22_X1 port map( A1 => n6595, A2 => n6390, B1 => n6470, B2 => 
                           n6372, ZN => n6348);
   U1533 : INV_X1 port map( A => n6344, ZN => n6346);
   U1534 : OAI22_X1 port map( A1 => n6335, A2 => n6399, B1 => n6401, B2 => 
                           n6334, ZN => n6345);
   U1535 : AOI22_X1 port map( A1 => n6335, A2 => n6352, B1 => n6334, B2 => 
                           n6351, ZN => n6336);
   U1536 : INV_X1 port map( A => n6336, ZN => n6343);
   U1537 : AOI21_X1 port map( B1 => n6633, B2 => DATA2(19), A => n6493, ZN => 
                           n6341);
   U1538 : OAI222_X1 port map( A1 => n6570, A2 => n6360, B1 => n6566, B2 => 
                           n6357, C1 => n6451, C2 => n6359, ZN => n6337);
   U1539 : AOI22_X1 port map( A1 => n6510, A2 => n6337, B1 => n6501, B2 => 
                           dataout_mul_19_port, ZN => n6339);
   U1540 : INV_X1 port map( A => DATA2(19), ZN => n6846);
   U1541 : NOR2_X1 port map( A1 => DATA1(19), A2 => n6846, ZN => n6742);
   U1542 : NOR2_X1 port map( A1 => n6340, A2 => DATA2(19), ZN => n6806);
   U1543 : OAI21_X1 port map( B1 => n6742, B2 => n6806, A => n6631, ZN => n6338
                           );
   U1544 : OAI211_X1 port map( C1 => n6341, C2 => n6340, A => n6339, B => n6338
                           , ZN => n6342);
   U1545 : AOI221_X1 port map( B1 => n6346, B2 => n6345, C1 => n6344, C2 => 
                           n6343, A => n6342, ZN => n6347);
   U1546 : OAI221_X1 port map( B1 => n6496, B2 => n6349, C1 => n6496, C2 => 
                           n6348, A => n6347, ZN => OUTALU(19));
   U1547 : AOI222_X1 port map( A1 => n6350, A2 => n6472, B1 => n6372, B2 => 
                           n6475, C1 => n6390, C2 => n6470, ZN => n6371);
   U1548 : INV_X1 port map( A => n6367, ZN => n6369);
   U1549 : AOI22_X1 port map( A1 => n6355, A2 => n6352, B1 => n6351, B2 => 
                           n6354, ZN => n6353);
   U1550 : INV_X1 port map( A => n6353, ZN => n6368);
   U1551 : OAI22_X1 port map( A1 => n6355, A2 => n6399, B1 => n6354, B2 => 
                           n6401, ZN => n6366);
   U1552 : INV_X1 port map( A => DATA2(18), ZN => n6847);
   U1553 : NOR2_X1 port map( A1 => DATA1(18), A2 => n6847, ZN => n6741);
   U1554 : NAND2_X1 port map( A1 => DATA1(18), A2 => n6847, ZN => n6670);
   U1555 : INV_X1 port map( A => n6670, ZN => n6736);
   U1556 : NOR2_X1 port map( A1 => n6741, A2 => n6736, ZN => n6795);
   U1557 : OAI21_X1 port map( B1 => n6389, B2 => n6847, A => n6388, ZN => n6356
                           );
   U1558 : AOI22_X1 port map( A1 => DATA1(18), A2 => n6356, B1 => n6501, B2 => 
                           dataout_mul_18_port, ZN => n6364);
   U1559 : OAI22_X1 port map( A1 => n6358, A2 => n5224, B1 => n6357, B2 => 
                           n6570, ZN => n6362);
   U1560 : OAI22_X1 port map( A1 => n6360, A2 => n6451, B1 => n6359, B2 => 
                           n6450, ZN => n6361);
   U1561 : OAI21_X1 port map( B1 => n6362, B2 => n6361, A => n6510, ZN => n6363
                           );
   U1562 : OAI211_X1 port map( C1 => n6795, C2 => n6531, A => n6364, B => n6363
                           , ZN => n6365);
   U1563 : AOI221_X1 port map( B1 => n6369, B2 => n6368, C1 => n6367, C2 => 
                           n6366, A => n6365, ZN => n6370);
   U1564 : OAI21_X1 port map( B1 => n6371, B2 => n6496, A => n6370, ZN => 
                           OUTALU(18));
   U1565 : AOI22_X1 port map( A1 => n6472, A2 => n6372, B1 => n6475, B2 => 
                           n6390, ZN => n6385);
   U1566 : INV_X1 port map( A => n6374, ZN => n6386);
   U1567 : OAI22_X1 port map( A1 => n6373, A2 => n6399, B1 => n6401, B2 => 
                           n6386, ZN => n6382);
   U1568 : OAI22_X1 port map( A1 => n6374, A2 => n6401, B1 => n6387, B2 => 
                           n6399, ZN => n6380);
   U1569 : NOR2_X1 port map( A1 => DATA2(17), A2 => n6375, ZN => n6737);
   U1570 : INV_X1 port map( A => DATA2(17), ZN => n6848);
   U1571 : NOR2_X1 port map( A1 => n6848, A2 => DATA1(17), ZN => n6643);
   U1572 : NOR2_X1 port map( A1 => n6737, A2 => n6643, ZN => n6777);
   U1573 : NOR3_X1 port map( A1 => n6391, A2 => n6830, A3 => n6410, ZN => n6376
                           );
   U1574 : AOI21_X1 port map( B1 => dataout_mul_17_port, B2 => n6501, A => 
                           n6376, ZN => n6378);
   U1575 : NAND3_X1 port map( A1 => DATA2(17), A2 => DATA1(17), A3 => n6528, ZN
                           => n6377);
   U1576 : OAI211_X1 port map( C1 => n6777, C2 => n6492, A => n6378, B => n6377
                           , ZN => n6379);
   U1577 : AOI221_X1 port map( B1 => n6383, B2 => n6382, C1 => n6381, C2 => 
                           n6380, A => n6379, ZN => n6384);
   U1578 : OAI21_X1 port map( B1 => n6385, B2 => n6496, A => n6384, ZN => 
                           OUTALU(17));
   U1579 : NAND2_X1 port map( A1 => n6387, A2 => n6386, ZN => n6400);
   U1580 : INV_X1 port map( A => n6400, ZN => n6402);
   U1581 : INV_X1 port map( A => DATA2(16), ZN => n6849);
   U1582 : OAI21_X1 port map( B1 => n6389, B2 => n6849, A => n6388, ZN => n6397
                           );
   U1583 : AND3_X1 port map( A1 => n6390, A2 => n6527, A3 => n6472, ZN => n6396
                           );
   U1584 : NOR2_X1 port map( A1 => DATA2(16), A2 => n6735, ZN => n6731);
   U1585 : AOI21_X1 port map( B1 => DATA2(16), B2 => n6735, A => n6731, ZN => 
                           n6667);
   U1586 : OAI22_X1 port map( A1 => n6392, A2 => n6410, B1 => n6391, B2 => 
                           n6409, ZN => n6393);
   U1587 : AOI22_X1 port map( A1 => n6510, A2 => n6393, B1 => n6641, B2 => 
                           dataout_mul_16_port, ZN => n6394);
   U1588 : OAI21_X1 port map( B1 => n6667, B2 => n6531, A => n6394, ZN => n6395
                           );
   U1589 : AOI211_X1 port map( C1 => DATA1(16), C2 => n6397, A => n6396, B => 
                           n6395, ZN => n6398);
   U1590 : OAI221_X1 port map( B1 => n6402, B2 => n6401, C1 => n6400, C2 => 
                           n6399, A => n6398, ZN => OUTALU(16));
   U1591 : NAND2_X1 port map( A1 => DATA2(15), A2 => n6403, ZN => n6732);
   U1592 : INV_X1 port map( A => DATA2(15), ZN => n6850);
   U1593 : NAND2_X1 port map( A1 => n6850, A2 => DATA1(15), ZN => n6644);
   U1594 : AOI21_X1 port map( B1 => n6732, B2 => n6644, A => n6492, ZN => n6408
                           );
   U1595 : INV_X1 port map( A => n6405, ZN => n6419);
   U1596 : INV_X1 port map( A => n6404, ZN => n6406);
   U1597 : INV_X1 port map( A => n6504, ZN => n6521);
   U1598 : AOI221_X1 port map( B1 => n6419, B2 => n6406, C1 => n6405, C2 => 
                           n6404, A => n6521, ZN => n6407);
   U1599 : AOI211_X1 port map( C1 => dataout_mul_15_port, C2 => n6501, A => 
                           n6408, B => n6407, ZN => n6426);
   U1600 : OAI22_X1 port map( A1 => n6411, A2 => n6410, B1 => n6431, B2 => 
                           n6409, ZN => n6422);
   U1601 : INV_X1 port map( A => n6519, ZN => n6413);
   U1602 : INV_X1 port map( A => n6520, ZN => n6412);
   U1603 : OAI21_X1 port map( B1 => n6413, B2 => n6537, A => n6412, ZN => n6534
                           );
   U1604 : NAND2_X1 port map( A1 => n6414, A2 => n6534, ZN => n6503);
   U1605 : INV_X1 port map( A => n6503, ZN => n6502);
   U1606 : OAI21_X1 port map( B1 => n6416, B2 => n6502, A => n6415, ZN => n6486
                           );
   U1607 : AOI21_X1 port map( B1 => n6418, B2 => n6486, A => n6417, ZN => n6436
                           );
   U1608 : NAND2_X1 port map( A1 => n6436, A2 => n6435, ZN => n6433);
   U1609 : AOI22_X1 port map( A1 => DATA1(14), A2 => DATA2_I_14_port, B1 => 
                           n6439, B2 => n6433, ZN => n6420);
   U1610 : XNOR2_X1 port map( A => n6420, B => n6419, ZN => n6421);
   U1611 : AOI22_X1 port map( A1 => n6527, A2 => n6422, B1 => n6535, B2 => 
                           n6421, ZN => n6425);
   U1612 : NAND3_X1 port map( A1 => n6510, A2 => n6472, A3 => n6473, ZN => 
                           n6424);
   U1613 : NAND3_X1 port map( A1 => DATA2(15), A2 => DATA1(15), A3 => n6528, ZN
                           => n6423);
   U1614 : NAND4_X1 port map( A1 => n6426, A2 => n6425, A3 => n6424, A4 => 
                           n6423, ZN => OUTALU(15));
   U1615 : NAND2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           ZN => n7096);
   U1616 : OAI21_X1 port map( B1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, B2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           A => n7096, ZN => n7098);
   U1617 : NOR3_X1 port map( A1 => n5126, A2 => n5134, A3 => n7098, ZN => n3087
                           );
   U1618 : AOI22_X1 port map( A1 => n6472, A2 => n6469, B1 => n6475, B2 => 
                           n6473, ZN => n6446);
   U1619 : AOI221_X1 port map( B1 => n5134, B2 => n5126, C1 => n7098, C2 => 
                           n5126, A => n3087, ZN => n6444);
   U1620 : NAND2_X1 port map( A1 => n6582, A2 => n6527, ZN => n6430);
   U1621 : NOR2_X1 port map( A1 => DATA2(14), A2 => n6427, ZN => n6725);
   U1622 : INV_X1 port map( A => DATA2(14), ZN => n6851);
   U1623 : NOR2_X1 port map( A1 => n6851, A2 => DATA1(14), ZN => n6729);
   U1624 : OAI21_X1 port map( B1 => n6725, B2 => n6729, A => n6631, ZN => n6429
                           );
   U1625 : NAND3_X1 port map( A1 => DATA2(14), A2 => n7169, A3 => n6528, ZN => 
                           n6428);
   U1626 : OAI211_X1 port map( C1 => n6431, C2 => n6430, A => n6429, B => n6428
                           , ZN => n6443);
   U1627 : AOI22_X1 port map( A1 => n6535, A2 => n6433, B1 => n6504, B2 => 
                           n6432, ZN => n6434);
   U1628 : INV_X1 port map( A => n6434, ZN => n6441);
   U1629 : INV_X1 port map( A => n6435, ZN => n6438);
   U1630 : AOI22_X1 port map( A1 => n6437, A2 => n6504, B1 => n6535, B2 => 
                           n6436, ZN => n6465);
   U1631 : NOR2_X1 port map( A1 => n6438, A2 => n6465, ZN => n6440);
   U1632 : MUX2_X1 port map( A => n6441, B => n6440, S => n6439, Z => n6442);
   U1633 : AOI211_X1 port map( C1 => n6641, C2 => n6444, A => n6443, B => n6442
                           , ZN => n6445);
   U1634 : OAI21_X1 port map( B1 => n6446, B2 => n6830, A => n6445, ZN => 
                           OUTALU(14));
   U1635 : NOR2_X1 port map( A1 => DATA2(13), A2 => n6447, ZN => n6724);
   U1636 : NOR2_X1 port map( A1 => n6852, A2 => DATA1(13), ZN => n6692);
   U1637 : NOR2_X1 port map( A1 => n6724, A2 => n6692, ZN => n6776);
   U1638 : OAI22_X1 port map( A1 => n6449, A2 => n6566, B1 => n6448, B2 => 
                           n6570, ZN => n6454);
   U1639 : OAI22_X1 port map( A1 => n6452, A2 => n6451, B1 => n6466, B2 => 
                           n6450, ZN => n6453);
   U1640 : OAI21_X1 port map( B1 => n6454, B2 => n6453, A => n6527, ZN => n6456
                           );
   U1641 : OAI211_X1 port map( C1 => n6493, C2 => n6633, A => DATA2(13), B => 
                           DATA1(13), ZN => n6455);
   U1642 : OAI211_X1 port map( C1 => n6776, C2 => n6492, A => n6456, B => n6455
                           , ZN => n6461);
   U1643 : AOI222_X1 port map( A1 => n6474, A2 => n6472, B1 => n6469, B2 => 
                           n6475, C1 => n6473, C2 => n6470, ZN => n6459);
   U1644 : INV_X1 port map( A => n6479, ZN => n6487);
   U1645 : NAND2_X1 port map( A1 => n6487, A2 => n6486, ZN => n6485);
   U1646 : OAI211_X1 port map( C1 => n6478, C2 => n6457, A => n6833, B => n6463
                           , ZN => n6458);
   U1647 : OAI22_X1 port map( A1 => n6459, A2 => n6830, B1 => n6485, B2 => 
                           n6458, ZN => n6460);
   U1648 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_13_port, A => 
                           n6461, B => n6460, ZN => n6462);
   U1649 : OAI221_X1 port map( B1 => n6465, B2 => n6464, C1 => n6465, C2 => 
                           n6463, A => n6462, ZN => OUTALU(13));
   U1650 : INV_X1 port map( A => n6466, ZN => n6525);
   U1651 : AOI222_X1 port map( A1 => n6525, A2 => n6468, B1 => n6494, B2 => 
                           n6495, C1 => n6467, C2 => n6526, ZN => n6490);
   U1652 : AOI22_X1 port map( A1 => n6472, A2 => n6471, B1 => n6470, B2 => 
                           n6469, ZN => n6477);
   U1653 : AOI22_X1 port map( A1 => n6475, A2 => n6474, B1 => n6595, B2 => 
                           n6473, ZN => n6476);
   U1654 : AOI21_X1 port map( B1 => n6477, B2 => n6476, A => n6830, ZN => n6484
                           );
   U1655 : OAI22_X1 port map( A1 => n6693, A2 => DATA2(12), B1 => n6853, B2 => 
                           n7168, ZN => n6812);
   U1656 : INV_X1 port map( A => n6812, ZN => n6722);
   U1657 : NAND3_X1 port map( A1 => DATA2(12), A2 => n7168, A3 => n6528, ZN => 
                           n6482);
   U1658 : INV_X1 port map( A => n6478, ZN => n6480);
   U1659 : OAI221_X1 port map( B1 => n6480, B2 => n6479, C1 => n6478, C2 => 
                           n6487, A => n6504, ZN => n6481);
   U1660 : OAI211_X1 port map( C1 => n6722, C2 => n6531, A => n6482, B => n6481
                           , ZN => n6483);
   U1661 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_12_port, A => 
                           n6484, B => n6483, ZN => n6489);
   U1662 : OAI211_X1 port map( C1 => n6487, C2 => n6486, A => n6535, B => n6485
                           , ZN => n6488);
   U1663 : OAI211_X1 port map( C1 => n6490, C2 => n6496, A => n6489, B => n6488
                           , ZN => OUTALU(12));
   U1664 : NAND2_X1 port map( A1 => DATA1(11), A2 => n6854, ZN => n6721);
   U1665 : NAND2_X1 port map( A1 => DATA2(11), A2 => n6491, ZN => n6720);
   U1666 : AOI21_X1 port map( B1 => n6721, B2 => n6720, A => n6492, ZN => n6500
                           );
   U1667 : AOI21_X1 port map( B1 => n6633, B2 => DATA1(11), A => n6493, ZN => 
                           n6498);
   U1668 : AOI22_X1 port map( A1 => n6495, A2 => n6525, B1 => n6526, B2 => 
                           n6494, ZN => n6497);
   U1669 : OAI22_X1 port map( A1 => n6498, A2 => n6854, B1 => n6497, B2 => 
                           n6496, ZN => n6499);
   U1670 : AOI211_X1 port map( C1 => dataout_mul_11_port, C2 => n6501, A => 
                           n6500, B => n6499, ZN => n6514);
   U1671 : INV_X1 port map( A => n6507, ZN => n6505);
   U1672 : OAI221_X1 port map( B1 => n6505, B2 => n6503, C1 => n6507, C2 => 
                           n6502, A => n6535, ZN => n6513);
   U1673 : INV_X1 port map( A => n6508, ZN => n6506);
   U1674 : OAI221_X1 port map( B1 => n6508, B2 => n6507, C1 => n6506, C2 => 
                           n6505, A => n6504, ZN => n6512);
   U1675 : NAND3_X1 port map( A1 => n6510, A2 => n6509, A3 => n6517, ZN => 
                           n6511);
   U1676 : NAND4_X1 port map( A1 => n6514, A2 => n6513, A3 => n6512, A4 => 
                           n6511, ZN => OUTALU(11));
   U1677 : AOI22_X1 port map( A1 => n6518, A2 => n6517, B1 => n6516, B2 => 
                           n6515, ZN => n6540);
   U1678 : NAND2_X1 port map( A1 => n6520, A2 => n6519, ZN => n6536);
   U1679 : INV_X1 port map( A => n6536, ZN => n6524);
   U1680 : AOI211_X1 port map( C1 => n6524, C2 => n6523, A => n6522, B => n6521
                           , ZN => n6533);
   U1681 : OAI22_X1 port map( A1 => n6662, A2 => n6855, B1 => DATA2(10), B2 => 
                           n7167, ZN => n6659);
   U1682 : NAND3_X1 port map( A1 => n6527, A2 => n6526, A3 => n6525, ZN => 
                           n6530);
   U1683 : NAND3_X1 port map( A1 => DATA2(10), A2 => n7167, A3 => n6528, ZN => 
                           n6529);
   U1684 : OAI211_X1 port map( C1 => n6659, C2 => n6531, A => n6530, B => n6529
                           , ZN => n6532);
   U1685 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_10_port, A => 
                           n6533, B => n6532, ZN => n6539);
   U1686 : OAI211_X1 port map( C1 => n6537, C2 => n6536, A => n6535, B => n6534
                           , ZN => n6538);
   U1687 : OAI211_X1 port map( C1 => n6540, C2 => n6830, A => n6539, B => n6538
                           , ZN => OUTALU(10));
   U1688 : INV_X1 port map( A => n6541, ZN => n6626);
   U1689 : AOI22_X1 port map( A1 => n6542, A2 => DATA1(3), B1 => n5185, B2 => 
                           DATA1(0), ZN => n6546);
   U1690 : NAND4_X1 port map( A1 => n6546, A2 => n6545, A3 => n6544, A4 => 
                           n6543, ZN => n6550);
   U1691 : AOI222_X1 port map( A1 => n6552, A2 => n6551, B1 => n6550, B2 => 
                           n6549, C1 => n6548, C2 => n6547, ZN => n6556);
   U1692 : INV_X1 port map( A => n6553, ZN => n6555);
   U1693 : OAI22_X1 port map( A1 => n6557, A2 => n6556, B1 => n6555, B2 => 
                           n6554, ZN => n6563);
   U1694 : OAI22_X1 port map( A1 => n6561, A2 => n6560, B1 => n6559, B2 => 
                           n6558, ZN => n6562);
   U1695 : AOI211_X1 port map( C1 => n6565, C2 => n6564, A => n6563, B => n6562
                           , ZN => n6567);
   U1696 : OAI22_X1 port map( A1 => n6569, A2 => n6568, B1 => n6567, B2 => 
                           n6566, ZN => n6575);
   U1697 : OAI22_X1 port map( A1 => n6573, A2 => n6572, B1 => n6571, B2 => 
                           n6570, ZN => n6574);
   U1698 : AOI211_X1 port map( C1 => n6577, C2 => n6576, A => n6575, B => n6574
                           , ZN => n6578);
   U1699 : INV_X1 port map( A => n6578, ZN => n6581);
   U1700 : AOI222_X1 port map( A1 => n6584, A2 => n6583, B1 => n6582, B2 => 
                           n6581, C1 => n6580, C2 => n6579, ZN => n6587);
   U1701 : OAI22_X1 port map( A1 => n6588, A2 => n6587, B1 => n6586, B2 => 
                           n6585, ZN => n6594);
   U1702 : OAI22_X1 port map( A1 => n6592, A2 => n6591, B1 => n6590, B2 => 
                           n6589, ZN => n6593);
   U1703 : AOI211_X1 port map( C1 => n6596, C2 => n6595, A => n6594, B => n6593
                           , ZN => n6597);
   U1704 : OAI22_X1 port map( A1 => n6600, A2 => n6599, B1 => n6598, B2 => 
                           n6597, ZN => n6601);
   U1705 : INV_X1 port map( A => n6601, ZN => n6607);
   U1706 : AOI22_X1 port map( A1 => n6605, A2 => n6604, B1 => n6603, B2 => 
                           n6602, ZN => n6606);
   U1707 : OAI211_X1 port map( C1 => n6609, C2 => n6608, A => n6607, B => n6606
                           , ZN => n6611);
   U1708 : AOI222_X1 port map( A1 => n6615, A2 => n6614, B1 => n6613, B2 => 
                           n6612, C1 => n6611, C2 => n6610, ZN => n6617);
   U1709 : OAI22_X1 port map( A1 => n6619, A2 => n6618, B1 => n6617, B2 => 
                           n6616, ZN => n6625);
   U1710 : OAI22_X1 port map( A1 => n6623, A2 => n6622, B1 => n6621, B2 => 
                           n6620, ZN => n6624);
   U1711 : AOI211_X1 port map( C1 => n6627, C2 => n6626, A => n6625, B => n6624
                           , ZN => n6831);
   U1712 : NOR3_X1 port map( A1 => n6629, A2 => n6832, A3 => n6628, ZN => n6640
                           );
   U1713 : OAI21_X1 port map( B1 => DATA1(0), B2 => DATA2_I_0_port, A => n6630,
                           ZN => n6638);
   U1714 : AOI22_X1 port map( A1 => DATA2(0), A2 => DATA1(0), B1 => n6696, B2 
                           => n6867, ZN => n6803);
   U1715 : AOI22_X1 port map( A1 => n6632, A2 => n6638, B1 => n6631, B2 => 
                           n6803, ZN => n6636);
   U1716 : OAI221_X1 port map( B1 => n6634, B2 => DATA2(0), C1 => n6634, C2 => 
                           n6633, A => DATA1(0), ZN => n6635);
   U1717 : OAI211_X1 port map( C1 => n6638, C2 => n6637, A => n6636, B => n6635
                           , ZN => n6639);
   U1718 : AOI211_X1 port map( C1 => n6641, C2 => dataout_mul_0_port, A => 
                           n6640, B => n6639, ZN => n6829);
   U1719 : AOI21_X1 port map( B1 => DATA1(26), B2 => n6839, A => n6764, ZN => 
                           n6802);
   U1720 : NOR2_X1 port map( A1 => n6742, A2 => n6642, ZN => n6785);
   U1721 : INV_X1 port map( A => n6643, ZN => n6738);
   U1722 : INV_X1 port map( A => n6644, ZN => n6730);
   U1723 : NOR2_X1 port map( A1 => n6725, A2 => n6730, ZN => n6796);
   U1724 : NOR2_X1 port map( A1 => DATA2(8), A2 => n6715, ZN => n6658);
   U1725 : AOI21_X1 port map( B1 => DATA1(6), B2 => n6861, A => n6712, ZN => 
                           n6797);
   U1726 : INV_X1 port map( A => n6704, ZN => n6655);
   U1727 : NAND2_X1 port map( A1 => DATA1(0), A2 => n6867, ZN => n6646);
   U1728 : INV_X1 port map( A => n6699, ZN => n6645);
   U1729 : OAI21_X1 port map( B1 => n6647, B2 => n6646, A => n6645, ZN => n6651
                           );
   U1730 : NOR2_X1 port map( A1 => DATA2(2), A2 => n6648, ZN => n6650);
   U1731 : INV_X1 port map( A => n6705, ZN => n6649);
   U1732 : AOI211_X1 port map( C1 => n6703, C2 => n6651, A => n6650, B => n6649
                           , ZN => n6653);
   U1733 : NAND2_X1 port map( A1 => n6652, A2 => n6707, ZN => n6815);
   U1734 : OAI21_X1 port map( B1 => n6653, B2 => n6815, A => n6710, ZN => n6654
                           );
   U1735 : OAI211_X1 port map( C1 => n6655, C2 => n6654, A => n6711, B => n6706
                           , ZN => n6656);
   U1736 : AOI211_X1 port map( C1 => n6797, C2 => n6656, A => n6694, B => n6813
                           , ZN => n6657);
   U1737 : OAI21_X1 port map( B1 => n6658, B2 => n6657, A => n6718, ZN => n6660
                           );
   U1738 : INV_X1 port map( A => n6659, ZN => n6716);
   U1739 : AOI21_X1 port map( B1 => n6661, B2 => n6660, A => n6716, ZN => n6663
                           );
   U1740 : OAI21_X1 port map( B1 => DATA2(10), B2 => n6662, A => n6721, ZN => 
                           n6799);
   U1741 : OAI211_X1 port map( C1 => n6663, C2 => n6799, A => n6722, B => n6720
                           , ZN => n6664);
   U1742 : OAI21_X1 port map( B1 => DATA2(12), B2 => n6693, A => n6664, ZN => 
                           n6666);
   U1743 : INV_X1 port map( A => n6729, ZN => n6793);
   U1744 : INV_X1 port map( A => n6692, ZN => n6665);
   U1745 : OAI211_X1 port map( C1 => n6724, C2 => n6666, A => n6793, B => n6665
                           , ZN => n6668);
   U1746 : NAND2_X1 port map( A1 => n6667, A2 => n6732, ZN => n6791);
   U1747 : AOI21_X1 port map( B1 => n6796, B2 => n6668, A => n6791, ZN => n6669
                           );
   U1748 : AOI221_X1 port map( B1 => n6731, B2 => n6738, C1 => n6669, C2 => 
                           n6738, A => n6737, ZN => n6672);
   U1749 : INV_X1 port map( A => n6806, ZN => n6671);
   U1750 : OAI211_X1 port map( C1 => n6741, C2 => n6672, A => n6671, B => n6670
                           , ZN => n6674);
   U1751 : INV_X1 port map( A => n6673, ZN => n6743);
   U1752 : AOI211_X1 port map( C1 => n6785, C2 => n6674, A => n6743, B => n6749
                           , ZN => n6676);
   U1753 : NOR3_X1 port map( A1 => n6676, A2 => n6675, A3 => n6748, ZN => n6678
                           );
   U1754 : OAI21_X1 port map( B1 => DATA2(22), B2 => n6677, A => n6754, ZN => 
                           n6801);
   U1755 : OAI211_X1 port map( C1 => n6678, C2 => n6801, A => n6755, B => n6752
                           , ZN => n6679);
   U1756 : OAI211_X1 port map( C1 => DATA2(24), C2 => n6680, A => n6679, B => 
                           n6759, ZN => n6681);
   U1757 : NAND3_X1 port map( A1 => n6758, A2 => n6681, A3 => n6690, ZN => 
                           n6682);
   U1758 : AOI211_X1 port map( C1 => n6802, C2 => n6682, A => n6762, B => n6810
                           , ZN => n6683);
   U1759 : AOI211_X1 port map( C1 => DATA1(28), C2 => n6837, A => n6683, B => 
                           n6770, ZN => n6685);
   U1760 : INV_X1 port map( A => n6684, ZN => n6771);
   U1761 : NOR3_X1 port map( A1 => n6685, A2 => n6766, A3 => n6771, ZN => n6688
                           );
   U1762 : NAND2_X1 port map( A1 => DATA1(31), A2 => n6834, ZN => n6687);
   U1763 : NAND2_X1 port map( A1 => DATA2(31), A2 => n6689, ZN => n6772);
   U1764 : OAI21_X1 port map( B1 => DATA2(30), B2 => n6686, A => n6772, ZN => 
                           n6804);
   U1765 : AOI221_X1 port map( B1 => n6688, B2 => n6687, C1 => n6804, C2 => 
                           n6687, A => FUNC(2), ZN => n6827);
   U1766 : OAI22_X1 port map( A1 => n6689, A2 => DATA2(31), B1 => n6835, B2 => 
                           DATA1(30), ZN => n6781);
   U1767 : OAI21_X1 port map( B1 => n6841, B2 => n6691, A => n6690, ZN => n6761
                           );
   U1768 : AOI21_X1 port map( B1 => DATA2(12), B2 => n6693, A => n6692, ZN => 
                           n6727);
   U1769 : AOI21_X1 port map( B1 => n6695, B2 => DATA2(6), A => n6694, ZN => 
                           n6807);
   U1770 : NAND2_X1 port map( A1 => DATA2(0), A2 => n6696, ZN => n6698);
   U1771 : OAI21_X1 port map( B1 => n6699, B2 => n6698, A => n6697, ZN => n6702
                           );
   U1772 : NOR2_X1 port map( A1 => DATA1(2), A2 => n6865, ZN => n6700);
   U1773 : AOI211_X1 port map( C1 => n6703, C2 => n6702, A => n6701, B => n6700
                           , ZN => n6708);
   U1774 : NAND2_X1 port map( A1 => n6705, A2 => n6704, ZN => n6809);
   U1775 : OAI211_X1 port map( C1 => n6708, C2 => n6809, A => n6707, B => n6706
                           , ZN => n6709);
   U1776 : NAND3_X1 port map( A1 => n6711, A2 => n6710, A3 => n6709, ZN => 
                           n6713);
   U1777 : AOI211_X1 port map( C1 => n6807, C2 => n6713, A => n6712, B => n6813
                           , ZN => n6714);
   U1778 : AOI21_X1 port map( B1 => DATA2(8), B2 => n6715, A => n6714, ZN => 
                           n6719);
   U1779 : AOI211_X1 port map( C1 => n6719, C2 => n6718, A => n6717, B => n6716
                           , ZN => n6723);
   U1780 : OAI21_X1 port map( B1 => n6855, B2 => n7167, A => n6720, ZN => n6784
                           );
   U1781 : OAI211_X1 port map( C1 => n6723, C2 => n6784, A => n6722, B => n6721
                           , ZN => n6726);
   U1782 : AOI211_X1 port map( C1 => n6727, C2 => n6726, A => n6725, B => n6724
                           , ZN => n6728);
   U1783 : NOR2_X1 port map( A1 => n6729, A2 => n6728, ZN => n6733);
   U1784 : AOI211_X1 port map( C1 => n6733, C2 => n6732, A => n6731, B => n6730
                           , ZN => n6734);
   U1785 : AOI21_X1 port map( B1 => DATA2(16), B2 => n6735, A => n6734, ZN => 
                           n6739);
   U1786 : AOI211_X1 port map( C1 => n6739, C2 => n6738, A => n6737, B => n6736
                           , ZN => n6740);
   U1787 : NOR2_X1 port map( A1 => n6741, A2 => n6740, ZN => n6745);
   U1788 : INV_X1 port map( A => n6742, ZN => n6744);
   U1789 : AOI211_X1 port map( C1 => n6745, C2 => n6744, A => n6743, B => n6806
                           , ZN => n6746);
   U1790 : AOI21_X1 port map( B1 => DATA2(20), B2 => n6747, A => n6746, ZN => 
                           n6751);
   U1791 : AOI211_X1 port map( C1 => n6751, C2 => n6750, A => n6749, B => n6748
                           , ZN => n6756);
   U1792 : OAI21_X1 port map( B1 => n6843, B2 => n6753, A => n6752, ZN => n6783
                           );
   U1793 : OAI211_X1 port map( C1 => n6756, C2 => n6783, A => n6755, B => n6754
                           , ZN => n6757);
   U1794 : INV_X1 port map( A => n6757, ZN => n6760);
   U1795 : OAI211_X1 port map( C1 => n6761, C2 => n6760, A => n6759, B => n6758
                           , ZN => n6765);
   U1796 : AOI21_X1 port map( B1 => DATA2(26), B2 => n6763, A => n6762, ZN => 
                           n6780);
   U1797 : AOI211_X1 port map( C1 => n6765, C2 => n6780, A => n6810, B => n6764
                           , ZN => n6767);
   U1798 : AOI211_X1 port map( C1 => n6768, C2 => DATA2(28), A => n6767, B => 
                           n6766, ZN => n6769);
   U1799 : NOR3_X1 port map( A1 => n6771, A2 => n6770, A3 => n6769, ZN => n6774
                           );
   U1800 : OAI211_X1 port map( C1 => n6781, C2 => n6774, A => n6773, B => n6772
                           , ZN => n6775);
   U1801 : INV_X1 port map( A => n6775, ZN => n6825);
   U1802 : NAND4_X1 port map( A1 => n6779, A2 => n6778, A3 => n6777, A4 => 
                           n6776, ZN => n6823);
   U1803 : INV_X1 port map( A => n6780, ZN => n6782);
   U1804 : OR4_X1 port map( A1 => n6784, A2 => n6783, A3 => n6782, A4 => n6781,
                           ZN => n6822);
   U1805 : INV_X1 port map( A => n6785, ZN => n6792);
   U1806 : NAND4_X1 port map( A1 => n6789, A2 => n6788, A3 => n6787, A4 => 
                           n6786, ZN => n6790);
   U1807 : NOR3_X1 port map( A1 => n6792, A2 => n6791, A3 => n6790, ZN => n6794
                           );
   U1808 : NAND4_X1 port map( A1 => FUNC(2), A2 => n6795, A3 => n6794, A4 => 
                           n6793, ZN => n6821);
   U1809 : INV_X1 port map( A => n6796, ZN => n6800);
   U1810 : INV_X1 port map( A => n6797, ZN => n6798);
   U1811 : NOR4_X1 port map( A1 => n6801, A2 => n6800, A3 => n6799, A4 => n6798
                           , ZN => n6819);
   U1812 : INV_X1 port map( A => n6802, ZN => n6805);
   U1813 : NOR4_X1 port map( A1 => n6806, A2 => n6805, A3 => n6804, A4 => n6803
                           , ZN => n6818);
   U1814 : INV_X1 port map( A => n6807, ZN => n6808);
   U1815 : NOR4_X1 port map( A1 => n6811, A2 => n6810, A3 => n6809, A4 => n6808
                           , ZN => n6817);
   U1816 : NOR4_X1 port map( A1 => n6815, A2 => n6814, A3 => n6813, A4 => n6812
                           , ZN => n6816);
   U1817 : NAND4_X1 port map( A1 => n6819, A2 => n6818, A3 => n6817, A4 => 
                           n6816, ZN => n6820);
   U1818 : NOR4_X1 port map( A1 => n6823, A2 => n6822, A3 => n6821, A4 => n6820
                           , ZN => n6824);
   U1819 : AOI211_X1 port map( C1 => n6832, C2 => n6825, A => n6824, B => 
                           FUNC(1), ZN => n6826);
   U1820 : OAI211_X1 port map( C1 => n6827, C2 => n6832, A => FUNC(0), B => 
                           n6826, ZN => n6828);
   U1821 : OAI211_X1 port map( C1 => n6831, C2 => n6830, A => n6829, B => n6828
                           , ZN => OUTALU(0));
   U1822 : NAND2_X1 port map( A1 => n6833, A2 => n6832, ZN => n6869);
   U1823 : CLKBUF_X1 port map( A => n6869, Z => n6859);
   U1824 : NAND2_X1 port map( A1 => FUNC(3), A2 => n6833, ZN => n6868);
   U1825 : AOI22_X1 port map( A1 => DATA2(31), A2 => n6859, B1 => n6858, B2 => 
                           n6834, ZN => N2548);
   U1826 : AOI22_X1 port map( A1 => DATA2(30), A2 => n6869, B1 => n6868, B2 => 
                           n6835, ZN => N2547);
   U1827 : AOI22_X1 port map( A1 => DATA2(29), A2 => n6859, B1 => n6858, B2 => 
                           n6836, ZN => N2546);
   U1828 : AOI22_X1 port map( A1 => DATA2(28), A2 => n6869, B1 => n6868, B2 => 
                           n6837, ZN => N2545);
   U1829 : AOI22_X1 port map( A1 => DATA2(27), A2 => n6859, B1 => n6858, B2 => 
                           n6838, ZN => N2544);
   U1830 : AOI22_X1 port map( A1 => DATA2(26), A2 => n6869, B1 => n6868, B2 => 
                           n6839, ZN => N2543);
   U1831 : AOI22_X1 port map( A1 => DATA2(25), A2 => n6859, B1 => n6858, B2 => 
                           n6840, ZN => N2542);
   U1832 : AOI22_X1 port map( A1 => DATA2(24), A2 => n6869, B1 => n6868, B2 => 
                           n6841, ZN => N2541);
   U1833 : AOI22_X1 port map( A1 => DATA2(23), A2 => n6859, B1 => n6858, B2 => 
                           n6842, ZN => N2540);
   U1834 : AOI22_X1 port map( A1 => DATA2(22), A2 => n6869, B1 => n6868, B2 => 
                           n6843, ZN => N2539);
   U1835 : INV_X1 port map( A => DATA2(21), ZN => n6844);
   U1836 : AOI22_X1 port map( A1 => DATA2(21), A2 => n6869, B1 => n6868, B2 => 
                           n6844, ZN => N2538);
   U1837 : AOI22_X1 port map( A1 => DATA2(20), A2 => n6869, B1 => n6868, B2 => 
                           n6845, ZN => N2537);
   U1838 : AOI22_X1 port map( A1 => DATA2(19), A2 => n6859, B1 => n6858, B2 => 
                           n6846, ZN => N2536);
   U1839 : AOI22_X1 port map( A1 => DATA2(18), A2 => n6859, B1 => n6858, B2 => 
                           n6847, ZN => N2535);
   U1840 : AOI22_X1 port map( A1 => DATA2(17), A2 => n6859, B1 => n6858, B2 => 
                           n6848, ZN => N2534);
   U1841 : AOI22_X1 port map( A1 => DATA2(16), A2 => n6859, B1 => n6858, B2 => 
                           n6849, ZN => N2533);
   U1842 : AOI22_X1 port map( A1 => DATA2(15), A2 => n6859, B1 => n6858, B2 => 
                           n6850, ZN => N2532);
   U1843 : AOI22_X1 port map( A1 => DATA2(14), A2 => n6859, B1 => n6858, B2 => 
                           n6851, ZN => N2531);
   U1844 : AOI22_X1 port map( A1 => DATA2(13), A2 => n6859, B1 => n6858, B2 => 
                           n6852, ZN => N2530);
   U1845 : AOI22_X1 port map( A1 => DATA2(12), A2 => n6859, B1 => n6858, B2 => 
                           n6853, ZN => N2529);
   U1846 : AOI22_X1 port map( A1 => DATA2(11), A2 => n6859, B1 => n6858, B2 => 
                           n6854, ZN => N2528);
   U1847 : AOI22_X1 port map( A1 => DATA2(10), A2 => n6859, B1 => n6858, B2 => 
                           n6855, ZN => N2527);
   U1848 : INV_X1 port map( A => DATA2(9), ZN => n6856);
   U1849 : AOI22_X1 port map( A1 => DATA2(9), A2 => n6859, B1 => n6858, B2 => 
                           n6856, ZN => N2526);
   U1850 : AOI22_X1 port map( A1 => DATA2(8), A2 => n6859, B1 => n6858, B2 => 
                           n6857, ZN => N2525);
   U1851 : AOI22_X1 port map( A1 => DATA2(7), A2 => n6869, B1 => n6868, B2 => 
                           n6860, ZN => N2524);
   U1852 : AOI22_X1 port map( A1 => DATA2(6), A2 => n6869, B1 => n6868, B2 => 
                           n6861, ZN => N2523);
   U1853 : AOI22_X1 port map( A1 => DATA2(5), A2 => n6869, B1 => n6868, B2 => 
                           n6862, ZN => N2522);
   U1854 : AOI22_X1 port map( A1 => DATA2(4), A2 => n6869, B1 => n6868, B2 => 
                           n6863, ZN => N2521);
   U1855 : AOI22_X1 port map( A1 => DATA2(3), A2 => n6869, B1 => n6868, B2 => 
                           n6864, ZN => N2520);
   U1856 : AOI22_X1 port map( A1 => DATA2(2), A2 => n6869, B1 => n6868, B2 => 
                           n6865, ZN => N2519);
   U1857 : AOI22_X1 port map( A1 => DATA2(1), A2 => n6869, B1 => n6868, B2 => 
                           n6866, ZN => N2518);
   U1858 : AOI22_X1 port map( A1 => DATA2(0), A2 => n6869, B1 => n6868, B2 => 
                           n6867, ZN => N2517);
   U1859 : NOR2_X1 port map( A1 => n6870, A2 => n1990, ZN => 
                           boothmul_pipelined_i_sum_out_1_0_port);
   U1860 : NAND2_X1 port map( A1 => n6911, A2 => data2_mul_3_port, ZN => n6874)
                           ;
   U1861 : INV_X1 port map( A => data2_mul_3_port, ZN => n6907);
   U1862 : NAND3_X1 port map( A1 => data2_mul_2_port, A2 => data2_mul_1_port, 
                           A3 => n6907, ZN => n6906);
   U1863 : INV_X1 port map( A => n6871, ZN => n6872);
   U1864 : NOR2_X1 port map( A1 => n6872, A2 => n6907, ZN => n6909);
   U1865 : NOR2_X1 port map( A1 => data2_mul_3_port, A2 => n6872, ZN => n6899);
   U1866 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n6909, B1 => data1_mul_1_port, B2 => n6899, ZN
                           => n6873);
   U1867 : OAI221_X1 port map( B1 => n1990, B2 => n6874, C1 => n1990, C2 => 
                           n6906, A => n6873, ZN => 
                           boothmul_pipelined_i_mux_out_1_3_port);
   U1868 : INV_X1 port map( A => n6874, ZN => n6908);
   U1869 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n6899, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n6908, ZN => n6876);
   U1870 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n6909, ZN => n6875);
   U1871 : OAI211_X1 port map( C1 => n1989, C2 => n6906, A => n6876, B => n6875
                           , ZN => boothmul_pipelined_i_mux_out_1_4_port);
   U1872 : CLKBUF_X1 port map( A => n6899, Z => n6903);
   U1873 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n6908, B1 => n6903, B2 => data1_mul_3_port, ZN
                           => n6878);
   U1874 : CLKBUF_X1 port map( A => n6909, Z => n6900);
   U1875 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, ZN => 
                           n6877);
   U1876 : OAI211_X1 port map( C1 => n6906, C2 => n1987, A => n6878, B => n6877
                           , ZN => boothmul_pipelined_i_mux_out_1_5_port);
   U1877 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_114_port, B1 => 
                           n6903, B2 => data1_mul_4_port, ZN => n6880);
   U1878 : NAND2_X1 port map( A1 => n6909, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, ZN => 
                           n6879);
   U1879 : OAI211_X1 port map( C1 => n1986, C2 => n6906, A => n6880, B => n6879
                           , ZN => boothmul_pipelined_i_mux_out_1_6_port);
   U1880 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_113_port, B1 => 
                           n6903, B2 => data1_mul_5_port, ZN => n6882);
   U1881 : NAND2_X1 port map( A1 => n6909, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, ZN => 
                           n6881);
   U1882 : OAI211_X1 port map( C1 => n1984, C2 => n6906, A => n6882, B => n6881
                           , ZN => boothmul_pipelined_i_mux_out_1_7_port);
   U1883 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_112_port, B1 => 
                           n6903, B2 => data1_mul_6_port, ZN => n6884);
   U1884 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, ZN => 
                           n6883);
   U1885 : OAI211_X1 port map( C1 => n1982, C2 => n6906, A => n6884, B => n6883
                           , ZN => boothmul_pipelined_i_mux_out_1_8_port);
   U1886 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_111_port, B1 => 
                           n6899, B2 => data1_mul_7_port, ZN => n6886);
   U1887 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, ZN => 
                           n6885);
   U1888 : OAI211_X1 port map( C1 => n1980, C2 => n6906, A => n6886, B => n6885
                           , ZN => boothmul_pipelined_i_mux_out_1_9_port);
   U1889 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_110_port, B1 => 
                           n6899, B2 => data1_mul_8_port, ZN => n6888);
   U1890 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, ZN => 
                           n6887);
   U1891 : OAI211_X1 port map( C1 => n1978, C2 => n6906, A => n6888, B => n6887
                           , ZN => boothmul_pipelined_i_mux_out_1_10_port);
   U1892 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_109_port, B1 => 
                           n6903, B2 => data1_mul_9_port, ZN => n6890);
   U1893 : NAND2_X1 port map( A1 => n6909, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, ZN => 
                           n6889);
   U1894 : OAI211_X1 port map( C1 => n1976, C2 => n6906, A => n6890, B => n6889
                           , ZN => boothmul_pipelined_i_mux_out_1_11_port);
   U1895 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_108_port, B1 => 
                           n6899, B2 => data1_mul_10_port, ZN => n6892);
   U1896 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, ZN => 
                           n6891);
   U1897 : OAI211_X1 port map( C1 => n1974, C2 => n6906, A => n6892, B => n6891
                           , ZN => boothmul_pipelined_i_mux_out_1_12_port);
   U1898 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_107_port, B1 => 
                           n6903, B2 => data1_mul_11_port, ZN => n6894);
   U1899 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, ZN => 
                           n6893);
   U1900 : OAI211_X1 port map( C1 => n1972, C2 => n6906, A => n6894, B => n6893
                           , ZN => boothmul_pipelined_i_mux_out_1_13_port);
   U1901 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_106_port, B1 => 
                           n6903, B2 => data1_mul_12_port, ZN => n6896);
   U1902 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, ZN => 
                           n6895);
   U1903 : OAI211_X1 port map( C1 => n1970, C2 => n6906, A => n6896, B => n6895
                           , ZN => boothmul_pipelined_i_mux_out_1_14_port);
   U1904 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_105_port, B1 => 
                           n6899, B2 => data1_mul_13_port, ZN => n6898);
   U1905 : NAND2_X1 port map( A1 => n6909, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, ZN => 
                           n6897);
   U1906 : OAI211_X1 port map( C1 => n1968, C2 => n6906, A => n6898, B => n6897
                           , ZN => boothmul_pipelined_i_mux_out_1_15_port);
   U1907 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_104_port, B1 => 
                           n6899, B2 => data1_mul_14_port, ZN => n6902);
   U1908 : NAND2_X1 port map( A1 => n6900, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n6901);
   U1909 : OAI211_X1 port map( C1 => n1966, C2 => n6906, A => n6902, B => n6901
                           , ZN => boothmul_pipelined_i_mux_out_1_16_port);
   U1910 : AOI22_X1 port map( A1 => n6908, A2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, B1 => 
                           n6903, B2 => data1_mul_15_port, ZN => n6905);
   U1911 : NAND2_X1 port map( A1 => n6909, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n6904);
   U1912 : OAI211_X1 port map( C1 => n1964, C2 => n6906, A => n6905, B => n6904
                           , ZN => boothmul_pipelined_i_mux_out_1_17_port);
   U1913 : NAND2_X1 port map( A1 => data1_mul_15_port, A2 => n6907, ZN => n6912
                           );
   U1914 : AOI22_X1 port map( A1 => n6909, A2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, B1 => 
                           n6908, B2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, ZN => 
                           n6910);
   U1915 : OAI21_X1 port map( B1 => n6912, B2 => n6911, A => n6910, ZN => 
                           boothmul_pipelined_i_mux_out_1_18_port);
   U1916 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n6951);
   U1917 : NAND2_X1 port map( A1 => n6951, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, ZN 
                           => n6915);
   U1918 : NAND3_X1 port map( A1 => n3076, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_2_4_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_2_3_port, 
                           ZN => n6947);
   U1919 : NOR2_X1 port map( A1 => n3076, A2 => n6913, ZN => n6928);
   U1920 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_2_5_port, A2 
                           => n6913, ZN => n6941);
   U1921 : CLKBUF_X1 port map( A => n6941, Z => n6944);
   U1922 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_116_port, 
                           A2 => n6928, B1 => data1_mul_1_port, B2 => n6944, ZN
                           => n6914);
   U1923 : OAI221_X1 port map( B1 => n1990, B2 => n6915, C1 => n1990, C2 => 
                           n6947, A => n6914, ZN => 
                           boothmul_pipelined_i_mux_out_2_5_port);
   U1924 : INV_X1 port map( A => n6915, ZN => n6949);
   U1925 : AOI22_X1 port map( A1 => data1_mul_2_port, A2 => n6941, B1 => 
                           boothmul_pipelined_i_muxes_in_0_116_port, B2 => 
                           n6949, ZN => n6917);
   U1926 : CLKBUF_X1 port map( A => n6928, Z => n6948);
   U1927 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n6948, ZN => n6916);
   U1928 : OAI211_X1 port map( C1 => n6947, C2 => n1989, A => n6917, B => n6916
                           , ZN => boothmul_pipelined_i_mux_out_2_6_port);
   U1929 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_115_port, 
                           A2 => n6949, B1 => data1_mul_3_port, B2 => n6944, ZN
                           => n6919);
   U1930 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n6928, ZN => n6918);
   U1931 : OAI211_X1 port map( C1 => n6947, C2 => n1987, A => n6919, B => n6918
                           , ZN => boothmul_pipelined_i_mux_out_2_7_port);
   U1932 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_114_port, 
                           A2 => n6949, B1 => data1_mul_4_port, B2 => n6944, ZN
                           => n6921);
   U1933 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n6928, ZN => n6920);
   U1934 : OAI211_X1 port map( C1 => n6947, C2 => n1986, A => n6921, B => n6920
                           , ZN => boothmul_pipelined_i_mux_out_2_8_port);
   U1935 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_113_port, 
                           A2 => n6949, B1 => data1_mul_5_port, B2 => n6941, ZN
                           => n6923);
   U1936 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n6928, ZN => n6922);
   U1937 : OAI211_X1 port map( C1 => n6947, C2 => n1984, A => n6923, B => n6922
                           , ZN => boothmul_pipelined_i_mux_out_2_9_port);
   U1938 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_112_port, 
                           A2 => n6949, B1 => data1_mul_6_port, B2 => n6944, ZN
                           => n6925);
   U1939 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n6928, ZN => n6924);
   U1940 : OAI211_X1 port map( C1 => n6947, C2 => n1982, A => n6925, B => n6924
                           , ZN => boothmul_pipelined_i_mux_out_2_10_port);
   U1941 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_111_port, 
                           A2 => n6949, B1 => data1_mul_7_port, B2 => n6941, ZN
                           => n6927);
   U1942 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n6928, ZN => n6926);
   U1943 : OAI211_X1 port map( C1 => n6947, C2 => n1980, A => n6927, B => n6926
                           , ZN => boothmul_pipelined_i_mux_out_2_11_port);
   U1944 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_110_port, 
                           A2 => n6949, B1 => data1_mul_8_port, B2 => n6944, ZN
                           => n6930);
   U1945 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n6928, ZN => n6929);
   U1946 : OAI211_X1 port map( C1 => n6947, C2 => n1978, A => n6930, B => n6929
                           , ZN => boothmul_pipelined_i_mux_out_2_12_port);
   U1947 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_109_port, 
                           A2 => n6949, B1 => data1_mul_9_port, B2 => n6944, ZN
                           => n6932);
   U1948 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n6948, ZN => n6931);
   U1949 : OAI211_X1 port map( C1 => n6947, C2 => n1976, A => n6932, B => n6931
                           , ZN => boothmul_pipelined_i_mux_out_2_13_port);
   U1950 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_108_port, 
                           A2 => n6949, B1 => data1_mul_10_port, B2 => n6941, 
                           ZN => n6934);
   U1951 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n6948, ZN => n6933);
   U1952 : OAI211_X1 port map( C1 => n6947, C2 => n1974, A => n6934, B => n6933
                           , ZN => boothmul_pipelined_i_mux_out_2_14_port);
   U1953 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_107_port, 
                           A2 => n6949, B1 => data1_mul_11_port, B2 => n6941, 
                           ZN => n6936);
   U1954 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n6948, ZN => n6935);
   U1955 : OAI211_X1 port map( C1 => n6947, C2 => n1972, A => n6936, B => n6935
                           , ZN => boothmul_pipelined_i_mux_out_2_15_port);
   U1956 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_106_port, 
                           A2 => n6949, B1 => data1_mul_12_port, B2 => n6944, 
                           ZN => n6938);
   U1957 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n6948, ZN => n6937);
   U1958 : OAI211_X1 port map( C1 => n6947, C2 => n1970, A => n6938, B => n6937
                           , ZN => boothmul_pipelined_i_mux_out_2_16_port);
   U1959 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_105_port, 
                           A2 => n6949, B1 => data1_mul_13_port, B2 => n6941, 
                           ZN => n6940);
   U1960 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n6948, ZN => n6939);
   U1961 : OAI211_X1 port map( C1 => n6947, C2 => n1968, A => n6940, B => n6939
                           , ZN => boothmul_pipelined_i_mux_out_2_17_port);
   U1962 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_104_port, 
                           A2 => n6949, B1 => data1_mul_14_port, B2 => n6941, 
                           ZN => n6943);
   U1963 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n6948, ZN => n6942);
   U1964 : OAI211_X1 port map( C1 => n6947, C2 => n1966, A => n6943, B => n6942
                           , ZN => boothmul_pipelined_i_mux_out_2_18_port);
   U1965 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_103_port, 
                           A2 => n6949, B1 => data1_mul_15_port, B2 => n6944, 
                           ZN => n6946);
   U1966 : NAND2_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n6948, ZN => n6945);
   U1967 : OAI211_X1 port map( C1 => n6947, C2 => n1964, A => n6946, B => n6945
                           , ZN => boothmul_pipelined_i_mux_out_2_19_port);
   U1968 : NAND2_X1 port map( A1 => n3076, A2 => data1_mul_15_port, ZN => n6952
                           );
   U1969 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_0_102_port, 
                           A2 => n6949, B1 => n6948, B2 => 
                           boothmul_pipelined_i_muxes_in_0_119_port, ZN => 
                           n6950);
   U1970 : OAI21_X1 port map( B1 => n6952, B2 => n6951, A => n6950, ZN => 
                           boothmul_pipelined_i_mux_out_2_20_port);
   U1971 : NAND3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n7162);
   U1972 : NOR3_X1 port map( A1 => n3082, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_3_6_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_3_5_port, 
                           ZN => n7160);
   U1973 : INV_X1 port map( A => n7160, ZN => n6955);
   U1974 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_3_7_port, A2 
                           => n6953, ZN => n7158);
   U1975 : CLKBUF_X1 port map( A => n7158, Z => n6985);
   U1976 : NOR2_X1 port map( A1 => n3082, A2 => n6953, ZN => n6968);
   U1977 : CLKBUF_X1 port map( A => n6968, Z => n7159);
   U1978 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_60_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_176_port, ZN
                           => n6954);
   U1979 : OAI221_X1 port map( B1 => n3077, B2 => n7162, C1 => n3077, C2 => 
                           n6955, A => n6954, ZN => 
                           boothmul_pipelined_i_mux_out_3_7_port);
   U1980 : INV_X1 port map( A => n7162, ZN => n6984);
   U1981 : CLKBUF_X1 port map( A => n7160, Z => n6981);
   U1982 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_3_60_port, A2
                           => n6984, B1 => n6981, B2 => 
                           boothmul_pipelined_i_muxes_in_3_176_port, ZN => 
                           n6957);
   U1983 : AOI22_X1 port map( A1 => n7158, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n6968
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n6956);
   U1984 : NAND2_X1 port map( A1 => n6957, A2 => n6956, ZN => 
                           boothmul_pipelined_i_mux_out_3_8_port);
   U1985 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_59_port, B1 => n7160
                           , B2 => boothmul_pipelined_i_muxes_in_3_175_port, ZN
                           => n6959);
   U1986 : AOI22_X1 port map( A1 => n7158, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n6968
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n6958);
   U1987 : NAND2_X1 port map( A1 => n6959, A2 => n6958, ZN => 
                           boothmul_pipelined_i_mux_out_3_9_port);
   U1988 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_58_port, B1 => n7160
                           , B2 => boothmul_pipelined_i_muxes_in_3_174_port, ZN
                           => n6961);
   U1989 : AOI22_X1 port map( A1 => n7158, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n6968
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n6960);
   U1990 : NAND2_X1 port map( A1 => n6961, A2 => n6960, ZN => 
                           boothmul_pipelined_i_mux_out_3_10_port);
   U1991 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_57_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_173_port, ZN
                           => n6963);
   U1992 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n6968
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n6962);
   U1993 : NAND2_X1 port map( A1 => n6963, A2 => n6962, ZN => 
                           boothmul_pipelined_i_mux_out_3_11_port);
   U1994 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_56_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_172_port, ZN
                           => n6965);
   U1995 : AOI22_X1 port map( A1 => n7158, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n6968
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n6964);
   U1996 : NAND2_X1 port map( A1 => n6965, A2 => n6964, ZN => 
                           boothmul_pipelined_i_mux_out_3_12_port);
   U1997 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_55_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_171_port, ZN
                           => n6967);
   U1998 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n6968
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n6966);
   U1999 : NAND2_X1 port map( A1 => n6967, A2 => n6966, ZN => 
                           boothmul_pipelined_i_mux_out_3_13_port);
   U2000 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_54_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_170_port, ZN
                           => n6970);
   U2001 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n6968
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n6969);
   U2002 : NAND2_X1 port map( A1 => n6970, A2 => n6969, ZN => 
                           boothmul_pipelined_i_mux_out_3_14_port);
   U2003 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_53_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_169_port, ZN
                           => n6972);
   U2004 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n6971);
   U2005 : NAND2_X1 port map( A1 => n6972, A2 => n6971, ZN => 
                           boothmul_pipelined_i_mux_out_3_15_port);
   U2006 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_52_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_168_port, ZN
                           => n6974);
   U2007 : AOI22_X1 port map( A1 => n7158, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n6973);
   U2008 : NAND2_X1 port map( A1 => n6974, A2 => n6973, ZN => 
                           boothmul_pipelined_i_mux_out_3_16_port);
   U2009 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_51_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_167_port, ZN
                           => n6976);
   U2010 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n6975);
   U2011 : NAND2_X1 port map( A1 => n6976, A2 => n6975, ZN => 
                           boothmul_pipelined_i_mux_out_3_17_port);
   U2012 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_50_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_166_port, ZN
                           => n6978);
   U2013 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n6977);
   U2014 : NAND2_X1 port map( A1 => n6978, A2 => n6977, ZN => 
                           boothmul_pipelined_i_mux_out_3_18_port);
   U2015 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_49_port, B1 => n7160
                           , B2 => boothmul_pipelined_i_muxes_in_3_165_port, ZN
                           => n6980);
   U2016 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n6979);
   U2017 : NAND2_X1 port map( A1 => n6980, A2 => n6979, ZN => 
                           boothmul_pipelined_i_mux_out_3_19_port);
   U2018 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_48_port, B1 => n6981
                           , B2 => boothmul_pipelined_i_muxes_in_3_164_port, ZN
                           => n6983);
   U2019 : AOI22_X1 port map( A1 => n7158, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n6982);
   U2020 : NAND2_X1 port map( A1 => n6983, A2 => n6982, ZN => 
                           boothmul_pipelined_i_mux_out_3_20_port);
   U2021 : AOI22_X1 port map( A1 => n6984, A2 => 
                           boothmul_pipelined_i_muxes_in_3_47_port, B1 => n7160
                           , B2 => boothmul_pipelined_i_muxes_in_3_163_port, ZN
                           => n6987);
   U2022 : AOI22_X1 port map( A1 => n6985, A2 => 
                           boothmul_pipelined_i_muxes_in_3_46_port, B1 => n7159
                           , B2 => boothmul_pipelined_i_muxes_in_3_162_port, ZN
                           => n6986);
   U2023 : NAND2_X1 port map( A1 => n6987, A2 => n6986, ZN => 
                           boothmul_pipelined_i_mux_out_3_21_port);
   U2024 : NAND3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n7146);
   U2025 : NOR3_X1 port map( A1 => n3078, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_4_8_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_4_7_port, 
                           ZN => n7144);
   U2026 : INV_X1 port map( A => n7144, ZN => n6991);
   U2027 : INV_X1 port map( A => n6989, ZN => n6988);
   U2028 : NAND2_X1 port map( A1 => n3078, A2 => n6988, ZN => n7147);
   U2029 : INV_X1 port map( A => n7147, ZN => n7017);
   U2030 : NOR2_X1 port map( A1 => n3078, A2 => n6989, ZN => n7021);
   U2031 : CLKBUF_X1 port map( A => n7021, Z => n7143);
   U2032 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_64_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_190_port, ZN
                           => n6990);
   U2033 : OAI221_X1 port map( B1 => n5121, B2 => n7146, C1 => n5121, C2 => 
                           n6991, A => n6990, ZN => 
                           boothmul_pipelined_i_mux_out_4_9_port);
   U2034 : INV_X1 port map( A => n7146, ZN => n7020);
   U2035 : CLKBUF_X1 port map( A => n7144, Z => n7016);
   U2036 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_4_64_port, A2
                           => n7020, B1 => n7016, B2 => 
                           boothmul_pipelined_i_muxes_in_4_190_port, ZN => 
                           n6993);
   U2037 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n7021
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n6992);
   U2038 : NAND2_X1 port map( A1 => n6993, A2 => n6992, ZN => 
                           boothmul_pipelined_i_mux_out_4_10_port);
   U2039 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_63_port, B1 => n7144
                           , B2 => boothmul_pipelined_i_muxes_in_4_189_port, ZN
                           => n6995);
   U2040 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n7021
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n6994);
   U2041 : NAND2_X1 port map( A1 => n6995, A2 => n6994, ZN => 
                           boothmul_pipelined_i_mux_out_4_11_port);
   U2042 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_62_port, B1 => n7144
                           , B2 => boothmul_pipelined_i_muxes_in_4_188_port, ZN
                           => n6997);
   U2043 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n7021
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n6996);
   U2044 : NAND2_X1 port map( A1 => n6997, A2 => n6996, ZN => 
                           boothmul_pipelined_i_mux_out_4_12_port);
   U2045 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_61_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_187_port, ZN
                           => n6999);
   U2046 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n6998);
   U2047 : NAND2_X1 port map( A1 => n6999, A2 => n6998, ZN => 
                           boothmul_pipelined_i_mux_out_4_13_port);
   U2048 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_60_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_186_port, ZN
                           => n7001);
   U2049 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n7021
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n7000);
   U2050 : NAND2_X1 port map( A1 => n7001, A2 => n7000, ZN => 
                           boothmul_pipelined_i_mux_out_4_14_port);
   U2051 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_59_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_185_port, ZN
                           => n7003);
   U2052 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n7002);
   U2053 : NAND2_X1 port map( A1 => n7003, A2 => n7002, ZN => 
                           boothmul_pipelined_i_mux_out_4_15_port);
   U2054 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_58_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_184_port, ZN
                           => n7005);
   U2055 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n7004);
   U2056 : NAND2_X1 port map( A1 => n7005, A2 => n7004, ZN => 
                           boothmul_pipelined_i_mux_out_4_16_port);
   U2057 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_57_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_183_port, ZN
                           => n7007);
   U2058 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n7006);
   U2059 : NAND2_X1 port map( A1 => n7007, A2 => n7006, ZN => 
                           boothmul_pipelined_i_mux_out_4_17_port);
   U2060 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_56_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_182_port, ZN
                           => n7009);
   U2061 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n7021
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n7008);
   U2062 : NAND2_X1 port map( A1 => n7009, A2 => n7008, ZN => 
                           boothmul_pipelined_i_mux_out_4_18_port);
   U2063 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_55_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_181_port, ZN
                           => n7011);
   U2064 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n7010);
   U2065 : NAND2_X1 port map( A1 => n7011, A2 => n7010, ZN => 
                           boothmul_pipelined_i_mux_out_4_19_port);
   U2066 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_54_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_180_port, ZN
                           => n7013);
   U2067 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n7012);
   U2068 : NAND2_X1 port map( A1 => n7013, A2 => n7012, ZN => 
                           boothmul_pipelined_i_mux_out_4_20_port);
   U2069 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_53_port, B1 => n7144
                           , B2 => boothmul_pipelined_i_muxes_in_4_179_port, ZN
                           => n7015);
   U2070 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n7143
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n7014);
   U2071 : NAND2_X1 port map( A1 => n7015, A2 => n7014, ZN => 
                           boothmul_pipelined_i_mux_out_4_21_port);
   U2072 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_52_port, B1 => n7016
                           , B2 => boothmul_pipelined_i_muxes_in_4_178_port, ZN
                           => n7019);
   U2073 : AOI22_X1 port map( A1 => n7017, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n7021
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n7018);
   U2074 : NAND2_X1 port map( A1 => n7019, A2 => n7018, ZN => 
                           boothmul_pipelined_i_mux_out_4_22_port);
   U2075 : AOI22_X1 port map( A1 => n7020, A2 => 
                           boothmul_pipelined_i_muxes_in_4_51_port, B1 => n7144
                           , B2 => boothmul_pipelined_i_muxes_in_4_177_port, ZN
                           => n7023);
   U2076 : NAND2_X1 port map( A1 => n7021, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, ZN => 
                           n7022);
   U2077 : OAI211_X1 port map( C1 => n5127, C2 => n7147, A => n7023, B => n7022
                           , ZN => boothmul_pipelined_i_mux_out_4_23_port);
   U2078 : NAND3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n7151);
   U2079 : NOR3_X1 port map( A1 => n3079, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_5_10_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_5_9_port, 
                           ZN => n7149);
   U2080 : INV_X1 port map( A => n7149, ZN => n7027);
   U2081 : INV_X1 port map( A => n7025, ZN => n7024);
   U2082 : NAND2_X1 port map( A1 => n3079, A2 => n7024, ZN => n7152);
   U2083 : INV_X1 port map( A => n7152, ZN => n7053);
   U2084 : NOR2_X1 port map( A1 => n3079, A2 => n7025, ZN => n7057);
   U2085 : CLKBUF_X1 port map( A => n7057, Z => n7148);
   U2086 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_68_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_204_port, ZN
                           => n7026);
   U2087 : OAI221_X1 port map( B1 => n5122, B2 => n7151, C1 => n5122, C2 => 
                           n7027, A => n7026, ZN => 
                           boothmul_pipelined_i_mux_out_5_11_port);
   U2088 : INV_X1 port map( A => n7151, ZN => n7056);
   U2089 : CLKBUF_X1 port map( A => n7149, Z => n7052);
   U2090 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_5_68_port, A2
                           => n7056, B1 => n7052, B2 => 
                           boothmul_pipelined_i_muxes_in_5_204_port, ZN => 
                           n7029);
   U2091 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n7057
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n7028);
   U2092 : NAND2_X1 port map( A1 => n7029, A2 => n7028, ZN => 
                           boothmul_pipelined_i_mux_out_5_12_port);
   U2093 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_67_port, B1 => n7149
                           , B2 => boothmul_pipelined_i_muxes_in_5_203_port, ZN
                           => n7031);
   U2094 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n7057
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n7030);
   U2095 : NAND2_X1 port map( A1 => n7031, A2 => n7030, ZN => 
                           boothmul_pipelined_i_mux_out_5_13_port);
   U2096 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_66_port, B1 => n7149
                           , B2 => boothmul_pipelined_i_muxes_in_5_202_port, ZN
                           => n7033);
   U2097 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n7057
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n7032);
   U2098 : NAND2_X1 port map( A1 => n7033, A2 => n7032, ZN => 
                           boothmul_pipelined_i_mux_out_5_14_port);
   U2099 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_65_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_201_port, ZN
                           => n7035);
   U2100 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n7034);
   U2101 : NAND2_X1 port map( A1 => n7035, A2 => n7034, ZN => 
                           boothmul_pipelined_i_mux_out_5_15_port);
   U2102 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_64_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_200_port, ZN
                           => n7037);
   U2103 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n7057
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n7036);
   U2104 : NAND2_X1 port map( A1 => n7037, A2 => n7036, ZN => 
                           boothmul_pipelined_i_mux_out_5_16_port);
   U2105 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_63_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_199_port, ZN
                           => n7039);
   U2106 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n7038);
   U2107 : NAND2_X1 port map( A1 => n7039, A2 => n7038, ZN => 
                           boothmul_pipelined_i_mux_out_5_17_port);
   U2108 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_62_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_198_port, ZN
                           => n7041);
   U2109 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n7040);
   U2110 : NAND2_X1 port map( A1 => n7041, A2 => n7040, ZN => 
                           boothmul_pipelined_i_mux_out_5_18_port);
   U2111 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_61_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_197_port, ZN
                           => n7043);
   U2112 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n7042);
   U2113 : NAND2_X1 port map( A1 => n7043, A2 => n7042, ZN => 
                           boothmul_pipelined_i_mux_out_5_19_port);
   U2114 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_60_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_196_port, ZN
                           => n7045);
   U2115 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n7057
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n7044);
   U2116 : NAND2_X1 port map( A1 => n7045, A2 => n7044, ZN => 
                           boothmul_pipelined_i_mux_out_5_20_port);
   U2117 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_59_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_195_port, ZN
                           => n7047);
   U2118 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n7046);
   U2119 : NAND2_X1 port map( A1 => n7047, A2 => n7046, ZN => 
                           boothmul_pipelined_i_mux_out_5_21_port);
   U2120 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_58_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_194_port, ZN
                           => n7049);
   U2121 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n7048);
   U2122 : NAND2_X1 port map( A1 => n7049, A2 => n7048, ZN => 
                           boothmul_pipelined_i_mux_out_5_22_port);
   U2123 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_57_port, B1 => n7149
                           , B2 => boothmul_pipelined_i_muxes_in_5_193_port, ZN
                           => n7051);
   U2124 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n7148
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n7050);
   U2125 : NAND2_X1 port map( A1 => n7051, A2 => n7050, ZN => 
                           boothmul_pipelined_i_mux_out_5_23_port);
   U2126 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_56_port, B1 => n7052
                           , B2 => boothmul_pipelined_i_muxes_in_5_192_port, ZN
                           => n7055);
   U2127 : AOI22_X1 port map( A1 => n7053, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n7057
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n7054);
   U2128 : NAND2_X1 port map( A1 => n7055, A2 => n7054, ZN => 
                           boothmul_pipelined_i_mux_out_5_24_port);
   U2129 : AOI22_X1 port map( A1 => n7056, A2 => 
                           boothmul_pipelined_i_muxes_in_5_55_port, B1 => n7149
                           , B2 => boothmul_pipelined_i_muxes_in_5_191_port, ZN
                           => n7059);
   U2130 : NAND2_X1 port map( A1 => n7057, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, ZN => 
                           n7058);
   U2131 : OAI211_X1 port map( C1 => n5128, C2 => n7152, A => n7059, B => n7058
                           , ZN => boothmul_pipelined_i_mux_out_5_25_port);
   U2132 : NAND3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n7156);
   U2133 : NOR3_X1 port map( A1 => n3080, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_6_12_port, A3 
                           => boothmul_pipelined_i_multiplicand_pip_6_11_port, 
                           ZN => n7154);
   U2134 : INV_X1 port map( A => n7154, ZN => n7063);
   U2135 : INV_X1 port map( A => n7061, ZN => n7060);
   U2136 : NAND2_X1 port map( A1 => n3080, A2 => n7060, ZN => n7157);
   U2137 : INV_X1 port map( A => n7157, ZN => n7089);
   U2138 : NOR2_X1 port map( A1 => n3080, A2 => n7061, ZN => n7093);
   U2139 : CLKBUF_X1 port map( A => n7093, Z => n7153);
   U2140 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_72_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_218_port, ZN
                           => n7062);
   U2141 : OAI221_X1 port map( B1 => n5123, B2 => n7156, C1 => n5123, C2 => 
                           n7063, A => n7062, ZN => 
                           boothmul_pipelined_i_mux_out_6_13_port);
   U2142 : INV_X1 port map( A => n7156, ZN => n7092);
   U2143 : CLKBUF_X1 port map( A => n7154, Z => n7088);
   U2144 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_6_72_port, A2
                           => n7092, B1 => n7088, B2 => 
                           boothmul_pipelined_i_muxes_in_6_218_port, ZN => 
                           n7065);
   U2145 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n7093
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n7064);
   U2146 : NAND2_X1 port map( A1 => n7065, A2 => n7064, ZN => 
                           boothmul_pipelined_i_mux_out_6_14_port);
   U2147 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_71_port, B1 => n7154
                           , B2 => boothmul_pipelined_i_muxes_in_6_217_port, ZN
                           => n7067);
   U2148 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n7093
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n7066);
   U2149 : NAND2_X1 port map( A1 => n7067, A2 => n7066, ZN => 
                           boothmul_pipelined_i_mux_out_6_15_port);
   U2150 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_70_port, B1 => n7154
                           , B2 => boothmul_pipelined_i_muxes_in_6_216_port, ZN
                           => n7069);
   U2151 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n7093
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n7068);
   U2152 : NAND2_X1 port map( A1 => n7069, A2 => n7068, ZN => 
                           boothmul_pipelined_i_mux_out_6_16_port);
   U2153 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_69_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_215_port, ZN
                           => n7071);
   U2154 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n7070);
   U2155 : NAND2_X1 port map( A1 => n7071, A2 => n7070, ZN => 
                           boothmul_pipelined_i_mux_out_6_17_port);
   U2156 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_68_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_214_port, ZN
                           => n7073);
   U2157 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n7093
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n7072);
   U2158 : NAND2_X1 port map( A1 => n7073, A2 => n7072, ZN => 
                           boothmul_pipelined_i_mux_out_6_18_port);
   U2159 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_67_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_213_port, ZN
                           => n7075);
   U2160 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n7074);
   U2161 : NAND2_X1 port map( A1 => n7075, A2 => n7074, ZN => 
                           boothmul_pipelined_i_mux_out_6_19_port);
   U2162 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_66_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_212_port, ZN
                           => n7077);
   U2163 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n7076);
   U2164 : NAND2_X1 port map( A1 => n7077, A2 => n7076, ZN => 
                           boothmul_pipelined_i_mux_out_6_20_port);
   U2165 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_65_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_211_port, ZN
                           => n7079);
   U2166 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n7078);
   U2167 : NAND2_X1 port map( A1 => n7079, A2 => n7078, ZN => 
                           boothmul_pipelined_i_mux_out_6_21_port);
   U2168 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_64_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_210_port, ZN
                           => n7081);
   U2169 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n7093
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n7080);
   U2170 : NAND2_X1 port map( A1 => n7081, A2 => n7080, ZN => 
                           boothmul_pipelined_i_mux_out_6_22_port);
   U2171 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_63_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_209_port, ZN
                           => n7083);
   U2172 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n7082);
   U2173 : NAND2_X1 port map( A1 => n7083, A2 => n7082, ZN => 
                           boothmul_pipelined_i_mux_out_6_23_port);
   U2174 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_62_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_208_port, ZN
                           => n7085);
   U2175 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n7084);
   U2176 : NAND2_X1 port map( A1 => n7085, A2 => n7084, ZN => 
                           boothmul_pipelined_i_mux_out_6_24_port);
   U2177 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_61_port, B1 => n7154
                           , B2 => boothmul_pipelined_i_muxes_in_6_207_port, ZN
                           => n7087);
   U2178 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n7153
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n7086);
   U2179 : NAND2_X1 port map( A1 => n7087, A2 => n7086, ZN => 
                           boothmul_pipelined_i_mux_out_6_25_port);
   U2180 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_60_port, B1 => n7088
                           , B2 => boothmul_pipelined_i_muxes_in_6_206_port, ZN
                           => n7091);
   U2181 : AOI22_X1 port map( A1 => n7089, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n7093
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n7090);
   U2182 : NAND2_X1 port map( A1 => n7091, A2 => n7090, ZN => 
                           boothmul_pipelined_i_mux_out_6_26_port);
   U2183 : AOI22_X1 port map( A1 => n7092, A2 => 
                           boothmul_pipelined_i_muxes_in_6_59_port, B1 => n7154
                           , B2 => boothmul_pipelined_i_muxes_in_6_205_port, ZN
                           => n7095);
   U2184 : NAND2_X1 port map( A1 => n7093, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, ZN => 
                           n7094);
   U2185 : OAI211_X1 port map( C1 => n5129, C2 => n7157, A => n7095, B => n7094
                           , ZN => boothmul_pipelined_i_mux_out_6_27_port);
   U2186 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, A2 
                           => n7096, ZN => n7114);
   U2187 : INV_X1 port map( A => n7114, ZN => n7100);
   U2188 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_13_port, A2 
                           => boothmul_pipelined_i_multiplicand_pip_7_14_port, 
                           ZN => n7097);
   U2189 : NAND2_X1 port map( A1 => n7097, A2 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, ZN 
                           => n7101);
   U2190 : NOR2_X1 port map( A1 => 
                           boothmul_pipelined_i_multiplicand_pip_7_15_port, A2 
                           => n7098, ZN => n7115);
   U2191 : CLKBUF_X1 port map( A => n7115, Z => n7134);
   U2192 : NOR2_X1 port map( A1 => n7098, A2 => n7165, ZN => n7135);
   U2193 : CLKBUF_X1 port map( A => n7135, Z => n7126);
   U2194 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_76_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_232_port, ZN
                           => n7099);
   U2195 : OAI221_X1 port map( B1 => n5134, B2 => n7100, C1 => n5134, C2 => 
                           n7101, A => n7099, ZN => 
                           boothmul_pipelined_i_mux_out_7_15_port);
   U2196 : INV_X1 port map( A => n7101, ZN => n7136);
   U2197 : AOI22_X1 port map( A1 => boothmul_pipelined_i_muxes_in_7_76_port, A2
                           => n7114, B1 => n7136, B2 => 
                           boothmul_pipelined_i_muxes_in_7_232_port, ZN => 
                           n7103);
   U2198 : AOI22_X1 port map( A1 => n7115, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_231_port, ZN
                           => n7102);
   U2199 : NAND2_X1 port map( A1 => n7103, A2 => n7102, ZN => 
                           boothmul_pipelined_i_mux_out_7_16_port);
   U2200 : CLKBUF_X1 port map( A => n7114, Z => n7133);
   U2201 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_75_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_231_port, ZN
                           => n7105);
   U2202 : AOI22_X1 port map( A1 => n7115, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_230_port, ZN
                           => n7104);
   U2203 : NAND2_X1 port map( A1 => n7105, A2 => n7104, ZN => 
                           boothmul_pipelined_i_mux_out_7_17_port);
   U2204 : AOI22_X1 port map( A1 => n7114, A2 => 
                           boothmul_pipelined_i_muxes_in_7_74_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_230_port, ZN
                           => n7107);
   U2205 : AOI22_X1 port map( A1 => n7115, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_229_port, ZN
                           => n7106);
   U2206 : NAND2_X1 port map( A1 => n7107, A2 => n7106, ZN => 
                           boothmul_pipelined_i_mux_out_7_18_port);
   U2207 : AOI22_X1 port map( A1 => n7114, A2 => 
                           boothmul_pipelined_i_muxes_in_7_73_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_229_port, ZN
                           => n7109);
   U2208 : AOI22_X1 port map( A1 => n7115, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_228_port, ZN
                           => n7108);
   U2209 : NAND2_X1 port map( A1 => n7109, A2 => n7108, ZN => 
                           boothmul_pipelined_i_mux_out_7_19_port);
   U2210 : AOI22_X1 port map( A1 => n7114, A2 => 
                           boothmul_pipelined_i_muxes_in_7_72_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_228_port, ZN
                           => n7111);
   U2211 : AOI22_X1 port map( A1 => n7115, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_227_port, ZN
                           => n7110);
   U2212 : NAND2_X1 port map( A1 => n7111, A2 => n7110, ZN => 
                           boothmul_pipelined_i_mux_out_7_20_port);
   U2213 : AOI22_X1 port map( A1 => n7114, A2 => 
                           boothmul_pipelined_i_muxes_in_7_71_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_227_port, ZN
                           => n7113);
   U2214 : AOI22_X1 port map( A1 => n7115, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => n7135
                           , B2 => boothmul_pipelined_i_muxes_in_7_226_port, ZN
                           => n7112);
   U2215 : NAND2_X1 port map( A1 => n7113, A2 => n7112, ZN => 
                           boothmul_pipelined_i_mux_out_7_21_port);
   U2216 : AOI22_X1 port map( A1 => n7114, A2 => 
                           boothmul_pipelined_i_muxes_in_7_70_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_226_port, ZN
                           => n7117);
   U2217 : AOI22_X1 port map( A1 => n7115, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_225_port, ZN
                           => n7116);
   U2218 : NAND2_X1 port map( A1 => n7117, A2 => n7116, ZN => 
                           boothmul_pipelined_i_mux_out_7_22_port);
   U2219 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_69_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_225_port, ZN
                           => n7119);
   U2220 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_224_port, ZN
                           => n7118);
   U2221 : NAND2_X1 port map( A1 => n7119, A2 => n7118, ZN => 
                           boothmul_pipelined_i_mux_out_7_23_port);
   U2222 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_68_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_224_port, ZN
                           => n7121);
   U2223 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => n7135
                           , B2 => boothmul_pipelined_i_muxes_in_7_223_port, ZN
                           => n7120);
   U2224 : NAND2_X1 port map( A1 => n7121, A2 => n7120, ZN => 
                           boothmul_pipelined_i_mux_out_7_24_port);
   U2225 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_67_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_223_port, ZN
                           => n7123);
   U2226 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => n7135
                           , B2 => boothmul_pipelined_i_muxes_in_7_222_port, ZN
                           => n7122);
   U2227 : NAND2_X1 port map( A1 => n7123, A2 => n7122, ZN => 
                           boothmul_pipelined_i_mux_out_7_25_port);
   U2228 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_66_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_222_port, ZN
                           => n7125);
   U2229 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => n7135
                           , B2 => boothmul_pipelined_i_muxes_in_7_221_port, ZN
                           => n7124);
   U2230 : NAND2_X1 port map( A1 => n7125, A2 => n7124, ZN => 
                           boothmul_pipelined_i_mux_out_7_26_port);
   U2231 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_65_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_221_port, ZN
                           => n7128);
   U2232 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => n7126
                           , B2 => boothmul_pipelined_i_muxes_in_7_220_port, ZN
                           => n7127);
   U2233 : NAND2_X1 port map( A1 => n7128, A2 => n7127, ZN => 
                           boothmul_pipelined_i_mux_out_7_27_port);
   U2234 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_64_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_220_port, ZN
                           => n7130);
   U2235 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => n7135
                           , B2 => boothmul_pipelined_i_muxes_in_7_219_port, ZN
                           => n7129);
   U2236 : NAND2_X1 port map( A1 => n7130, A2 => n7129, ZN => 
                           boothmul_pipelined_i_mux_out_7_28_port);
   U2237 : AOI22_X1 port map( A1 => n7133, A2 => 
                           boothmul_pipelined_i_muxes_in_7_63_port, B1 => n7136
                           , B2 => boothmul_pipelined_i_muxes_in_7_219_port, ZN
                           => n7132);
   U2238 : AOI22_X1 port map( A1 => n7134, A2 => 
                           boothmul_pipelined_i_muxes_in_7_62_port, B1 => n7135
                           , B2 => boothmul_pipelined_i_muxes_in_7_218_port, ZN
                           => n7131);
   U2239 : NAND2_X1 port map( A1 => n7132, A2 => n7131, ZN => 
                           boothmul_pipelined_i_mux_out_7_29_port);
   U2240 : OAI21_X1 port map( B1 => n7134, B2 => n7133, A => 
                           boothmul_pipelined_i_muxes_in_7_62_port, ZN => n7138
                           );
   U2241 : AOI22_X1 port map( A1 => n7136, A2 => 
                           boothmul_pipelined_i_muxes_in_7_218_port, B1 => 
                           n7135, B2 => 
                           boothmul_pipelined_i_muxes_in_7_217_port, ZN => 
                           n7137);
   U2242 : NAND2_X1 port map( A1 => n7138, A2 => n7137, ZN => 
                           boothmul_pipelined_i_mux_out_7_30_port);
   U2243 : AOI22_X1 port map( A1 => n7140, A2 => 
                           boothmul_pipelined_i_muxes_in_0_102_port, B1 => 
                           n7139, B2 => 
                           boothmul_pipelined_i_muxes_in_0_103_port, ZN => 
                           n7141);
   U2244 : OAI21_X1 port map( B1 => n7142, B2 => n1962, A => n7141, ZN => 
                           boothmul_pipelined_i_sum_B_in_1_15_port);
   U2245 : AOI22_X1 port map( A1 => n7144, A2 => 
                           boothmul_pipelined_i_muxes_in_4_176_port, B1 => 
                           n7143, B2 => 
                           boothmul_pipelined_i_muxes_in_4_175_port, ZN => 
                           n7145);
   U2246 : OAI221_X1 port map( B1 => n5127, B2 => n7147, C1 => n5127, C2 => 
                           n7146, A => n7145, ZN => n1997);
   U2247 : AOI22_X1 port map( A1 => n7149, A2 => 
                           boothmul_pipelined_i_muxes_in_5_190_port, B1 => 
                           n7148, B2 => 
                           boothmul_pipelined_i_muxes_in_5_189_port, ZN => 
                           n7150);
   U2248 : OAI221_X1 port map( B1 => n5128, B2 => n7152, C1 => n5128, C2 => 
                           n7151, A => n7150, ZN => n1996);
   U2249 : AOI22_X1 port map( A1 => n7154, A2 => 
                           boothmul_pipelined_i_muxes_in_6_204_port, B1 => 
                           n7153, B2 => 
                           boothmul_pipelined_i_muxes_in_6_203_port, ZN => 
                           n7155);
   U2250 : OAI221_X1 port map( B1 => n5129, B2 => n7157, C1 => n5129, C2 => 
                           n7156, A => n7155, ZN => n1995);
   U2251 : INV_X1 port map( A => n7158, ZN => n7163);
   U2252 : AOI22_X1 port map( A1 => n7160, A2 => 
                           boothmul_pipelined_i_muxes_in_3_162_port, B1 => 
                           n7159, B2 => 
                           boothmul_pipelined_i_muxes_in_3_161_port, ZN => 
                           n7161);
   U2253 : OAI221_X1 port map( B1 => n7164, B2 => n7163, C1 => n7164, C2 => 
                           n7162, A => n7161, ZN => n1991);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBITREG32_NBITADD5 is

   port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : 
         in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
         RESET_BAR : in std_logic);

end register_file_NBITREG32_NBITADD5;

architecture SYN_beh of register_file_NBITREG32_NBITADD5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N385, N386, N387, N388, N389, N390, N391, N392, N393
      , N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, 
      n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, 
      n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, 
      n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, 
      n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, 
      n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, 
      n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, 
      n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, 
      n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, 
      n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, 
      n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, 
      n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, 
      n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, 
      n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, 
      n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, 
      n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, 
      n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, 
      n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, 
      n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, 
      n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, 
      n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, 
      n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, 
      n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, 
      n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, 
      n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, 
      n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, 
      n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, 
      n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, 
      n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, 
      n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, 
      n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, 
      n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, 
      n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, 
      n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, 
      n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, 
      n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, 
      n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, 
      n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, 
      n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, 
      n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, 
      n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, 
      n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, 
      n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, 
      n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, 
      n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, 
      n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, 
      n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, 
      n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, 
      n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, 
      n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, 
      n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, 
      n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, 
      n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, 
      n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, 
      n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, 
      n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, 
      n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, 
      n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, 
      n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, 
      n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, 
      n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, 
      n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, 
      n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, 
      n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, 
      n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, 
      n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, 
      n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, 
      n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, 
      n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, 
      n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, 
      n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, 
      n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, 
      n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, 
      n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
      n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
      n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, 
      n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, 
      n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, 
      n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, 
      n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, 
      n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, 
      n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, 
      n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, 
      n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, 
      n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, 
      n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, 
      n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, 
      n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, 
      n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, 
      n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, 
      n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, 
      n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, 
      n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, 
      n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, 
      n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, 
      n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, 
      n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, 
      n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, 
      n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, 
      n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, 
      n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, 
      n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, 
      n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, 
      n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, 
      n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, 
      n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, 
      n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, 
      n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, 
      n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, 
      n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, 
      n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, 
      n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, 
      n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, 
      n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, 
      n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, 
      n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, 
      n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, 
      n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, 
      n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, 
      n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, 
      n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, 
      n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, 
      n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, 
      n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, 
      n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, 
      n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, 
      n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, 
      n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, 
      n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, 
      n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, 
      n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, 
      n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, 
      n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, 
      n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, 
      n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, 
      n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, 
      n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, 
      n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, 
      n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, 
      n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, 
      n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, 
      n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, 
      n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, 
      n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, 
      n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, 
      n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, 
      n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, 
      n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, 
      n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, 
      n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, 
      n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, 
      n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, 
      n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, 
      n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, 
      n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, 
      n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, 
      n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, 
      n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, 
      n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, 
      n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, 
      n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, 
      n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, 
      n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
      n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, 
      n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, 
      n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, 
      n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, 
      n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, 
      n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, 
      n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, 
      n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, 
      n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, 
      n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, 
      n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, 
      n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, 
      n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, 
      n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, 
      n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, 
      n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, 
      n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, 
      n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, 
      n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, 
      n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, 
      n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, 
      n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, 
      n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, 
      n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, 
      n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, 
      n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, 
      n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, 
      n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, 
      n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, 
      n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, 
      n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, 
      n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, 
      n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, 
      n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, 
      n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, 
      n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, 
      n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, 
      n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, 
      n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, 
      n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, 
      n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, 
      n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, 
      n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, 
      n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, 
      n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, 
      n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, 
      n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, 
      n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, 
      n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, 
      n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, 
      n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, 
      n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, 
      n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, 
      n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, 
      n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, 
      n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, 
      n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, 
      n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, 
      n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, 
      n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, 
      n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, 
      n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, 
      n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, 
      n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, 
      n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, 
      n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, 
      n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, 
      n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, 
      n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, 
      n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, 
      n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, 
      n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, 
      n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, 
      n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, 
      n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, 
      n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, 
      n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, 
      n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, 
      n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, 
      n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, 
      n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, 
      n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, 
      n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, 
      n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, 
      n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, 
      n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, 
      n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, 
      n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, 
      n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, 
      n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, 
      n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, 
      n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, 
      n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, 
      n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, 
      n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, 
      n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, 
      n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, 
      n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, 
      n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, 
      n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, 
      n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, 
      n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, 
      n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, 
      n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, 
      n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, 
      n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, 
      n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, 
      n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, 
      n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, 
      n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, 
      n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, 
      n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, 
      n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, 
      n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, 
      n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, 
      n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, 
      n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, 
      n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, 
      n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, 
      n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, 
      n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, 
      n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, 
      n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, 
      n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, 
      n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, 
      n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, 
      n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, 
      n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, 
      n11222, n11223, n11224, n11225, n_1349, n_1350, n_1351, n_1352, n_1353, 
      n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, 
      n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, 
      n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, 
      n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, 
      n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, 
      n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, 
      n_1408, n_1409, n_1410, n_1411, n_1412 : std_logic;

begin
   
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => 
                           REGISTERS_0_29_port, QN => n10722);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => 
                           REGISTERS_0_28_port, QN => n10723);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => 
                           REGISTERS_0_27_port, QN => n10453);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => 
                           REGISTERS_0_26_port, QN => n10724);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => 
                           REGISTERS_0_25_port, QN => n10454);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => 
                           REGISTERS_0_24_port, QN => n10455);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => 
                           REGISTERS_0_23_port, QN => n10456);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => 
                           REGISTERS_0_22_port, QN => n10457);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => 
                           REGISTERS_0_21_port, QN => n10458);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => 
                           REGISTERS_0_20_port, QN => n10208);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => 
                           REGISTERS_0_19_port, QN => n10459);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => 
                           REGISTERS_0_18_port, QN => n10209);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => 
                           REGISTERS_0_17_port, QN => n10460);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => 
                           REGISTERS_0_16_port, QN => n10725);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => 
                           REGISTERS_0_15_port, QN => n10461);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => 
                           REGISTERS_0_14_port, QN => n10462);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => 
                           REGISTERS_0_13_port, QN => n10210);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => 
                           REGISTERS_0_12_port, QN => n10463);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => 
                           REGISTERS_0_11_port, QN => n10211);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => 
                           REGISTERS_0_10_port, QN => n10464);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => 
                           REGISTERS_0_9_port, QN => n10465);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => 
                           REGISTERS_0_8_port, QN => n10466);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => 
                           REGISTERS_0_7_port, QN => n10987);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => 
                           REGISTERS_0_6_port, QN => n10212);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => 
                           REGISTERS_0_5_port, QN => n10467);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => 
                           REGISTERS_0_4_port, QN => n10468);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => 
                           REGISTERS_0_3_port, QN => n10213);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => 
                           REGISTERS_0_2_port, QN => n10726);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => 
                           REGISTERS_0_1_port, QN => n10469);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => 
                           REGISTERS_0_0_port, QN => n10470);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => 
                           REGISTERS_1_31_port, QN => n10471);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => 
                           REGISTERS_1_30_port, QN => n10472);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => 
                           REGISTERS_1_29_port, QN => n10214);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => 
                           REGISTERS_1_28_port, QN => n10473);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => 
                           REGISTERS_1_27_port, QN => n10215);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => 
                           REGISTERS_1_26_port, QN => n10216);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => 
                           REGISTERS_1_25_port, QN => n10988);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => 
                           REGISTERS_1_24_port, QN => n10727);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           REGISTERS_1_23_port, QN => n10728);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           REGISTERS_1_22_port, QN => n10217);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           REGISTERS_1_21_port, QN => n10218);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           REGISTERS_1_20_port, QN => n10474);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           REGISTERS_1_19_port, QN => n10219);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           REGISTERS_1_18_port, QN => n10989);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           REGISTERS_1_17_port, QN => n10990);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           REGISTERS_1_16_port, QN => n10220);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           REGISTERS_1_15_port, QN => n10221);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => 
                           REGISTERS_1_14_port, QN => n10475);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => 
                           REGISTERS_1_13_port, QN => n10476);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => 
                           REGISTERS_1_12_port, QN => n10222);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => 
                           REGISTERS_1_11_port, QN => n10477);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => 
                           REGISTERS_1_10_port, QN => n10478);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => 
                           REGISTERS_1_9_port, QN => n10991);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => 
                           REGISTERS_1_8_port, QN => n10729);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => 
                           REGISTERS_1_7_port, QN => n10223);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => 
                           REGISTERS_1_6_port, QN => n10479);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => 
                           REGISTERS_1_5_port, QN => n10992);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => 
                           REGISTERS_1_4_port, QN => n10730);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           REGISTERS_1_3_port, QN => n10480);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           REGISTERS_1_2_port, QN => n10481);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           REGISTERS_1_1_port, QN => n10993);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           REGISTERS_1_0_port, QN => n10224);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           REGISTERS_2_31_port, QN => n10482);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           REGISTERS_2_30_port, QN => n10225);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           REGISTERS_2_29_port, QN => n10483);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           REGISTERS_2_28_port, QN => n10226);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => 
                           REGISTERS_2_27_port, QN => n10484);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           REGISTERS_2_26_port, QN => n10227);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           REGISTERS_2_25_port, QN => n10485);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           REGISTERS_2_24_port, QN => n10486);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           REGISTERS_2_23_port, QN => n10228);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           REGISTERS_2_22_port, QN => n10229);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => 
                           REGISTERS_2_21_port, QN => n10230);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => 
                           REGISTERS_2_20_port, QN => n10487);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => 
                           REGISTERS_2_19_port, QN => n10231);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => 
                           REGISTERS_2_18_port, QN => n10232);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           REGISTERS_2_17_port, QN => n10233);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           REGISTERS_2_16_port, QN => n10488);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           REGISTERS_2_15_port, QN => n10234);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           REGISTERS_2_14_port, QN => n10235);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           REGISTERS_2_13_port, QN => n10489);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           REGISTERS_2_12_port, QN => n10490);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           REGISTERS_2_11_port, QN => n10491);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           REGISTERS_2_10_port, QN => n10492);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           REGISTERS_2_9_port, QN => n10236);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           REGISTERS_2_8_port, QN => n10237);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           REGISTERS_2_7_port, QN => n10493);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           REGISTERS_2_6_port, QN => n10238);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           REGISTERS_2_5_port, QN => n10239);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           REGISTERS_2_4_port, QN => n10240);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           REGISTERS_2_3_port, QN => n10494);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           REGISTERS_2_2_port, QN => n10241);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           REGISTERS_2_1_port, QN => n10242);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           REGISTERS_2_0_port, QN => n10495);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           REGISTERS_3_31_port, QN => n10731);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           REGISTERS_3_30_port, QN => n10994);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           REGISTERS_3_29_port, QN => n10995);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           REGISTERS_3_28_port, QN => n10732);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           REGISTERS_3_27_port, QN => n10243);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           REGISTERS_3_26_port, QN => n10496);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           REGISTERS_3_25_port, QN => n10244);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           REGISTERS_3_24_port, QN => n10497);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           REGISTERS_3_23_port, QN => n10733);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           REGISTERS_3_22_port, QN => n10498);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           REGISTERS_3_21_port, QN => n10245);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           REGISTERS_3_20_port, QN => n10734);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           REGISTERS_3_19_port, QN => n10246);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           REGISTERS_3_18_port, QN => n10499);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => 
                           REGISTERS_3_17_port, QN => n10735);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => 
                           REGISTERS_3_16_port, QN => n10500);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => 
                           REGISTERS_3_15_port, QN => n10996);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => 
                           REGISTERS_3_14_port, QN => n10247);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => 
                           REGISTERS_3_13_port, QN => n10997);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => 
                           REGISTERS_3_12_port, QN => n10736);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => 
                           REGISTERS_3_11_port, QN => n10737);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => 
                           REGISTERS_3_10_port, QN => n10738);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => 
                           REGISTERS_3_9_port, QN => n10998);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => 
                           REGISTERS_3_8_port, QN => n10999);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => 
                           REGISTERS_3_7_port, QN => n10248);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => 
                           REGISTERS_3_6_port, QN => n10501);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           REGISTERS_3_5_port, QN => n10249);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           REGISTERS_3_4_port, QN => n10502);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           REGISTERS_3_3_port, QN => n10250);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           REGISTERS_3_2_port, QN => n11000);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           REGISTERS_3_1_port, QN => n10251);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           REGISTERS_3_0_port, QN => n10739);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           REGISTERS_4_31_port, QN => n11001);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           REGISTERS_4_30_port, QN => n11002);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           REGISTERS_4_29_port, QN => n11003);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           REGISTERS_4_28_port, QN => n11004);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           REGISTERS_4_27_port, QN => n11005);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           REGISTERS_4_26_port, QN => n11006);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => 
                           REGISTERS_4_25_port, QN => n11007);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           REGISTERS_4_24_port, QN => n10740);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           REGISTERS_4_23_port, QN => n10741);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           REGISTERS_4_22_port, QN => n10742);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => 
                           REGISTERS_4_21_port, QN => n11008);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => 
                           REGISTERS_4_20_port, QN => n10743);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => 
                           REGISTERS_4_19_port, QN => n10744);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => 
                           REGISTERS_4_18_port, QN => n10745);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => 
                           REGISTERS_4_17_port, QN => n10503);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => 
                           REGISTERS_4_16_port, QN => n11009);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => 
                           REGISTERS_4_15_port, QN => n11010);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => 
                           REGISTERS_4_14_port, QN => n10746);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => 
                           REGISTERS_4_13_port, QN => n11011);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => 
                           REGISTERS_4_12_port, QN => n11012);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => 
                           REGISTERS_4_11_port, QN => n10747);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => 
                           REGISTERS_4_10_port, QN => n10252);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => 
                           REGISTERS_4_9_port, QN => n10253);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => 
                           REGISTERS_4_8_port, QN => n10504);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => 
                           REGISTERS_4_7_port, QN => n11013);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => 
                           REGISTERS_4_6_port, QN => n10748);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => 
                           REGISTERS_4_5_port, QN => n11014);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => 
                           REGISTERS_4_4_port, QN => n10749);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => 
                           REGISTERS_4_3_port, QN => n11015);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => 
                           REGISTERS_4_2_port, QN => n11016);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => 
                           REGISTERS_4_1_port, QN => n10750);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => 
                           REGISTERS_4_0_port, QN => n11017);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => 
                           REGISTERS_5_31_port, QN => n11018);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => 
                           REGISTERS_5_30_port, QN => n11019);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => 
                           REGISTERS_5_29_port, QN => n10254);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => 
                           REGISTERS_5_28_port, QN => n10505);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => 
                           REGISTERS_5_27_port, QN => n11020);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => 
                           REGISTERS_5_26_port, QN => n11021);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => 
                           REGISTERS_5_25_port, QN => n10751);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => 
                           REGISTERS_5_24_port, QN => n10255);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => 
                           REGISTERS_5_23_port, QN => n10506);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => 
                           REGISTERS_5_22_port, QN => n10752);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => 
                           REGISTERS_5_21_port, QN => n11022);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => 
                           REGISTERS_5_20_port, QN => n11023);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => 
                           REGISTERS_5_19_port, QN => n11024);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => 
                           REGISTERS_5_18_port, QN => n11025);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => 
                           REGISTERS_5_17_port, QN => n10753);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => 
                           REGISTERS_5_16_port, QN => n11026);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => 
                           REGISTERS_5_15_port, QN => n10754);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => 
                           REGISTERS_5_14_port, QN => n11027);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => 
                           REGISTERS_5_13_port, QN => n10755);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => 
                           REGISTERS_5_12_port, QN => n10256);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => 
                           REGISTERS_5_11_port, QN => n11028);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => 
                           REGISTERS_5_10_port, QN => n11029);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => 
                           REGISTERS_5_9_port, QN => n10756);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => 
                           REGISTERS_5_8_port, QN => n10757);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => 
                           REGISTERS_5_7_port, QN => n10758);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => 
                           REGISTERS_5_6_port, QN => n11030);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => 
                           REGISTERS_5_5_port, QN => n10759);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => 
                           REGISTERS_5_4_port, QN => n10760);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => 
                           REGISTERS_5_3_port, QN => n11031);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => 
                           REGISTERS_5_2_port, QN => n10507);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => 
                           REGISTERS_5_1_port, QN => n10761);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => 
                           REGISTERS_5_0_port, QN => n11032);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => 
                           REGISTERS_6_31_port, QN => n10762);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => 
                           REGISTERS_6_30_port, QN => n10763);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => 
                           REGISTERS_6_29_port, QN => n10764);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => 
                           REGISTERS_6_28_port, QN => n11033);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => 
                           REGISTERS_6_27_port, QN => n10765);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => 
                           REGISTERS_6_26_port, QN => n11034);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => 
                           REGISTERS_6_25_port, QN => n10766);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => 
                           REGISTERS_6_24_port, QN => n10767);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => 
                           REGISTERS_6_23_port, QN => n11035);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => 
                           REGISTERS_6_22_port, QN => n11036);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => 
                           REGISTERS_6_21_port, QN => n11037);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => 
                           REGISTERS_6_20_port, QN => n10768);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => 
                           REGISTERS_6_19_port, QN => n11038);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => 
                           REGISTERS_6_18_port, QN => n10769);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => 
                           REGISTERS_6_17_port, QN => n11039);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => 
                           REGISTERS_6_16_port, QN => n10770);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => 
                           REGISTERS_6_15_port, QN => n10771);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => 
                           REGISTERS_6_14_port, QN => n10772);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => 
                           REGISTERS_6_13_port, QN => n10773);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => 
                           REGISTERS_6_12_port, QN => n10774);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => 
                           REGISTERS_6_11_port, QN => n11040);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => 
                           REGISTERS_6_10_port, QN => n10775);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => 
                           REGISTERS_6_9_port, QN => n10776);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => 
                           REGISTERS_6_8_port, QN => n10777);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => 
                           REGISTERS_6_7_port, QN => n11041);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => 
                           REGISTERS_6_6_port, QN => n10778);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => 
                           REGISTERS_6_5_port, QN => n11042);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => 
                           REGISTERS_6_4_port, QN => n11043);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => 
                           REGISTERS_6_3_port, QN => n10779);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           REGISTERS_6_2_port, QN => n10780);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           REGISTERS_6_1_port, QN => n11044);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           REGISTERS_6_0_port, QN => n10781);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           REGISTERS_7_31_port, QN => n10257);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           REGISTERS_7_30_port, QN => n10258);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => 
                           REGISTERS_7_29_port, QN => n10508);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => 
                           REGISTERS_7_28_port, QN => n10259);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => 
                           REGISTERS_7_27_port, QN => n10782);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => 
                           REGISTERS_7_26_port, QN => n10260);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => 
                           REGISTERS_7_25_port, QN => n10261);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => 
                           REGISTERS_7_24_port, QN => n11045);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => 
                           REGISTERS_7_23_port, QN => n10509);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => 
                           REGISTERS_7_22_port, QN => n11046);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => 
                           REGISTERS_7_21_port, QN => n10783);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => 
                           REGISTERS_7_20_port, QN => n10510);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => 
                           REGISTERS_7_19_port, QN => n11047);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => 
                           REGISTERS_7_18_port, QN => n10511);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => 
                           REGISTERS_7_17_port, QN => n10262);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => 
                           REGISTERS_7_16_port, QN => n10263);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => 
                           REGISTERS_7_15_port, QN => n10512);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => 
                           REGISTERS_7_14_port, QN => n11048);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => 
                           REGISTERS_7_13_port, QN => n10264);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => 
                           REGISTERS_7_12_port, QN => n11049);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => 
                           REGISTERS_7_11_port, QN => n10265);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => 
                           REGISTERS_7_10_port, QN => n10784);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => 
                           REGISTERS_7_9_port, QN => n10513);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => 
                           REGISTERS_7_8_port, QN => n10514);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => 
                           REGISTERS_7_7_port, QN => n10266);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => 
                           REGISTERS_7_6_port, QN => n11050);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => 
                           REGISTERS_7_5_port, QN => n10267);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => 
                           REGISTERS_7_4_port, QN => n10515);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => 
                           REGISTERS_7_3_port, QN => n10785);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => 
                           REGISTERS_7_2_port, QN => n10268);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => 
                           REGISTERS_7_1_port, QN => n10516);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => 
                           REGISTERS_7_0_port, QN => n10269);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => 
                           REGISTERS_8_31_port, QN => n10270);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => 
                           REGISTERS_8_30_port, QN => n10517);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => 
                           REGISTERS_8_29_port, QN => n10786);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => 
                           REGISTERS_8_28_port, QN => n10518);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => 
                           REGISTERS_8_27_port, QN => n10787);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => 
                           REGISTERS_8_26_port, QN => n10271);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => 
                           REGISTERS_8_25_port, QN => n10519);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => 
                           REGISTERS_8_24_port, QN => n10520);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => 
                           REGISTERS_8_23_port, QN => n10521);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => 
                           REGISTERS_8_22_port, QN => n10272);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => 
                           REGISTERS_8_21_port, QN => n10788);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => 
                           REGISTERS_8_20_port, QN => n11051);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => 
                           REGISTERS_8_19_port, QN => n10273);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => 
                           REGISTERS_8_18_port, QN => n10522);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => 
                           REGISTERS_8_17_port, QN => n10274);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => 
                           REGISTERS_8_16_port, QN => n10523);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => 
                           REGISTERS_8_15_port, QN => n10275);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => 
                           REGISTERS_8_14_port, QN => n10276);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => 
                           REGISTERS_8_13_port, QN => n10277);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => 
                           REGISTERS_8_12_port, QN => n10278);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => 
                           REGISTERS_8_11_port, QN => n10524);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => 
                           REGISTERS_8_10_port, QN => n10279);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => 
                           REGISTERS_8_9_port, QN => n10525);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => 
                           REGISTERS_8_8_port, QN => n10526);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => 
                           REGISTERS_8_7_port, QN => n11052);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => 
                           REGISTERS_8_6_port, QN => n10280);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => 
                           REGISTERS_8_5_port, QN => n10281);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           REGISTERS_8_4_port, QN => n10282);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           REGISTERS_8_3_port, QN => n10527);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           REGISTERS_8_2_port, QN => n10528);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           REGISTERS_8_1_port, QN => n10283);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           REGISTERS_8_0_port, QN => n10284);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           REGISTERS_9_31_port, QN => n10529);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           REGISTERS_9_30_port, QN => n10530);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           REGISTERS_9_29_port, QN => n10285);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           REGISTERS_9_28_port, QN => n10531);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           REGISTERS_9_27_port, QN => n10532);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           REGISTERS_9_26_port, QN => n10533);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           REGISTERS_9_25_port, QN => n11053);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           REGISTERS_9_24_port, QN => n10286);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           REGISTERS_9_23_port, QN => n10789);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           REGISTERS_9_22_port, QN => n10287);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           REGISTERS_9_21_port, QN => n10288);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           REGISTERS_9_20_port, QN => n10534);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           REGISTERS_9_19_port, QN => n10535);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           REGISTERS_9_18_port, QN => n10536);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           REGISTERS_9_17_port, QN => n10289);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           REGISTERS_9_16_port, QN => n10290);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           REGISTERS_9_15_port, QN => n10537);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => 
                           REGISTERS_9_14_port, QN => n10790);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => 
                           REGISTERS_9_13_port, QN => n11054);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => 
                           REGISTERS_9_12_port, QN => n10291);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => 
                           REGISTERS_9_11_port, QN => n10292);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => 
                           REGISTERS_9_10_port, QN => n10538);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => 
                           REGISTERS_9_9_port, QN => n10791);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => 
                           REGISTERS_9_8_port, QN => n10792);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => 
                           REGISTERS_9_7_port, QN => n10293);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => 
                           REGISTERS_9_6_port, QN => n10294);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => 
                           REGISTERS_9_5_port, QN => n10539);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           REGISTERS_9_4_port, QN => n11055);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           REGISTERS_9_3_port, QN => n10540);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           REGISTERS_9_2_port, QN => n10793);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           REGISTERS_9_1_port, QN => n10794);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           REGISTERS_9_0_port, QN => n10795);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           REGISTERS_10_31_port, QN => n10295);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           REGISTERS_10_30_port, QN => n10296);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           REGISTERS_10_29_port, QN => n10297);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           REGISTERS_10_28_port, QN => n10541);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           REGISTERS_10_27_port, QN => n10298);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           REGISTERS_10_26_port, QN => n10542);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           REGISTERS_10_25_port, QN => n10299);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           REGISTERS_10_24_port, QN => n10300);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           REGISTERS_10_23_port, QN => n10543);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           REGISTERS_10_22_port, QN => n10544);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           REGISTERS_10_21_port, QN => n10301);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           REGISTERS_10_20_port, QN => n10545);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           REGISTERS_10_19_port, QN => n10302);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           REGISTERS_10_18_port, QN => n10303);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           REGISTERS_10_17_port, QN => n10546);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           REGISTERS_10_16_port, QN => n10547);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           REGISTERS_10_15_port, QN => n10548);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => 
                           REGISTERS_10_14_port, QN => n10549);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => 
                           REGISTERS_10_13_port, QN => n10304);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => 
                           REGISTERS_10_12_port, QN => n10550);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => 
                           REGISTERS_10_11_port, QN => n10551);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => 
                           REGISTERS_10_10_port, QN => n10552);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => 
                           REGISTERS_10_9_port, QN => n10305);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => 
                           REGISTERS_10_8_port, QN => n10553);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => 
                           REGISTERS_10_7_port, QN => n10554);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => 
                           REGISTERS_10_6_port, QN => n10555);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => 
                           REGISTERS_10_5_port, QN => n10556);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           REGISTERS_10_4_port, QN => n10306);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           REGISTERS_10_3_port, QN => n10307);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           REGISTERS_10_2_port, QN => n10557);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           REGISTERS_10_1_port, QN => n10308);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           REGISTERS_10_0_port, QN => n10558);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           REGISTERS_11_31_port, QN => n10796);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           REGISTERS_11_30_port, QN => n10309);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           REGISTERS_11_29_port, QN => n10310);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           REGISTERS_11_28_port, QN => n10797);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           REGISTERS_11_27_port, QN => n11056);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           REGISTERS_11_26_port, QN => n10798);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           REGISTERS_11_25_port, QN => n10311);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           REGISTERS_11_24_port, QN => n10799);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           REGISTERS_11_23_port, QN => n11057);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           REGISTERS_11_22_port, QN => n10800);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           REGISTERS_11_21_port, QN => n10801);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           REGISTERS_11_20_port, QN => n10312);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           REGISTERS_11_19_port, QN => n10802);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           REGISTERS_11_18_port, QN => n10803);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           REGISTERS_11_17_port, QN => n10559);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           REGISTERS_11_16_port, QN => n10804);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           REGISTERS_11_15_port, QN => n11058);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => 
                           REGISTERS_11_14_port, QN => n10560);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => 
                           REGISTERS_11_13_port, QN => n10561);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => 
                           REGISTERS_11_12_port, QN => n10805);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => 
                           REGISTERS_11_11_port, QN => n10313);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => 
                           REGISTERS_11_10_port, QN => n11059);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => 
                           REGISTERS_11_9_port, QN => n10562);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => 
                           REGISTERS_11_8_port, QN => n11060);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => 
                           REGISTERS_11_7_port, QN => n10563);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => 
                           REGISTERS_11_6_port, QN => n11061);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => 
                           REGISTERS_11_5_port, QN => n11062);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           REGISTERS_11_4_port, QN => n10564);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           REGISTERS_11_3_port, QN => n10806);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           REGISTERS_11_2_port, QN => n11063);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           REGISTERS_11_1_port, QN => n10565);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           REGISTERS_11_0_port, QN => n10314);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           REGISTERS_12_31_port, QN => n11064);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           REGISTERS_12_30_port, QN => n11065);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           REGISTERS_12_29_port, QN => n11066);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           REGISTERS_12_28_port, QN => n10807);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           REGISTERS_12_27_port, QN => n11067);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           REGISTERS_12_26_port, QN => n11068);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           REGISTERS_12_25_port, QN => n11069);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           REGISTERS_12_24_port, QN => n11070);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           REGISTERS_12_23_port, QN => n10315);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           REGISTERS_12_22_port, QN => n11071);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           REGISTERS_12_21_port, QN => n10566);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           REGISTERS_12_20_port, QN => n10808);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           REGISTERS_12_19_port, QN => n11072);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           REGISTERS_12_18_port, QN => n11073);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           REGISTERS_12_17_port, QN => n11074);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           REGISTERS_12_16_port, QN => n10809);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           REGISTERS_12_15_port, QN => n10567);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => 
                           REGISTERS_12_14_port, QN => n10810);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => 
                           REGISTERS_12_13_port, QN => n10568);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => 
                           REGISTERS_12_12_port, QN => n11075);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => 
                           REGISTERS_12_11_port, QN => n11076);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => 
                           REGISTERS_12_10_port, QN => n10811);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => 
                           REGISTERS_12_9_port, QN => n10812);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => 
                           REGISTERS_12_8_port, QN => n10316);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => 
                           REGISTERS_12_7_port, QN => n10813);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => 
                           REGISTERS_12_6_port, QN => n10814);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => 
                           REGISTERS_12_5_port, QN => n10815);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           REGISTERS_12_4_port, QN => n10816);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           REGISTERS_12_3_port, QN => n11077);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           REGISTERS_12_2_port, QN => n11078);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           REGISTERS_12_1_port, QN => n11079);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           REGISTERS_12_0_port, QN => n10569);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           REGISTERS_13_31_port, QN => n10817);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           REGISTERS_13_30_port, QN => n10818);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           REGISTERS_13_29_port, QN => n10570);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           REGISTERS_13_28_port, QN => n11080);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           REGISTERS_13_27_port, QN => n10317);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           REGISTERS_13_26_port, QN => n10819);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           REGISTERS_13_25_port, QN => n11081);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           REGISTERS_13_24_port, QN => n11082);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           REGISTERS_13_23_port, QN => n11083);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           REGISTERS_13_22_port, QN => n10820);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           REGISTERS_13_21_port, QN => n11084);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           REGISTERS_13_20_port, QN => n11085);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           REGISTERS_13_19_port, QN => n11086);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           REGISTERS_13_18_port, QN => n10821);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           REGISTERS_13_17_port, QN => n11087);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           REGISTERS_13_16_port, QN => n10822);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           REGISTERS_13_15_port, QN => n10823);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => 
                           REGISTERS_13_14_port, QN => n10571);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => 
                           REGISTERS_13_13_port, QN => n11088);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => 
                           REGISTERS_13_12_port, QN => n10572);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => 
                           REGISTERS_13_11_port, QN => n11089);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => 
                           REGISTERS_13_10_port, QN => n10318);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => 
                           REGISTERS_13_9_port, QN => n10319);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => 
                           REGISTERS_13_8_port, QN => n10824);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => 
                           REGISTERS_13_7_port, QN => n10825);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => 
                           REGISTERS_13_6_port, QN => n10826);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => 
                           REGISTERS_13_5_port, QN => n10827);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           REGISTERS_13_4_port, QN => n10828);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           REGISTERS_13_3_port, QN => n10573);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           REGISTERS_13_2_port, QN => n10320);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           REGISTERS_13_1_port, QN => n10574);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           REGISTERS_13_0_port, QN => n11090);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           REGISTERS_14_31_port, QN => n11091);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           REGISTERS_14_30_port, QN => n11092);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           REGISTERS_14_29_port, QN => n11093);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           REGISTERS_14_28_port, QN => n10829);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           REGISTERS_14_27_port, QN => n10830);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           REGISTERS_14_26_port, QN => n11094);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           REGISTERS_14_25_port, QN => n10831);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           REGISTERS_14_24_port, QN => n10832);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           REGISTERS_14_23_port, QN => n10833);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           REGISTERS_14_22_port, QN => n11095);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           REGISTERS_14_21_port, QN => n11096);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           REGISTERS_14_20_port, QN => n10834);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           REGISTERS_14_19_port, QN => n10835);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           REGISTERS_14_18_port, QN => n11097);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           REGISTERS_14_17_port, QN => n10836);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           REGISTERS_14_16_port, QN => n11098);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           REGISTERS_14_15_port, QN => n10837);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => 
                           REGISTERS_14_14_port, QN => n10838);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => 
                           REGISTERS_14_13_port, QN => n10839);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => 
                           REGISTERS_14_12_port, QN => n11099);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => 
                           REGISTERS_14_11_port, QN => n10840);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => 
                           REGISTERS_14_10_port, QN => n10841);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => 
                           REGISTERS_14_9_port, QN => n11100);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => 
                           REGISTERS_14_8_port, QN => n10842);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => 
                           REGISTERS_14_7_port, QN => n11101);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => 
                           REGISTERS_14_6_port, QN => n11102);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => 
                           REGISTERS_14_5_port, QN => n11103);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           REGISTERS_14_4_port, QN => n11104);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           REGISTERS_14_3_port, QN => n10843);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           REGISTERS_14_2_port, QN => n10844);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           REGISTERS_14_1_port, QN => n11105);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           REGISTERS_14_0_port, QN => n11106);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           REGISTERS_15_31_port, QN => n10575);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           REGISTERS_15_30_port, QN => n10845);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           REGISTERS_15_29_port, QN => n11107);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           REGISTERS_15_28_port, QN => n10321);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           REGISTERS_15_27_port, QN => n10576);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           REGISTERS_15_26_port, QN => n10322);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           REGISTERS_15_25_port, QN => n10323);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           REGISTERS_15_24_port, QN => n10577);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           REGISTERS_15_23_port, QN => n10324);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           REGISTERS_15_22_port, QN => n10578);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           REGISTERS_15_21_port, QN => n10579);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           REGISTERS_15_20_port, QN => n10325);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           REGISTERS_15_19_port, QN => n10580);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           REGISTERS_15_18_port, QN => n10326);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           REGISTERS_15_17_port, QN => n10846);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           REGISTERS_15_16_port, QN => n10581);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           REGISTERS_15_15_port, QN => n10847);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           REGISTERS_15_14_port, QN => n11108);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           REGISTERS_15_13_port, QN => n10848);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           REGISTERS_15_12_port, QN => n10849);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           REGISTERS_15_11_port, QN => n10850);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           REGISTERS_15_10_port, QN => n11109);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           REGISTERS_15_9_port, QN => n11110);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           REGISTERS_15_8_port, QN => n10582);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           REGISTERS_15_7_port, QN => n10327);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           REGISTERS_15_6_port, QN => n10583);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           REGISTERS_15_5_port, QN => n10328);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           REGISTERS_15_4_port, QN => n10584);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           REGISTERS_15_3_port, QN => n10851);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           REGISTERS_15_2_port, QN => n10329);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           REGISTERS_15_1_port, QN => n10852);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           REGISTERS_15_0_port, QN => n10853);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           REGISTERS_16_31_port, QN => n10445);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           REGISTERS_16_30_port, QN => n10330);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           REGISTERS_16_29_port, QN => n10585);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           REGISTERS_16_28_port, QN => n10586);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           REGISTERS_16_27_port, QN => n10587);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           REGISTERS_16_26_port, QN => n10588);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           REGISTERS_16_25_port, QN => n10854);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           REGISTERS_16_24_port, QN => n10589);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           REGISTERS_16_23_port, QN => n10590);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           REGISTERS_16_22_port, QN => n10591);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           REGISTERS_16_21_port, QN => n10592);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           REGISTERS_16_20_port, QN => n10593);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           REGISTERS_16_19_port, QN => n10594);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           REGISTERS_16_18_port, QN => n10595);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           REGISTERS_16_17_port, QN => n10855);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           REGISTERS_16_16_port, QN => n10331);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           REGISTERS_16_15_port, QN => n10332);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           REGISTERS_16_14_port, QN => n10596);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           REGISTERS_16_13_port, QN => n10597);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           REGISTERS_16_12_port, QN => n11111);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           REGISTERS_16_11_port, QN => n10333);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           REGISTERS_16_10_port, QN => n10334);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           REGISTERS_16_9_port, QN => n10598);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           REGISTERS_16_8_port, QN => n10335);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           REGISTERS_16_7_port, QN => n10599);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           REGISTERS_16_6_port, QN => n11112);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           REGISTERS_16_5_port, QN => n11113);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           REGISTERS_16_4_port, QN => n10600);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           REGISTERS_16_3_port, QN => n10336);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           REGISTERS_16_2_port, QN => n11114);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           REGISTERS_16_1_port, QN => n10601);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           REGISTERS_16_0_port, QN => n10337);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           REGISTERS_17_31_port, QN => n10202);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           REGISTERS_17_30_port, QN => n10338);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           REGISTERS_17_29_port, QN => n10602);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           REGISTERS_17_28_port, QN => n10339);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           REGISTERS_17_27_port, QN => n10603);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           REGISTERS_17_26_port, QN => n10604);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           REGISTERS_17_25_port, QN => n10605);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           REGISTERS_17_24_port, QN => n10340);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           REGISTERS_17_23_port, QN => n10606);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           REGISTERS_17_22_port, QN => n10607);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           REGISTERS_17_21_port, QN => n10341);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           REGISTERS_17_20_port, QN => n10608);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           REGISTERS_17_19_port, QN => n10609);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           REGISTERS_17_18_port, QN => n10610);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           REGISTERS_17_17_port, QN => n10611);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           REGISTERS_17_16_port, QN => n10342);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           REGISTERS_17_15_port, QN => n10612);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           REGISTERS_17_14_port, QN => n10343);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           REGISTERS_17_13_port, QN => n10344);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           REGISTERS_17_12_port, QN => n10345);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           REGISTERS_17_11_port, QN => n10613);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           REGISTERS_17_10_port, QN => n10614);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           REGISTERS_17_9_port, QN => n10615);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           REGISTERS_17_8_port, QN => n10616);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           REGISTERS_17_7_port, QN => n10346);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           REGISTERS_17_6_port, QN => n10347);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           REGISTERS_17_5_port, QN => n10348);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           REGISTERS_17_4_port, QN => n10617);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           REGISTERS_17_3_port, QN => n10618);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           REGISTERS_17_2_port, QN => n10619);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           REGISTERS_17_1_port, QN => n10349);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           REGISTERS_17_0_port, QN => n10620);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           REGISTERS_18_31_port, QN => n10446);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           REGISTERS_18_30_port, QN => n10350);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           REGISTERS_18_29_port, QN => n10621);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           REGISTERS_18_28_port, QN => n10351);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           REGISTERS_18_27_port, QN => n10352);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           REGISTERS_18_26_port, QN => n10353);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           REGISTERS_18_25_port, QN => n10354);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           REGISTERS_18_24_port, QN => n10355);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           REGISTERS_18_23_port, QN => n10356);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           REGISTERS_18_22_port, QN => n10357);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           REGISTERS_18_21_port, QN => n10358);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           REGISTERS_18_20_port, QN => n10622);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           REGISTERS_18_19_port, QN => n10359);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           REGISTERS_18_18_port, QN => n10360);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           REGISTERS_18_17_port, QN => n10623);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           REGISTERS_18_16_port, QN => n10361);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           REGISTERS_18_15_port, QN => n10362);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           REGISTERS_18_14_port, QN => n10363);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           REGISTERS_18_13_port, QN => n10624);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           REGISTERS_18_12_port, QN => n10364);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           REGISTERS_18_11_port, QN => n10365);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           REGISTERS_18_10_port, QN => n10366);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           REGISTERS_18_9_port, QN => n10367);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           REGISTERS_18_8_port, QN => n10856);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           REGISTERS_18_7_port, QN => n10625);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           REGISTERS_18_6_port, QN => n10626);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           REGISTERS_18_5_port, QN => n10627);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           REGISTERS_18_4_port, QN => n10368);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           REGISTERS_18_3_port, QN => n10628);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           REGISTERS_18_2_port, QN => n10369);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           REGISTERS_18_1_port, QN => n10629);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           REGISTERS_18_0_port, QN => n11115);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           REGISTERS_19_31_port, QN => n10718);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           REGISTERS_19_30_port, QN => n11116);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           REGISTERS_19_29_port, QN => n10857);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           REGISTERS_19_28_port, QN => n10630);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           REGISTERS_19_27_port, QN => n10858);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           REGISTERS_19_26_port, QN => n11117);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           REGISTERS_19_25_port, QN => n10859);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           REGISTERS_19_24_port, QN => n10860);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           REGISTERS_19_23_port, QN => n11118);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           REGISTERS_19_22_port, QN => n11119);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           REGISTERS_19_21_port, QN => n11120);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           REGISTERS_19_20_port, QN => n10861);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           REGISTERS_19_19_port, QN => n10631);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           REGISTERS_19_18_port, QN => n10862);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           REGISTERS_19_17_port, QN => n10863);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           REGISTERS_19_16_port, QN => n11121);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           REGISTERS_19_15_port, QN => n10370);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           REGISTERS_19_14_port, QN => n10864);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           REGISTERS_19_13_port, QN => n10865);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           REGISTERS_19_12_port, QN => n10371);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           REGISTERS_19_11_port, QN => n11122);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           REGISTERS_19_10_port, QN => n11123);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           REGISTERS_19_9_port, QN => n11124);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           REGISTERS_19_8_port, QN => n11125);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           REGISTERS_19_7_port, QN => n10372);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           REGISTERS_19_6_port, QN => n11126);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           REGISTERS_19_5_port, QN => n10632);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           REGISTERS_19_4_port, QN => n10866);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           REGISTERS_19_3_port, QN => n10633);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           REGISTERS_19_2_port, QN => n10867);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           REGISTERS_19_1_port, QN => n10373);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           REGISTERS_19_0_port, QN => n10868);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           REGISTERS_20_31_port, QN => n10447);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           REGISTERS_20_30_port, QN => n11127);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           REGISTERS_20_29_port, QN => n11128);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           REGISTERS_20_28_port, QN => n10869);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           REGISTERS_20_27_port, QN => n11129);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           REGISTERS_20_26_port, QN => n11130);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           REGISTERS_20_25_port, QN => n10634);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           REGISTERS_20_24_port, QN => n10635);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           REGISTERS_20_23_port, QN => n10870);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           REGISTERS_20_22_port, QN => n10374);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           REGISTERS_20_21_port, QN => n10636);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           REGISTERS_20_20_port, QN => n10871);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           REGISTERS_20_19_port, QN => n10872);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           REGISTERS_20_18_port, QN => n11131);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           REGISTERS_20_17_port, QN => n10637);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           REGISTERS_20_16_port, QN => n11132);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           REGISTERS_20_15_port, QN => n10638);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           REGISTERS_20_14_port, QN => n10873);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           REGISTERS_20_13_port, QN => n10874);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           REGISTERS_20_12_port, QN => n11133);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           REGISTERS_20_11_port, QN => n10875);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           REGISTERS_20_10_port, QN => n10876);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           REGISTERS_20_9_port, QN => n11134);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           REGISTERS_20_8_port, QN => n11135);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           REGISTERS_20_7_port, QN => n10877);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           REGISTERS_20_6_port, QN => n10375);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           REGISTERS_20_5_port, QN => n10878);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           REGISTERS_20_4_port, QN => n10879);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           REGISTERS_20_3_port, QN => n11136);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           REGISTERS_20_2_port, QN => n10376);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           REGISTERS_20_1_port, QN => n10880);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           REGISTERS_20_0_port, QN => n10639);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           REGISTERS_21_31_port, QN => n10719);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           REGISTERS_21_30_port, QN => n10881);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           REGISTERS_21_29_port, QN => n10377);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           REGISTERS_21_28_port, QN => n10882);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           REGISTERS_21_27_port, QN => n10883);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           REGISTERS_21_26_port, QN => n10884);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           REGISTERS_21_25_port, QN => n11137);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           REGISTERS_21_24_port, QN => n11138);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           REGISTERS_21_23_port, QN => n11139);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           REGISTERS_21_22_port, QN => n10885);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           REGISTERS_21_21_port, QN => n10886);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           REGISTERS_21_20_port, QN => n10887);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           REGISTERS_21_19_port, QN => n10888);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           REGISTERS_21_18_port, QN => n11140);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           REGISTERS_21_17_port, QN => n11141);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           REGISTERS_21_16_port, QN => n10378);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           REGISTERS_21_15_port, QN => n11142);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           REGISTERS_21_14_port, QN => n11143);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           REGISTERS_21_13_port, QN => n11144);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           REGISTERS_21_12_port, QN => n10640);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           REGISTERS_21_11_port, QN => n10889);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           REGISTERS_21_10_port, QN => n11145);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           REGISTERS_21_9_port, QN => n11146);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           REGISTERS_21_8_port, QN => n10890);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           REGISTERS_21_7_port, QN => n11147);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           REGISTERS_21_6_port, QN => n10891);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           REGISTERS_21_5_port, QN => n10892);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           REGISTERS_21_4_port, QN => n11148);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           REGISTERS_21_3_port, QN => n10893);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           REGISTERS_21_2_port, QN => n11149);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           REGISTERS_21_1_port, QN => n11150);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           REGISTERS_21_0_port, QN => n10379);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           REGISTERS_22_31_port, QN => n10448);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           REGISTERS_22_30_port, QN => n11151);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           REGISTERS_22_29_port, QN => n11152);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           REGISTERS_22_28_port, QN => n10894);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           REGISTERS_22_27_port, QN => n11153);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           REGISTERS_22_26_port, QN => n10641);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           REGISTERS_22_25_port, QN => n11154);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           REGISTERS_22_24_port, QN => n11155);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           REGISTERS_22_23_port, QN => n11156);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           REGISTERS_22_22_port, QN => n10895);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           REGISTERS_22_21_port, QN => n11157);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           REGISTERS_22_20_port, QN => n10896);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           REGISTERS_22_19_port, QN => n10897);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           REGISTERS_22_18_port, QN => n11158);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           REGISTERS_22_17_port, QN => n10898);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           REGISTERS_22_16_port, QN => n11159);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           REGISTERS_22_15_port, QN => n11160);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           REGISTERS_22_14_port, QN => n11161);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           REGISTERS_22_13_port, QN => n10899);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           REGISTERS_22_12_port, QN => n10900);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           REGISTERS_22_11_port, QN => n11162);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           REGISTERS_22_10_port, QN => n10642);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           REGISTERS_22_9_port, QN => n10901);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           REGISTERS_22_8_port, QN => n10643);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           REGISTERS_22_7_port, QN => n10902);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           REGISTERS_22_6_port, QN => n10903);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           REGISTERS_22_5_port, QN => n11163);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           REGISTERS_22_4_port, QN => n10904);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           REGISTERS_22_3_port, QN => n11164);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           REGISTERS_22_2_port, QN => n10380);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           REGISTERS_22_1_port, QN => n11165);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           REGISTERS_22_0_port, QN => n10905);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           REGISTERS_23_31_port, QN => n10203);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           REGISTERS_23_30_port, QN => n10906);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           REGISTERS_23_29_port, QN => n11166);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           REGISTERS_23_28_port, QN => n10381);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           REGISTERS_23_27_port, QN => n11167);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           REGISTERS_23_26_port, QN => n11168);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           REGISTERS_23_25_port, QN => n10382);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           REGISTERS_23_24_port, QN => n11169);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           REGISTERS_23_23_port, QN => n10383);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           REGISTERS_23_22_port, QN => n10644);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           REGISTERS_23_21_port, QN => n10907);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           REGISTERS_23_20_port, QN => n10645);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           REGISTERS_23_19_port, QN => n10384);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           REGISTERS_23_18_port, QN => n10646);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           REGISTERS_23_17_port, QN => n10385);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           REGISTERS_23_16_port, QN => n11170);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           REGISTERS_23_15_port, QN => n10908);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           REGISTERS_23_14_port, QN => n11171);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           REGISTERS_23_13_port, QN => n10909);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           REGISTERS_23_12_port, QN => n10647);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           REGISTERS_23_11_port, QN => n10648);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           REGISTERS_23_10_port, QN => n11172);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           REGISTERS_23_9_port, QN => n10910);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           REGISTERS_23_8_port, QN => n10649);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           REGISTERS_23_7_port, QN => n10386);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           REGISTERS_23_6_port, QN => n10650);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           REGISTERS_23_5_port, QN => n10651);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           REGISTERS_23_4_port, QN => n10911);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           REGISTERS_23_3_port, QN => n10387);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           REGISTERS_23_2_port, QN => n11173);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           REGISTERS_23_1_port, QN => n10912);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           REGISTERS_23_0_port, QN => n10388);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           REGISTERS_24_31_port, QN => n10449);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           REGISTERS_24_30_port, QN => n10389);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           REGISTERS_24_29_port, QN => n10390);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           REGISTERS_24_28_port, QN => n11174);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           REGISTERS_24_27_port, QN => n10652);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           REGISTERS_24_26_port, QN => n10913);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           REGISTERS_24_25_port, QN => n11175);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           REGISTERS_24_24_port, QN => n10653);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           REGISTERS_24_23_port, QN => n10654);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           REGISTERS_24_22_port, QN => n11176);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           REGISTERS_24_21_port, QN => n10655);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           REGISTERS_24_20_port, QN => n10391);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           REGISTERS_24_19_port, QN => n11177);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           REGISTERS_24_18_port, QN => n10914);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           REGISTERS_24_17_port, QN => n11178);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           REGISTERS_24_16_port, QN => n10656);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           REGISTERS_24_15_port, QN => n10915);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           REGISTERS_24_14_port, QN => n10392);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           REGISTERS_24_13_port, QN => n10657);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           REGISTERS_24_12_port, QN => n10916);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           REGISTERS_24_11_port, QN => n11179);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           REGISTERS_24_10_port, QN => n10658);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           REGISTERS_24_9_port, QN => n10393);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           REGISTERS_24_8_port, QN => n10394);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           REGISTERS_24_7_port, QN => n10659);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           REGISTERS_24_6_port, QN => n10395);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           REGISTERS_24_5_port, QN => n10396);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           REGISTERS_24_4_port, QN => n11180);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           REGISTERS_24_3_port, QN => n11181);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           REGISTERS_24_2_port, QN => n10397);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           REGISTERS_24_1_port, QN => n10660);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           REGISTERS_24_0_port, QN => n10398);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           REGISTERS_25_31_port, QN => n10450);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           REGISTERS_25_30_port, QN => n10917);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           REGISTERS_25_29_port, QN => n10918);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           REGISTERS_25_28_port, QN => n10919);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           REGISTERS_25_27_port, QN => n10399);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           REGISTERS_25_26_port, QN => n10920);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           REGISTERS_25_25_port, QN => n10661);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           REGISTERS_25_24_port, QN => n10400);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           REGISTERS_25_23_port, QN => n10401);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           REGISTERS_25_22_port, QN => n10921);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           REGISTERS_25_21_port, QN => n10922);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           REGISTERS_25_20_port, QN => n10662);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           REGISTERS_25_19_port, QN => n11182);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           REGISTERS_25_18_port, QN => n10663);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           REGISTERS_25_17_port, QN => n10402);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           REGISTERS_25_16_port, QN => n10403);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           REGISTERS_25_15_port, QN => n11183);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           REGISTERS_25_14_port, QN => n10923);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           REGISTERS_25_13_port, QN => n10664);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           REGISTERS_25_12_port, QN => n10665);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           REGISTERS_25_11_port, QN => n10924);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           REGISTERS_25_10_port, QN => n10925);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           REGISTERS_25_9_port, QN => n10404);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           REGISTERS_25_8_port, QN => n11184);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           REGISTERS_25_7_port, QN => n11185);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           REGISTERS_25_6_port, QN => n11186);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           REGISTERS_25_5_port, QN => n10405);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           REGISTERS_25_4_port, QN => n10666);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           REGISTERS_25_3_port, QN => n10406);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           REGISTERS_25_2_port, QN => n10926);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           REGISTERS_25_1_port, QN => n11187);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           REGISTERS_25_0_port, QN => n10927);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           REGISTERS_26_31_port, QN => n10720);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           REGISTERS_26_30_port, QN => n10667);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           REGISTERS_26_29_port, QN => n10668);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           REGISTERS_26_28_port, QN => n11188);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           REGISTERS_26_27_port, QN => n10407);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           REGISTERS_26_26_port, QN => n10669);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           REGISTERS_26_25_port, QN => n10408);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           REGISTERS_26_24_port, QN => n10670);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           REGISTERS_26_23_port, QN => n10671);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           REGISTERS_26_22_port, QN => n10409);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           REGISTERS_26_21_port, QN => n10672);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           REGISTERS_26_20_port, QN => n10410);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           REGISTERS_26_19_port, QN => n10673);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           REGISTERS_26_18_port, QN => n10674);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           REGISTERS_26_17_port, QN => n10411);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           REGISTERS_26_16_port, QN => n10675);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           REGISTERS_26_15_port, QN => n10412);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           REGISTERS_26_14_port, QN => n10676);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           REGISTERS_26_13_port, QN => n10677);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           REGISTERS_26_12_port, QN => n11189);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           REGISTERS_26_11_port, QN => n10413);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           REGISTERS_26_10_port, QN => n10928);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           REGISTERS_26_9_port, QN => n10414);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           REGISTERS_26_8_port, QN => n10415);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           REGISTERS_26_7_port, QN => n10678);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           REGISTERS_26_6_port, QN => n10416);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           REGISTERS_26_5_port, QN => n10679);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           REGISTERS_26_4_port, QN => n10680);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           REGISTERS_26_3_port, QN => n10929);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           REGISTERS_26_2_port, QN => n10417);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           REGISTERS_26_1_port, QN => n10418);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           REGISTERS_26_0_port, QN => n10681);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           REGISTERS_27_31_port, QN => n10204);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           REGISTERS_27_30_port, QN => n10682);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           REGISTERS_27_29_port, QN => n10683);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           REGISTERS_27_28_port, QN => n10684);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           REGISTERS_27_27_port, QN => n10930);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           REGISTERS_27_26_port, QN => n10419);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           REGISTERS_27_25_port, QN => n10685);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           REGISTERS_27_24_port, QN => n10686);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           REGISTERS_27_23_port, QN => n10420);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           REGISTERS_27_22_port, QN => n10421);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           REGISTERS_27_21_port, QN => n10422);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           REGISTERS_27_20_port, QN => n10687);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           REGISTERS_27_19_port, QN => n10423);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           REGISTERS_27_18_port, QN => n10424);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           REGISTERS_27_17_port, QN => n10425);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           REGISTERS_27_16_port, QN => n10688);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           REGISTERS_27_15_port, QN => n10426);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           REGISTERS_27_14_port, QN => n10689);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           REGISTERS_27_13_port, QN => n10427);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           REGISTERS_27_12_port, QN => n10690);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           REGISTERS_27_11_port, QN => n10691);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           REGISTERS_27_10_port, QN => n10692);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           REGISTERS_27_9_port, QN => n10693);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           REGISTERS_27_8_port, QN => n10428);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           REGISTERS_27_7_port, QN => n10429);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           REGISTERS_27_6_port, QN => n10694);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           REGISTERS_27_5_port, QN => n10695);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           REGISTERS_27_4_port, QN => n10696);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           REGISTERS_27_3_port, QN => n10697);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           REGISTERS_27_2_port, QN => n10698);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           REGISTERS_27_1_port, QN => n10430);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           REGISTERS_27_0_port, QN => n10699);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           REGISTERS_28_31_port, QN => n10451);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           REGISTERS_28_30_port, QN => n11190);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           REGISTERS_28_29_port, QN => n10931);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           REGISTERS_28_28_port, QN => n11191);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           REGISTERS_28_27_port, QN => n11192);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           REGISTERS_28_26_port, QN => n10932);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           REGISTERS_28_25_port, QN => n10933);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           REGISTERS_28_24_port, QN => n10934);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           REGISTERS_28_23_port, QN => n10935);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           REGISTERS_28_22_port, QN => n11193);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           REGISTERS_28_21_port, QN => n10936);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           REGISTERS_28_20_port, QN => n10937);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           REGISTERS_28_19_port, QN => n11194);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           REGISTERS_28_18_port, QN => n10938);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           REGISTERS_28_17_port, QN => n10700);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           REGISTERS_28_16_port, QN => n10939);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           REGISTERS_28_15_port, QN => n10940);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           REGISTERS_28_14_port, QN => n11195);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           REGISTERS_28_13_port, QN => n10941);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           REGISTERS_28_12_port, QN => n10942);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           REGISTERS_28_11_port, QN => n10943);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           REGISTERS_28_10_port, QN => n10944);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           REGISTERS_28_9_port, QN => n10945);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           REGISTERS_28_8_port, QN => n10946);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           REGISTERS_28_7_port, QN => n10947);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           REGISTERS_28_6_port, QN => n10948);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           REGISTERS_28_5_port, QN => n11196);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           REGISTERS_28_4_port, QN => n10949);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           REGISTERS_28_3_port, QN => n10950);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           REGISTERS_28_2_port, QN => n10951);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           REGISTERS_28_1_port, QN => n10952);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           REGISTERS_28_0_port, QN => n11197);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           REGISTERS_29_31_port, QN => n10452);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           REGISTERS_29_30_port, QN => n10701);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           REGISTERS_29_29_port, QN => n10431);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           REGISTERS_29_28_port, QN => n10702);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           REGISTERS_29_27_port, QN => n10432);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           REGISTERS_29_26_port, QN => n10433);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           REGISTERS_29_25_port, QN => n11198);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           REGISTERS_29_24_port, QN => n10953);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           REGISTERS_29_23_port, QN => n10954);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           REGISTERS_29_22_port, QN => n10955);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           REGISTERS_29_21_port, QN => n10956);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           REGISTERS_29_20_port, QN => n11199);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           REGISTERS_29_19_port, QN => n10957);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           REGISTERS_29_18_port, QN => n10958);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           REGISTERS_29_17_port, QN => n10959);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           REGISTERS_29_16_port, QN => n10960);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           REGISTERS_29_15_port, QN => n11200);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           REGISTERS_29_14_port, QN => n10703);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           REGISTERS_29_13_port, QN => n11201);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           REGISTERS_29_12_port, QN => n10961);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           REGISTERS_29_11_port, QN => n10434);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           REGISTERS_29_10_port, QN => n10435);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           REGISTERS_29_9_port, QN => n11202);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           REGISTERS_29_8_port, QN => n10704);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           REGISTERS_29_7_port, QN => n10962);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           REGISTERS_29_6_port, QN => n11203);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           REGISTERS_29_5_port, QN => n10963);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           REGISTERS_29_4_port, QN => n10436);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           REGISTERS_29_3_port, QN => n10964);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           REGISTERS_29_2_port, QN => n11204);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           REGISTERS_29_1_port, QN => n10705);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           REGISTERS_29_0_port, QN => n10965);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           REGISTERS_30_31_port, QN => n10721);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           REGISTERS_30_30_port, QN => n11205);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           REGISTERS_30_29_port, QN => n10966);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           REGISTERS_30_28_port, QN => n10967);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           REGISTERS_30_27_port, QN => n10968);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           REGISTERS_30_26_port, QN => n11206);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           REGISTERS_30_25_port, QN => n10969);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           REGISTERS_30_24_port, QN => n10970);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           REGISTERS_30_23_port, QN => n10971);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           REGISTERS_30_22_port, QN => n11207);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           REGISTERS_30_21_port, QN => n11208);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           REGISTERS_30_20_port, QN => n11209);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           REGISTERS_30_19_port, QN => n11210);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           REGISTERS_30_18_port, QN => n10972);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           REGISTERS_30_17_port, QN => n11211);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           REGISTERS_30_16_port, QN => n10973);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           REGISTERS_30_15_port, QN => n11212);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           REGISTERS_30_14_port, QN => n10974);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           REGISTERS_30_13_port, QN => n10975);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           REGISTERS_30_12_port, QN => n11213);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           REGISTERS_30_11_port, QN => n11214);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           REGISTERS_30_10_port, QN => n10976);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           REGISTERS_30_9_port, QN => n10977);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           REGISTERS_30_8_port, QN => n11215);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           REGISTERS_30_7_port, QN => n11216);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           REGISTERS_30_6_port, QN => n10978);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           REGISTERS_30_5_port, QN => n10979);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1179, CK => CLK, Q => 
                           REGISTERS_30_4_port, QN => n10980);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1178, CK => CLK, Q => 
                           REGISTERS_30_3_port, QN => n11217);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1177, CK => CLK, Q => 
                           REGISTERS_30_2_port, QN => n11218);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1176, CK => CLK, Q => 
                           REGISTERS_30_1_port, QN => n10981);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1175, CK => CLK, Q => 
                           REGISTERS_30_0_port, QN => n11219);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1174, CK => CLK, Q => 
                           REGISTERS_31_31_port, QN => n10205);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1173, CK => CLK, Q => 
                           REGISTERS_31_30_port, QN => n10437);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1172, CK => CLK, Q => 
                           REGISTERS_31_29_port, QN => n10982);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1171, CK => CLK, Q => 
                           REGISTERS_31_28_port, QN => n10706);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1170, CK => CLK, Q => 
                           REGISTERS_31_27_port, QN => n10707);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1169, CK => CLK, Q => 
                           REGISTERS_31_26_port, QN => n10438);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1168, CK => CLK, Q => 
                           REGISTERS_31_25_port, QN => n10439);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1167, CK => CLK, Q => 
                           REGISTERS_31_24_port, QN => n10983);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1166, CK => CLK, Q => 
                           REGISTERS_31_23_port, QN => n11220);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1165, CK => CLK, Q => 
                           REGISTERS_31_22_port, QN => n10708);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1164, CK => CLK, Q => 
                           REGISTERS_31_21_port, QN => n10709);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1163, CK => CLK, Q => 
                           REGISTERS_31_20_port, QN => n10984);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1162, CK => CLK, Q => 
                           REGISTERS_31_19_port, QN => n10440);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1161, CK => CLK, Q => 
                           REGISTERS_31_18_port, QN => n10441);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1160, CK => CLK, Q => 
                           REGISTERS_31_17_port, QN => n11221);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1159, CK => CLK, Q => 
                           REGISTERS_31_16_port, QN => n11222);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1158, CK => CLK, Q => 
                           REGISTERS_31_15_port, QN => n10710);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1157, CK => CLK, Q => 
                           REGISTERS_31_14_port, QN => n10442);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1156, CK => CLK, Q => 
                           REGISTERS_31_13_port, QN => n10711);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1155, CK => CLK, Q => 
                           REGISTERS_31_12_port, QN => n10443);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1154, CK => CLK, Q => 
                           REGISTERS_31_11_port, QN => n10712);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1153, CK => CLK, Q => 
                           REGISTERS_31_10_port, QN => n10713);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1152, CK => CLK, Q => 
                           REGISTERS_31_9_port, QN => n10714);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1151, CK => CLK, Q => 
                           REGISTERS_31_8_port, QN => n10985);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1150, CK => CLK, Q => 
                           REGISTERS_31_7_port, QN => n11223);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1149, CK => CLK, Q => 
                           REGISTERS_31_6_port, QN => n10715);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1148, CK => CLK, Q => 
                           REGISTERS_31_5_port, QN => n10986);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1147, CK => CLK, Q => 
                           REGISTERS_31_4_port, QN => n10716);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1146, CK => CLK, Q => 
                           REGISTERS_31_3_port, QN => n10444);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1145, CK => CLK, Q => 
                           REGISTERS_31_2_port, QN => n10717);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1144, CK => CLK, Q => 
                           REGISTERS_31_1_port, QN => n11224);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1143, CK => CLK, Q => 
                           REGISTERS_31_0_port, QN => n11225);
   OUT1_reg_31_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT1(31), QN 
                           => n_1349);
   OUT1_reg_30_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT1(30), QN 
                           => n_1350);
   OUT1_reg_29_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT1(29), QN 
                           => n_1351);
   OUT1_reg_28_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT1(28), QN 
                           => n_1352);
   OUT1_reg_27_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT1(27), QN 
                           => n_1353);
   OUT1_reg_26_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT1(26), QN 
                           => n_1354);
   OUT1_reg_25_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT1(25), QN 
                           => n_1355);
   OUT1_reg_24_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT1(24), QN 
                           => n_1356);
   OUT1_reg_23_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT1(23), QN 
                           => n_1357);
   OUT1_reg_22_inst : DFF_X1 port map( D => N407, CK => CLK, Q => OUT1(22), QN 
                           => n_1358);
   OUT1_reg_21_inst : DFF_X1 port map( D => N406, CK => CLK, Q => OUT1(21), QN 
                           => n_1359);
   OUT1_reg_20_inst : DFF_X1 port map( D => N405, CK => CLK, Q => OUT1(20), QN 
                           => n_1360);
   OUT1_reg_19_inst : DFF_X1 port map( D => N404, CK => CLK, Q => OUT1(19), QN 
                           => n_1361);
   OUT1_reg_18_inst : DFF_X1 port map( D => N403, CK => CLK, Q => OUT1(18), QN 
                           => n_1362);
   OUT1_reg_17_inst : DFF_X1 port map( D => N402, CK => CLK, Q => OUT1(17), QN 
                           => n_1363);
   OUT1_reg_16_inst : DFF_X1 port map( D => N401, CK => CLK, Q => OUT1(16), QN 
                           => n_1364);
   OUT1_reg_15_inst : DFF_X1 port map( D => N400, CK => CLK, Q => OUT1(15), QN 
                           => n_1365);
   OUT1_reg_14_inst : DFF_X1 port map( D => N399, CK => CLK, Q => OUT1(14), QN 
                           => n_1366);
   OUT1_reg_13_inst : DFF_X1 port map( D => N398, CK => CLK, Q => OUT1(13), QN 
                           => n_1367);
   OUT1_reg_12_inst : DFF_X1 port map( D => N397, CK => CLK, Q => OUT1(12), QN 
                           => n_1368);
   OUT1_reg_11_inst : DFF_X1 port map( D => N396, CK => CLK, Q => OUT1(11), QN 
                           => n_1369);
   OUT1_reg_10_inst : DFF_X1 port map( D => N395, CK => CLK, Q => OUT1(10), QN 
                           => n_1370);
   OUT1_reg_9_inst : DFF_X1 port map( D => N394, CK => CLK, Q => OUT1(9), QN =>
                           n_1371);
   OUT1_reg_8_inst : DFF_X1 port map( D => N393, CK => CLK, Q => OUT1(8), QN =>
                           n_1372);
   OUT1_reg_7_inst : DFF_X1 port map( D => N392, CK => CLK, Q => OUT1(7), QN =>
                           n_1373);
   OUT1_reg_6_inst : DFF_X1 port map( D => N391, CK => CLK, Q => OUT1(6), QN =>
                           n_1374);
   OUT1_reg_5_inst : DFF_X1 port map( D => N390, CK => CLK, Q => OUT1(5), QN =>
                           n_1375);
   OUT1_reg_4_inst : DFF_X1 port map( D => N389, CK => CLK, Q => OUT1(4), QN =>
                           n_1376);
   OUT1_reg_3_inst : DFF_X1 port map( D => N388, CK => CLK, Q => OUT1(3), QN =>
                           n_1377);
   OUT1_reg_2_inst : DFF_X1 port map( D => N387, CK => CLK, Q => OUT1(2), QN =>
                           n_1378);
   OUT1_reg_1_inst : DFF_X1 port map( D => N386, CK => CLK, Q => OUT1(1), QN =>
                           n_1379);
   OUT2_reg_31_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT2(31), QN 
                           => n_1380);
   OUT2_reg_30_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT2(30), QN 
                           => n_1381);
   OUT2_reg_29_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT2(29), QN 
                           => n_1382);
   OUT2_reg_28_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT2(28), QN 
                           => n_1383);
   OUT2_reg_27_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT2(27), QN 
                           => n_1384);
   OUT2_reg_26_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT2(26), QN 
                           => n_1385);
   OUT2_reg_25_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT2(25), QN 
                           => n_1386);
   OUT2_reg_24_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT2(24), QN 
                           => n_1387);
   OUT2_reg_23_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT2(23), QN 
                           => n_1388);
   OUT2_reg_22_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(22), QN 
                           => n_1389);
   OUT2_reg_21_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(21), QN 
                           => n_1390);
   OUT2_reg_20_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(20), QN 
                           => n_1391);
   OUT2_reg_19_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(19), QN 
                           => n_1392);
   OUT2_reg_18_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(18), QN 
                           => n_1393);
   OUT2_reg_17_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(17), QN 
                           => n_1394);
   OUT2_reg_16_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(16), QN 
                           => n_1395);
   OUT2_reg_15_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(15), QN 
                           => n_1396);
   OUT2_reg_14_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(14), QN 
                           => n_1397);
   OUT2_reg_13_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(13), QN 
                           => n_1398);
   OUT2_reg_12_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(12), QN 
                           => n_1399);
   OUT2_reg_11_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(11), QN 
                           => n_1400);
   OUT2_reg_10_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(10), QN 
                           => n_1401);
   OUT2_reg_9_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(9), QN =>
                           n_1402);
   OUT2_reg_8_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(8), QN =>
                           n_1403);
   OUT2_reg_7_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(7), QN =>
                           n_1404);
   OUT2_reg_6_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(6), QN =>
                           n_1405);
   OUT2_reg_5_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(5), QN =>
                           n_1406);
   OUT2_reg_4_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(4), QN =>
                           n_1407);
   OUT2_reg_3_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(3), QN =>
                           n_1408);
   OUT2_reg_2_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(2), QN =>
                           n_1409);
   OUT2_reg_1_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(1), QN =>
                           n_1410);
   OUT2_reg_0_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(0), QN =>
                           n_1411);
   OUT1_reg_0_inst : DFF_X1 port map( D => N385, CK => CLK, Q => OUT1(0), QN =>
                           n_1412);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => 
                           REGISTERS_0_31_port, QN => n10206);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => 
                           REGISTERS_0_30_port, QN => n10207);
   U3 : CLKBUF_X1 port map( A => RESET_BAR, Z => n8448);
   U4 : CLKBUF_X1 port map( A => RESET_BAR, Z => n8449);
   U5 : CLKBUF_X1 port map( A => RESET_BAR, Z => n8450);
   U6 : CLKBUF_X1 port map( A => RESET_BAR, Z => n8451);
   U7 : NAND2_X2 port map( A1 => n8448, A2 => n8625, ZN => n8637);
   U8 : NAND2_X2 port map( A1 => n8448, A2 => n8598, ZN => n8600);
   U9 : NAND2_X2 port map( A1 => n8448, A2 => n8594, ZN => n8596);
   U10 : NAND2_X2 port map( A1 => n8449, A2 => n8590, ZN => n8592);
   U11 : NAND2_X2 port map( A1 => n8451, A2 => n8586, ZN => n8588);
   U12 : NAND2_X2 port map( A1 => n8448, A2 => n8582, ZN => n8584);
   U13 : NAND2_X2 port map( A1 => n8451, A2 => n8573, ZN => n8575);
   U14 : NAND2_X2 port map( A1 => n8451, A2 => n8508, ZN => n8510);
   U15 : NAND2_X2 port map( A1 => n8448, A2 => n8504, ZN => n8506);
   U16 : NAND2_X2 port map( A1 => n8448, A2 => n8501, ZN => n8503);
   U17 : NAND2_X2 port map( A1 => n8451, A2 => n8498, ZN => n8500);
   U18 : NAND2_X2 port map( A1 => n8449, A2 => n8495, ZN => n8497);
   U19 : NAND2_X2 port map( A1 => n8448, A2 => n8488, ZN => n8490);
   U20 : NAND2_X2 port map( A1 => n8448, A2 => n8485, ZN => n8487);
   U21 : NAND2_X2 port map( A1 => n8451, A2 => n8567, ZN => n8569);
   U22 : NAND2_X2 port map( A1 => n8451, A2 => n8562, ZN => n8564);
   U23 : NAND2_X2 port map( A1 => n8448, A2 => n8555, ZN => n8557);
   U24 : NAND2_X2 port map( A1 => n8448, A2 => n8552, ZN => n8554);
   U25 : NAND2_X2 port map( A1 => n8450, A2 => n8539, ZN => n8551);
   U26 : NAND2_X2 port map( A1 => n8449, A2 => n8515, ZN => n8517);
   U27 : NAND2_X2 port map( A1 => n8448, A2 => n8512, ZN => n8514);
   U28 : NAND2_X2 port map( A1 => n8451, A2 => n8482, ZN => n8484);
   U29 : NAND2_X2 port map( A1 => n8448, A2 => n8476, ZN => n8478);
   U30 : NAND2_X2 port map( A1 => n8451, A2 => n8472, ZN => n8474);
   U31 : NAND2_X2 port map( A1 => n8451, A2 => n8468, ZN => n8470);
   U32 : INV_X1 port map( A => ADD_WR(4), ZN => n8571);
   U33 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n8570, ZN => n8507);
   U34 : NOR2_X1 port map( A1 => ADD_WR(4), A2 => n8511, ZN => n8481);
   U35 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(0), A3 => ADD_WR(1), 
                           ZN => n8572);
   U36 : CLKBUF_X1 port map( A => n9419, Z => n9365);
   U37 : CLKBUF_X1 port map( A => n10201, Z => n10148);
   U38 : CLKBUF_X1 port map( A => n8594, Z => n8595);
   U39 : NAND2_X1 port map( A1 => n8449, A2 => n8577, ZN => n8580);
   U40 : NAND2_X1 port map( A1 => n8449, A2 => n8558, ZN => n8561);
   U41 : CLKBUF_X1 port map( A => n8504, Z => n8505);
   U42 : CLKBUF_X1 port map( A => n8544, Z => n8630);
   U43 : CLKBUF_X1 port map( A => n8528, Z => n8614);
   U44 : NAND2_X1 port map( A1 => n8449, A2 => n8491, ZN => n8494);
   U45 : NAND2_X1 port map( A1 => n8450, A2 => n8464, ZN => n8467);
   U46 : NAND2_X1 port map( A1 => n8449, A2 => n8457, ZN => n8460);
   U47 : CLKBUF_X1 port map( A => n8454, Z => n8455);
   U48 : INV_X1 port map( A => ADD_WR(3), ZN => n8452);
   U49 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n8452, ZN => n8511);
   U50 : NAND2_X1 port map( A1 => n8572, A2 => n8481, ZN => n8454);
   U51 : NAND2_X1 port map( A1 => n8449, A2 => n8455, ZN => n8456);
   U52 : CLKBUF_X1 port map( A => n8456, Z => n8453);
   U53 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(31), ZN => n8603);
   U54 : CLKBUF_X1 port map( A => n8603, Z => n8566);
   U55 : OAI22_X1 port map( A1 => n10206, A2 => n8453, B1 => n8566, B2 => n8455
                           , ZN => n2166);
   U56 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(30), ZN => n8518);
   U57 : OAI22_X1 port map( A1 => n10207, A2 => n8456, B1 => n8455, B2 => n8518
                           , ZN => n2165);
   U58 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(29), ZN => n8519);
   U59 : OAI22_X1 port map( A1 => n10722, A2 => n8453, B1 => n8455, B2 => n8519
                           , ZN => n2164);
   U60 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(28), ZN => n8520);
   U61 : OAI22_X1 port map( A1 => n10723, A2 => n8456, B1 => n8455, B2 => n8520
                           , ZN => n2163);
   U62 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(27), ZN => n8521);
   U63 : OAI22_X1 port map( A1 => n10453, A2 => n8453, B1 => n8455, B2 => n8521
                           , ZN => n2162);
   U64 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(26), ZN => n8522);
   U65 : OAI22_X1 port map( A1 => n10724, A2 => n8456, B1 => n8455, B2 => n8522
                           , ZN => n2161);
   U66 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(25), ZN => n8523);
   U67 : OAI22_X1 port map( A1 => n10454, A2 => n8453, B1 => n8455, B2 => n8523
                           , ZN => n2160);
   U68 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(24), ZN => n8524);
   U69 : OAI22_X1 port map( A1 => n10455, A2 => n8456, B1 => n8455, B2 => n8524
                           , ZN => n2159);
   U70 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(23), ZN => n8525);
   U71 : OAI22_X1 port map( A1 => n10456, A2 => n8453, B1 => n8454, B2 => n8525
                           , ZN => n2158);
   U72 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(22), ZN => n8526);
   U73 : OAI22_X1 port map( A1 => n10457, A2 => n8456, B1 => n8454, B2 => n8526
                           , ZN => n2157);
   U74 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(21), ZN => n8527);
   U75 : OAI22_X1 port map( A1 => n10458, A2 => n8456, B1 => n8454, B2 => n8527
                           , ZN => n2156);
   U76 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(20), ZN => n8528);
   U77 : OAI22_X1 port map( A1 => n10208, A2 => n8456, B1 => n8454, B2 => n8528
                           , ZN => n2155);
   U78 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(19), ZN => n8529);
   U79 : OAI22_X1 port map( A1 => n10459, A2 => n8453, B1 => n8454, B2 => n8529
                           , ZN => n2154);
   U80 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(18), ZN => n8530);
   U81 : OAI22_X1 port map( A1 => n10209, A2 => n8453, B1 => n8454, B2 => n8530
                           , ZN => n2153);
   U82 : NAND2_X1 port map( A1 => n8451, A2 => DATAIN(17), ZN => n8531);
   U83 : OAI22_X1 port map( A1 => n10460, A2 => n8453, B1 => n8454, B2 => n8531
                           , ZN => n2152);
   U84 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(16), ZN => n8532);
   U85 : OAI22_X1 port map( A1 => n10725, A2 => n8453, B1 => n8454, B2 => n8532
                           , ZN => n2151);
   U86 : NAND2_X1 port map( A1 => n8451, A2 => DATAIN(15), ZN => n8533);
   U87 : OAI22_X1 port map( A1 => n10461, A2 => n8453, B1 => n8455, B2 => n8533
                           , ZN => n2150);
   U88 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(14), ZN => n8534);
   U89 : OAI22_X1 port map( A1 => n10462, A2 => n8453, B1 => n8454, B2 => n8534
                           , ZN => n2149);
   U90 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(13), ZN => n8535);
   U91 : OAI22_X1 port map( A1 => n10210, A2 => n8453, B1 => n8455, B2 => n8535
                           , ZN => n2148);
   U92 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(12), ZN => n8536);
   U93 : OAI22_X1 port map( A1 => n10463, A2 => n8453, B1 => n8454, B2 => n8536
                           , ZN => n2147);
   U94 : NAND2_X1 port map( A1 => n8451, A2 => DATAIN(11), ZN => n8537);
   U95 : OAI22_X1 port map( A1 => n10211, A2 => n8453, B1 => n8454, B2 => n8537
                           , ZN => n2146);
   U96 : NAND2_X1 port map( A1 => n8449, A2 => DATAIN(10), ZN => n8538);
   U97 : OAI22_X1 port map( A1 => n10464, A2 => n8453, B1 => n8454, B2 => n8538
                           , ZN => n2145);
   U98 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(9), ZN => n8540);
   U99 : OAI22_X1 port map( A1 => n10465, A2 => n8453, B1 => n8455, B2 => n8540
                           , ZN => n2144);
   U100 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(8), ZN => n8541);
   U101 : OAI22_X1 port map( A1 => n10466, A2 => n8453, B1 => n8454, B2 => 
                           n8541, ZN => n2143);
   U102 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(7), ZN => n8542);
   U103 : OAI22_X1 port map( A1 => n10987, A2 => n8456, B1 => n8455, B2 => 
                           n8542, ZN => n2142);
   U104 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(6), ZN => n8543);
   U105 : OAI22_X1 port map( A1 => n10212, A2 => n8456, B1 => n8454, B2 => 
                           n8543, ZN => n2141);
   U106 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(5), ZN => n8544);
   U107 : OAI22_X1 port map( A1 => n10467, A2 => n8456, B1 => n8455, B2 => 
                           n8544, ZN => n2140);
   U108 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(4), ZN => n8545);
   U109 : OAI22_X1 port map( A1 => n10468, A2 => n8456, B1 => n8454, B2 => 
                           n8545, ZN => n2139);
   U110 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(3), ZN => n8546);
   U111 : OAI22_X1 port map( A1 => n10213, A2 => n8456, B1 => n8455, B2 => 
                           n8546, ZN => n2138);
   U112 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(2), ZN => n8547);
   U113 : OAI22_X1 port map( A1 => n10726, A2 => n8456, B1 => n8454, B2 => 
                           n8547, ZN => n2137);
   U114 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(1), ZN => n8548);
   U115 : OAI22_X1 port map( A1 => n10469, A2 => n8456, B1 => n8455, B2 => 
                           n8548, ZN => n2136);
   U116 : NAND2_X1 port map( A1 => n8450, A2 => DATAIN(0), ZN => n8550);
   U117 : OAI22_X1 port map( A1 => n10470, A2 => n8456, B1 => n8455, B2 => 
                           n8550, ZN => n2135);
   U118 : INV_X1 port map( A => ADD_WR(0), ZN => n8471);
   U119 : NOR3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), A3 => n8471, ZN 
                           => n8576);
   U120 : NAND2_X1 port map( A1 => n8481, A2 => n8576, ZN => n8457);
   U121 : CLKBUF_X1 port map( A => n8460, Z => n8458);
   U122 : CLKBUF_X1 port map( A => n8457, Z => n8459);
   U123 : OAI22_X1 port map( A1 => n10471, A2 => n8458, B1 => n8603, B2 => 
                           n8459, ZN => n2134);
   U124 : OAI22_X1 port map( A1 => n10472, A2 => n8460, B1 => n8518, B2 => 
                           n8457, ZN => n2133);
   U125 : OAI22_X1 port map( A1 => n10214, A2 => n8458, B1 => n8519, B2 => 
                           n8459, ZN => n2132);
   U126 : OAI22_X1 port map( A1 => n10473, A2 => n8460, B1 => n8520, B2 => 
                           n8457, ZN => n2131);
   U127 : OAI22_X1 port map( A1 => n10215, A2 => n8458, B1 => n8521, B2 => 
                           n8459, ZN => n2130);
   U128 : OAI22_X1 port map( A1 => n10216, A2 => n8460, B1 => n8522, B2 => 
                           n8457, ZN => n2129);
   U129 : OAI22_X1 port map( A1 => n10988, A2 => n8458, B1 => n8523, B2 => 
                           n8459, ZN => n2128);
   U130 : OAI22_X1 port map( A1 => n10727, A2 => n8460, B1 => n8524, B2 => 
                           n8457, ZN => n2127);
   U131 : OAI22_X1 port map( A1 => n10728, A2 => n8458, B1 => n8525, B2 => 
                           n8459, ZN => n2126);
   U132 : OAI22_X1 port map( A1 => n10217, A2 => n8460, B1 => n8526, B2 => 
                           n8457, ZN => n2125);
   U133 : OAI22_X1 port map( A1 => n10218, A2 => n8460, B1 => n8527, B2 => 
                           n8457, ZN => n2124);
   U134 : OAI22_X1 port map( A1 => n10474, A2 => n8460, B1 => n8528, B2 => 
                           n8459, ZN => n2123);
   U135 : OAI22_X1 port map( A1 => n10219, A2 => n8458, B1 => n8529, B2 => 
                           n8457, ZN => n2122);
   U136 : OAI22_X1 port map( A1 => n10989, A2 => n8458, B1 => n8530, B2 => 
                           n8459, ZN => n2121);
   U137 : OAI22_X1 port map( A1 => n10990, A2 => n8458, B1 => n8531, B2 => 
                           n8457, ZN => n2120);
   U138 : OAI22_X1 port map( A1 => n10220, A2 => n8458, B1 => n8532, B2 => 
                           n8459, ZN => n2119);
   U139 : OAI22_X1 port map( A1 => n10221, A2 => n8458, B1 => n8533, B2 => 
                           n8457, ZN => n2118);
   U140 : OAI22_X1 port map( A1 => n10475, A2 => n8458, B1 => n8534, B2 => 
                           n8457, ZN => n2117);
   U141 : OAI22_X1 port map( A1 => n10476, A2 => n8458, B1 => n8535, B2 => 
                           n8457, ZN => n2116);
   U142 : OAI22_X1 port map( A1 => n10222, A2 => n8458, B1 => n8536, B2 => 
                           n8457, ZN => n2115);
   U143 : OAI22_X1 port map( A1 => n10477, A2 => n8458, B1 => n8537, B2 => 
                           n8457, ZN => n2114);
   U144 : OAI22_X1 port map( A1 => n10478, A2 => n8458, B1 => n8538, B2 => 
                           n8457, ZN => n2113);
   U145 : OAI22_X1 port map( A1 => n10991, A2 => n8458, B1 => n8540, B2 => 
                           n8457, ZN => n2112);
   U146 : OAI22_X1 port map( A1 => n10729, A2 => n8458, B1 => n8541, B2 => 
                           n8459, ZN => n2111);
   U147 : OAI22_X1 port map( A1 => n10223, A2 => n8460, B1 => n8542, B2 => 
                           n8459, ZN => n2110);
   U148 : OAI22_X1 port map( A1 => n10479, A2 => n8460, B1 => n8543, B2 => 
                           n8459, ZN => n2109);
   U149 : OAI22_X1 port map( A1 => n10992, A2 => n8460, B1 => n8544, B2 => 
                           n8459, ZN => n2108);
   U150 : OAI22_X1 port map( A1 => n10730, A2 => n8460, B1 => n8545, B2 => 
                           n8459, ZN => n2107);
   U151 : OAI22_X1 port map( A1 => n10480, A2 => n8460, B1 => n8546, B2 => 
                           n8459, ZN => n2106);
   U152 : OAI22_X1 port map( A1 => n10481, A2 => n8460, B1 => n8547, B2 => 
                           n8459, ZN => n2105);
   U153 : OAI22_X1 port map( A1 => n10993, A2 => n8460, B1 => n8548, B2 => 
                           n8459, ZN => n2104);
   U154 : OAI22_X1 port map( A1 => n10224, A2 => n8460, B1 => n8550, B2 => 
                           n8459, ZN => n2103);
   U155 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n8471, ZN => n8475);
   U156 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n8475, ZN => n8581);
   U157 : NAND2_X1 port map( A1 => n8481, A2 => n8581, ZN => n8461);
   U158 : NAND2_X2 port map( A1 => n8448, A2 => n8461, ZN => n8463);
   U159 : CLKBUF_X1 port map( A => n8461, Z => n8462);
   U160 : OAI22_X1 port map( A1 => n10482, A2 => n8463, B1 => n8566, B2 => 
                           n8462, ZN => n2102);
   U161 : OAI22_X1 port map( A1 => n10225, A2 => n8463, B1 => n8518, B2 => 
                           n8461, ZN => n2101);
   U162 : OAI22_X1 port map( A1 => n10483, A2 => n8463, B1 => n8519, B2 => 
                           n8462, ZN => n2100);
   U163 : OAI22_X1 port map( A1 => n10226, A2 => n8463, B1 => n8520, B2 => 
                           n8461, ZN => n2099);
   U164 : OAI22_X1 port map( A1 => n10484, A2 => n8463, B1 => n8521, B2 => 
                           n8462, ZN => n2098);
   U165 : OAI22_X1 port map( A1 => n10227, A2 => n8463, B1 => n8522, B2 => 
                           n8461, ZN => n2097);
   U166 : OAI22_X1 port map( A1 => n10485, A2 => n8463, B1 => n8523, B2 => 
                           n8462, ZN => n2096);
   U167 : OAI22_X1 port map( A1 => n10486, A2 => n8463, B1 => n8524, B2 => 
                           n8461, ZN => n2095);
   U168 : OAI22_X1 port map( A1 => n10228, A2 => n8463, B1 => n8525, B2 => 
                           n8462, ZN => n2094);
   U169 : OAI22_X1 port map( A1 => n10229, A2 => n8463, B1 => n8526, B2 => 
                           n8461, ZN => n2093);
   U170 : OAI22_X1 port map( A1 => n10230, A2 => n8463, B1 => n8527, B2 => 
                           n8461, ZN => n2092);
   U171 : OAI22_X1 port map( A1 => n10487, A2 => n8463, B1 => n8528, B2 => 
                           n8462, ZN => n2091);
   U172 : OAI22_X1 port map( A1 => n10231, A2 => n8463, B1 => n8529, B2 => 
                           n8461, ZN => n2090);
   U173 : OAI22_X1 port map( A1 => n10232, A2 => n8463, B1 => n8530, B2 => 
                           n8462, ZN => n2089);
   U174 : OAI22_X1 port map( A1 => n10233, A2 => n8463, B1 => n8531, B2 => 
                           n8461, ZN => n2088);
   U175 : OAI22_X1 port map( A1 => n10488, A2 => n8463, B1 => n8532, B2 => 
                           n8462, ZN => n2087);
   U176 : OAI22_X1 port map( A1 => n10234, A2 => n8463, B1 => n8533, B2 => 
                           n8461, ZN => n2086);
   U177 : OAI22_X1 port map( A1 => n10235, A2 => n8463, B1 => n8534, B2 => 
                           n8461, ZN => n2085);
   U178 : OAI22_X1 port map( A1 => n10489, A2 => n8463, B1 => n8535, B2 => 
                           n8461, ZN => n2084);
   U179 : OAI22_X1 port map( A1 => n10490, A2 => n8463, B1 => n8536, B2 => 
                           n8461, ZN => n2083);
   U180 : OAI22_X1 port map( A1 => n10491, A2 => n8463, B1 => n8537, B2 => 
                           n8461, ZN => n2082);
   U181 : OAI22_X1 port map( A1 => n10492, A2 => n8463, B1 => n8538, B2 => 
                           n8461, ZN => n2081);
   U182 : OAI22_X1 port map( A1 => n10236, A2 => n8463, B1 => n8540, B2 => 
                           n8461, ZN => n2080);
   U183 : OAI22_X1 port map( A1 => n10237, A2 => n8463, B1 => n8541, B2 => 
                           n8462, ZN => n2079);
   U184 : OAI22_X1 port map( A1 => n10493, A2 => n8463, B1 => n8542, B2 => 
                           n8462, ZN => n2078);
   U185 : OAI22_X1 port map( A1 => n10238, A2 => n8463, B1 => n8543, B2 => 
                           n8462, ZN => n2077);
   U186 : OAI22_X1 port map( A1 => n10239, A2 => n8463, B1 => n8544, B2 => 
                           n8462, ZN => n2076);
   U187 : OAI22_X1 port map( A1 => n10240, A2 => n8463, B1 => n8545, B2 => 
                           n8462, ZN => n2075);
   U188 : OAI22_X1 port map( A1 => n10494, A2 => n8463, B1 => n8546, B2 => 
                           n8462, ZN => n2074);
   U189 : OAI22_X1 port map( A1 => n10241, A2 => n8463, B1 => n8547, B2 => 
                           n8462, ZN => n2073);
   U190 : OAI22_X1 port map( A1 => n10242, A2 => n8463, B1 => n8548, B2 => 
                           n8462, ZN => n2072);
   U191 : OAI22_X1 port map( A1 => n10495, A2 => n8463, B1 => n8550, B2 => 
                           n8462, ZN => n2071);
   U192 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n8479);
   U193 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => n8479, ZN => n8585);
   U194 : NAND2_X1 port map( A1 => n8481, A2 => n8585, ZN => n8464);
   U195 : CLKBUF_X1 port map( A => n8467, Z => n8465);
   U196 : CLKBUF_X1 port map( A => n8464, Z => n8466);
   U197 : OAI22_X1 port map( A1 => n10731, A2 => n8465, B1 => n8603, B2 => 
                           n8466, ZN => n2070);
   U198 : OAI22_X1 port map( A1 => n10994, A2 => n8467, B1 => n8518, B2 => 
                           n8464, ZN => n2069);
   U199 : OAI22_X1 port map( A1 => n10995, A2 => n8465, B1 => n8519, B2 => 
                           n8466, ZN => n2068);
   U200 : OAI22_X1 port map( A1 => n10732, A2 => n8467, B1 => n8520, B2 => 
                           n8464, ZN => n2067);
   U201 : OAI22_X1 port map( A1 => n10243, A2 => n8465, B1 => n8521, B2 => 
                           n8466, ZN => n2066);
   U202 : OAI22_X1 port map( A1 => n10496, A2 => n8467, B1 => n8522, B2 => 
                           n8464, ZN => n2065);
   U203 : OAI22_X1 port map( A1 => n10244, A2 => n8465, B1 => n8523, B2 => 
                           n8466, ZN => n2064);
   U204 : OAI22_X1 port map( A1 => n10497, A2 => n8467, B1 => n8524, B2 => 
                           n8464, ZN => n2063);
   U205 : OAI22_X1 port map( A1 => n10733, A2 => n8465, B1 => n8525, B2 => 
                           n8466, ZN => n2062);
   U206 : OAI22_X1 port map( A1 => n10498, A2 => n8467, B1 => n8526, B2 => 
                           n8464, ZN => n2061);
   U207 : OAI22_X1 port map( A1 => n10245, A2 => n8467, B1 => n8527, B2 => 
                           n8464, ZN => n2060);
   U208 : OAI22_X1 port map( A1 => n10734, A2 => n8467, B1 => n8528, B2 => 
                           n8466, ZN => n2059);
   U209 : OAI22_X1 port map( A1 => n10246, A2 => n8465, B1 => n8529, B2 => 
                           n8464, ZN => n2058);
   U210 : OAI22_X1 port map( A1 => n10499, A2 => n8465, B1 => n8530, B2 => 
                           n8466, ZN => n2057);
   U211 : OAI22_X1 port map( A1 => n10735, A2 => n8465, B1 => n8531, B2 => 
                           n8464, ZN => n2056);
   U212 : OAI22_X1 port map( A1 => n10500, A2 => n8465, B1 => n8532, B2 => 
                           n8466, ZN => n2055);
   U213 : OAI22_X1 port map( A1 => n10996, A2 => n8465, B1 => n8533, B2 => 
                           n8464, ZN => n2054);
   U214 : OAI22_X1 port map( A1 => n10247, A2 => n8465, B1 => n8534, B2 => 
                           n8464, ZN => n2053);
   U215 : OAI22_X1 port map( A1 => n10997, A2 => n8465, B1 => n8535, B2 => 
                           n8464, ZN => n2052);
   U216 : OAI22_X1 port map( A1 => n10736, A2 => n8465, B1 => n8536, B2 => 
                           n8464, ZN => n2051);
   U217 : OAI22_X1 port map( A1 => n10737, A2 => n8465, B1 => n8537, B2 => 
                           n8464, ZN => n2050);
   U218 : OAI22_X1 port map( A1 => n10738, A2 => n8465, B1 => n8538, B2 => 
                           n8464, ZN => n2049);
   U219 : OAI22_X1 port map( A1 => n10998, A2 => n8465, B1 => n8540, B2 => 
                           n8464, ZN => n2048);
   U220 : OAI22_X1 port map( A1 => n10999, A2 => n8465, B1 => n8541, B2 => 
                           n8466, ZN => n2047);
   U221 : OAI22_X1 port map( A1 => n10248, A2 => n8467, B1 => n8542, B2 => 
                           n8466, ZN => n2046);
   U222 : OAI22_X1 port map( A1 => n10501, A2 => n8467, B1 => n8543, B2 => 
                           n8466, ZN => n2045);
   U223 : OAI22_X1 port map( A1 => n10249, A2 => n8467, B1 => n8544, B2 => 
                           n8466, ZN => n2044);
   U224 : OAI22_X1 port map( A1 => n10502, A2 => n8467, B1 => n8545, B2 => 
                           n8466, ZN => n2043);
   U225 : OAI22_X1 port map( A1 => n10250, A2 => n8467, B1 => n8546, B2 => 
                           n8466, ZN => n2042);
   U226 : OAI22_X1 port map( A1 => n11000, A2 => n8467, B1 => n8547, B2 => 
                           n8466, ZN => n2041);
   U227 : OAI22_X1 port map( A1 => n10251, A2 => n8467, B1 => n8548, B2 => 
                           n8466, ZN => n2040);
   U228 : OAI22_X1 port map( A1 => n10739, A2 => n8467, B1 => n8550, B2 => 
                           n8466, ZN => n2039);
   U229 : INV_X1 port map( A => ADD_WR(2), ZN => n8480);
   U230 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n8480, ZN 
                           => n8589);
   U231 : NAND2_X1 port map( A1 => n8481, A2 => n8589, ZN => n8468);
   U232 : CLKBUF_X1 port map( A => n8468, Z => n8469);
   U233 : OAI22_X1 port map( A1 => n11001, A2 => n8470, B1 => n8566, B2 => 
                           n8469, ZN => n2038);
   U234 : OAI22_X1 port map( A1 => n11002, A2 => n8470, B1 => n8518, B2 => 
                           n8468, ZN => n2037);
   U235 : OAI22_X1 port map( A1 => n11003, A2 => n8470, B1 => n8519, B2 => 
                           n8469, ZN => n2036);
   U236 : OAI22_X1 port map( A1 => n11004, A2 => n8470, B1 => n8520, B2 => 
                           n8468, ZN => n2035);
   U237 : OAI22_X1 port map( A1 => n11005, A2 => n8470, B1 => n8521, B2 => 
                           n8469, ZN => n2034);
   U238 : OAI22_X1 port map( A1 => n11006, A2 => n8470, B1 => n8522, B2 => 
                           n8468, ZN => n2033);
   U239 : OAI22_X1 port map( A1 => n11007, A2 => n8470, B1 => n8523, B2 => 
                           n8469, ZN => n2032);
   U240 : OAI22_X1 port map( A1 => n10740, A2 => n8470, B1 => n8524, B2 => 
                           n8468, ZN => n2031);
   U241 : OAI22_X1 port map( A1 => n10741, A2 => n8470, B1 => n8525, B2 => 
                           n8469, ZN => n2030);
   U242 : OAI22_X1 port map( A1 => n10742, A2 => n8470, B1 => n8526, B2 => 
                           n8468, ZN => n2029);
   U243 : OAI22_X1 port map( A1 => n11008, A2 => n8470, B1 => n8527, B2 => 
                           n8468, ZN => n2028);
   U244 : OAI22_X1 port map( A1 => n10743, A2 => n8470, B1 => n8528, B2 => 
                           n8469, ZN => n2027);
   U245 : OAI22_X1 port map( A1 => n10744, A2 => n8470, B1 => n8529, B2 => 
                           n8468, ZN => n2026);
   U246 : OAI22_X1 port map( A1 => n10745, A2 => n8470, B1 => n8530, B2 => 
                           n8469, ZN => n2025);
   U247 : OAI22_X1 port map( A1 => n10503, A2 => n8470, B1 => n8531, B2 => 
                           n8468, ZN => n2024);
   U248 : OAI22_X1 port map( A1 => n11009, A2 => n8470, B1 => n8532, B2 => 
                           n8469, ZN => n2023);
   U249 : OAI22_X1 port map( A1 => n11010, A2 => n8470, B1 => n8533, B2 => 
                           n8468, ZN => n2022);
   U250 : OAI22_X1 port map( A1 => n10746, A2 => n8470, B1 => n8534, B2 => 
                           n8468, ZN => n2021);
   U251 : OAI22_X1 port map( A1 => n11011, A2 => n8470, B1 => n8535, B2 => 
                           n8468, ZN => n2020);
   U252 : OAI22_X1 port map( A1 => n11012, A2 => n8470, B1 => n8536, B2 => 
                           n8468, ZN => n2019);
   U253 : OAI22_X1 port map( A1 => n10747, A2 => n8470, B1 => n8537, B2 => 
                           n8468, ZN => n2018);
   U254 : OAI22_X1 port map( A1 => n10252, A2 => n8470, B1 => n8538, B2 => 
                           n8468, ZN => n2017);
   U255 : OAI22_X1 port map( A1 => n10253, A2 => n8470, B1 => n8540, B2 => 
                           n8468, ZN => n2016);
   U256 : OAI22_X1 port map( A1 => n10504, A2 => n8470, B1 => n8541, B2 => 
                           n8469, ZN => n2015);
   U257 : OAI22_X1 port map( A1 => n11013, A2 => n8470, B1 => n8542, B2 => 
                           n8469, ZN => n2014);
   U258 : OAI22_X1 port map( A1 => n10748, A2 => n8470, B1 => n8543, B2 => 
                           n8469, ZN => n2013);
   U259 : OAI22_X1 port map( A1 => n11014, A2 => n8470, B1 => n8544, B2 => 
                           n8469, ZN => n2012);
   U260 : OAI22_X1 port map( A1 => n10749, A2 => n8470, B1 => n8545, B2 => 
                           n8469, ZN => n2011);
   U261 : OAI22_X1 port map( A1 => n11015, A2 => n8470, B1 => n8546, B2 => 
                           n8469, ZN => n2010);
   U262 : OAI22_X1 port map( A1 => n11016, A2 => n8470, B1 => n8547, B2 => 
                           n8469, ZN => n2009);
   U263 : OAI22_X1 port map( A1 => n10750, A2 => n8470, B1 => n8548, B2 => 
                           n8469, ZN => n2008);
   U264 : OAI22_X1 port map( A1 => n11017, A2 => n8470, B1 => n8550, B2 => 
                           n8469, ZN => n2007);
   U265 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => n8471, A3 => n8480, ZN => 
                           n8593);
   U266 : NAND2_X1 port map( A1 => n8481, A2 => n8593, ZN => n8472);
   U267 : CLKBUF_X1 port map( A => n8472, Z => n8473);
   U268 : OAI22_X1 port map( A1 => n11018, A2 => n8474, B1 => n8603, B2 => 
                           n8473, ZN => n2006);
   U269 : OAI22_X1 port map( A1 => n11019, A2 => n8474, B1 => n8518, B2 => 
                           n8472, ZN => n2005);
   U270 : OAI22_X1 port map( A1 => n10254, A2 => n8474, B1 => n8519, B2 => 
                           n8473, ZN => n2004);
   U271 : OAI22_X1 port map( A1 => n10505, A2 => n8474, B1 => n8520, B2 => 
                           n8472, ZN => n2003);
   U272 : OAI22_X1 port map( A1 => n11020, A2 => n8474, B1 => n8521, B2 => 
                           n8473, ZN => n2002);
   U273 : OAI22_X1 port map( A1 => n11021, A2 => n8474, B1 => n8522, B2 => 
                           n8472, ZN => n2001);
   U274 : OAI22_X1 port map( A1 => n10751, A2 => n8474, B1 => n8523, B2 => 
                           n8473, ZN => n2000);
   U275 : OAI22_X1 port map( A1 => n10255, A2 => n8474, B1 => n8524, B2 => 
                           n8472, ZN => n1999);
   U276 : OAI22_X1 port map( A1 => n10506, A2 => n8474, B1 => n8525, B2 => 
                           n8473, ZN => n1998);
   U277 : OAI22_X1 port map( A1 => n10752, A2 => n8474, B1 => n8526, B2 => 
                           n8472, ZN => n1997);
   U278 : OAI22_X1 port map( A1 => n11022, A2 => n8474, B1 => n8527, B2 => 
                           n8472, ZN => n1996);
   U279 : OAI22_X1 port map( A1 => n11023, A2 => n8474, B1 => n8528, B2 => 
                           n8473, ZN => n1995);
   U280 : OAI22_X1 port map( A1 => n11024, A2 => n8474, B1 => n8529, B2 => 
                           n8472, ZN => n1994);
   U281 : OAI22_X1 port map( A1 => n11025, A2 => n8474, B1 => n8530, B2 => 
                           n8473, ZN => n1993);
   U282 : OAI22_X1 port map( A1 => n10753, A2 => n8474, B1 => n8531, B2 => 
                           n8472, ZN => n1992);
   U283 : OAI22_X1 port map( A1 => n11026, A2 => n8474, B1 => n8532, B2 => 
                           n8473, ZN => n1991);
   U284 : OAI22_X1 port map( A1 => n10754, A2 => n8474, B1 => n8533, B2 => 
                           n8472, ZN => n1990);
   U285 : OAI22_X1 port map( A1 => n11027, A2 => n8474, B1 => n8534, B2 => 
                           n8472, ZN => n1989);
   U286 : OAI22_X1 port map( A1 => n10755, A2 => n8474, B1 => n8535, B2 => 
                           n8472, ZN => n1988);
   U287 : OAI22_X1 port map( A1 => n10256, A2 => n8474, B1 => n8536, B2 => 
                           n8472, ZN => n1987);
   U288 : OAI22_X1 port map( A1 => n11028, A2 => n8474, B1 => n8537, B2 => 
                           n8472, ZN => n1986);
   U289 : OAI22_X1 port map( A1 => n11029, A2 => n8474, B1 => n8538, B2 => 
                           n8472, ZN => n1985);
   U290 : OAI22_X1 port map( A1 => n10756, A2 => n8474, B1 => n8540, B2 => 
                           n8472, ZN => n1984);
   U291 : OAI22_X1 port map( A1 => n10757, A2 => n8474, B1 => n8541, B2 => 
                           n8473, ZN => n1983);
   U292 : OAI22_X1 port map( A1 => n10758, A2 => n8474, B1 => n8542, B2 => 
                           n8473, ZN => n1982);
   U293 : OAI22_X1 port map( A1 => n11030, A2 => n8474, B1 => n8543, B2 => 
                           n8473, ZN => n1981);
   U294 : OAI22_X1 port map( A1 => n10759, A2 => n8474, B1 => n8544, B2 => 
                           n8473, ZN => n1980);
   U295 : OAI22_X1 port map( A1 => n10760, A2 => n8474, B1 => n8545, B2 => 
                           n8473, ZN => n1979);
   U296 : OAI22_X1 port map( A1 => n11031, A2 => n8474, B1 => n8546, B2 => 
                           n8473, ZN => n1978);
   U297 : OAI22_X1 port map( A1 => n10507, A2 => n8474, B1 => n8547, B2 => 
                           n8473, ZN => n1977);
   U298 : OAI22_X1 port map( A1 => n10761, A2 => n8474, B1 => n8548, B2 => 
                           n8473, ZN => n1976);
   U299 : OAI22_X1 port map( A1 => n11032, A2 => n8474, B1 => n8550, B2 => 
                           n8473, ZN => n1975);
   U300 : NOR2_X1 port map( A1 => n8480, A2 => n8475, ZN => n8597);
   U301 : NAND2_X1 port map( A1 => n8481, A2 => n8597, ZN => n8476);
   U302 : CLKBUF_X1 port map( A => n8476, Z => n8477);
   U303 : OAI22_X1 port map( A1 => n10762, A2 => n8478, B1 => n8566, B2 => 
                           n8477, ZN => n1974);
   U304 : OAI22_X1 port map( A1 => n10763, A2 => n8478, B1 => n8518, B2 => 
                           n8476, ZN => n1973);
   U305 : OAI22_X1 port map( A1 => n10764, A2 => n8478, B1 => n8519, B2 => 
                           n8477, ZN => n1972);
   U306 : OAI22_X1 port map( A1 => n11033, A2 => n8478, B1 => n8520, B2 => 
                           n8476, ZN => n1971);
   U307 : OAI22_X1 port map( A1 => n10765, A2 => n8478, B1 => n8521, B2 => 
                           n8477, ZN => n1970);
   U308 : OAI22_X1 port map( A1 => n11034, A2 => n8478, B1 => n8522, B2 => 
                           n8476, ZN => n1969);
   U309 : OAI22_X1 port map( A1 => n10766, A2 => n8478, B1 => n8523, B2 => 
                           n8477, ZN => n1968);
   U310 : OAI22_X1 port map( A1 => n10767, A2 => n8478, B1 => n8524, B2 => 
                           n8476, ZN => n1967);
   U311 : OAI22_X1 port map( A1 => n11035, A2 => n8478, B1 => n8525, B2 => 
                           n8477, ZN => n1966);
   U312 : OAI22_X1 port map( A1 => n11036, A2 => n8478, B1 => n8526, B2 => 
                           n8476, ZN => n1965);
   U313 : OAI22_X1 port map( A1 => n11037, A2 => n8478, B1 => n8527, B2 => 
                           n8476, ZN => n1964);
   U314 : OAI22_X1 port map( A1 => n10768, A2 => n8478, B1 => n8528, B2 => 
                           n8477, ZN => n1963);
   U315 : OAI22_X1 port map( A1 => n11038, A2 => n8478, B1 => n8529, B2 => 
                           n8476, ZN => n1962);
   U316 : OAI22_X1 port map( A1 => n10769, A2 => n8478, B1 => n8530, B2 => 
                           n8477, ZN => n1961);
   U317 : OAI22_X1 port map( A1 => n11039, A2 => n8478, B1 => n8531, B2 => 
                           n8476, ZN => n1960);
   U318 : OAI22_X1 port map( A1 => n10770, A2 => n8478, B1 => n8532, B2 => 
                           n8477, ZN => n1959);
   U319 : OAI22_X1 port map( A1 => n10771, A2 => n8478, B1 => n8533, B2 => 
                           n8476, ZN => n1958);
   U320 : OAI22_X1 port map( A1 => n10772, A2 => n8478, B1 => n8534, B2 => 
                           n8476, ZN => n1957);
   U321 : OAI22_X1 port map( A1 => n10773, A2 => n8478, B1 => n8535, B2 => 
                           n8476, ZN => n1956);
   U322 : OAI22_X1 port map( A1 => n10774, A2 => n8478, B1 => n8536, B2 => 
                           n8476, ZN => n1955);
   U323 : OAI22_X1 port map( A1 => n11040, A2 => n8478, B1 => n8537, B2 => 
                           n8476, ZN => n1954);
   U324 : OAI22_X1 port map( A1 => n10775, A2 => n8478, B1 => n8538, B2 => 
                           n8476, ZN => n1953);
   U325 : OAI22_X1 port map( A1 => n10776, A2 => n8478, B1 => n8540, B2 => 
                           n8476, ZN => n1952);
   U326 : OAI22_X1 port map( A1 => n10777, A2 => n8478, B1 => n8541, B2 => 
                           n8477, ZN => n1951);
   U327 : OAI22_X1 port map( A1 => n11041, A2 => n8478, B1 => n8542, B2 => 
                           n8477, ZN => n1950);
   U328 : OAI22_X1 port map( A1 => n10778, A2 => n8478, B1 => n8543, B2 => 
                           n8477, ZN => n1949);
   U329 : OAI22_X1 port map( A1 => n11042, A2 => n8478, B1 => n8544, B2 => 
                           n8477, ZN => n1948);
   U330 : OAI22_X1 port map( A1 => n11043, A2 => n8478, B1 => n8545, B2 => 
                           n8477, ZN => n1947);
   U331 : OAI22_X1 port map( A1 => n10779, A2 => n8478, B1 => n8546, B2 => 
                           n8477, ZN => n1946);
   U332 : OAI22_X1 port map( A1 => n10780, A2 => n8478, B1 => n8547, B2 => 
                           n8477, ZN => n1945);
   U333 : OAI22_X1 port map( A1 => n11044, A2 => n8478, B1 => n8548, B2 => 
                           n8477, ZN => n1944);
   U334 : OAI22_X1 port map( A1 => n10781, A2 => n8478, B1 => n8550, B2 => 
                           n8477, ZN => n1943);
   U335 : NOR2_X1 port map( A1 => n8480, A2 => n8479, ZN => n8602);
   U336 : NAND2_X1 port map( A1 => n8481, A2 => n8602, ZN => n8482);
   U337 : CLKBUF_X1 port map( A => n8482, Z => n8483);
   U338 : OAI22_X1 port map( A1 => n10257, A2 => n8484, B1 => n8603, B2 => 
                           n8483, ZN => n1942);
   U339 : OAI22_X1 port map( A1 => n10258, A2 => n8484, B1 => n8518, B2 => 
                           n8482, ZN => n1941);
   U340 : OAI22_X1 port map( A1 => n10508, A2 => n8484, B1 => n8519, B2 => 
                           n8483, ZN => n1940);
   U341 : OAI22_X1 port map( A1 => n10259, A2 => n8484, B1 => n8520, B2 => 
                           n8482, ZN => n1939);
   U342 : OAI22_X1 port map( A1 => n10782, A2 => n8484, B1 => n8521, B2 => 
                           n8483, ZN => n1938);
   U343 : OAI22_X1 port map( A1 => n10260, A2 => n8484, B1 => n8522, B2 => 
                           n8482, ZN => n1937);
   U344 : OAI22_X1 port map( A1 => n10261, A2 => n8484, B1 => n8523, B2 => 
                           n8483, ZN => n1936);
   U345 : OAI22_X1 port map( A1 => n11045, A2 => n8484, B1 => n8524, B2 => 
                           n8482, ZN => n1935);
   U346 : OAI22_X1 port map( A1 => n10509, A2 => n8484, B1 => n8525, B2 => 
                           n8483, ZN => n1934);
   U347 : OAI22_X1 port map( A1 => n11046, A2 => n8484, B1 => n8526, B2 => 
                           n8482, ZN => n1933);
   U348 : OAI22_X1 port map( A1 => n10783, A2 => n8484, B1 => n8527, B2 => 
                           n8482, ZN => n1932);
   U349 : OAI22_X1 port map( A1 => n10510, A2 => n8484, B1 => n8528, B2 => 
                           n8483, ZN => n1931);
   U350 : OAI22_X1 port map( A1 => n11047, A2 => n8484, B1 => n8529, B2 => 
                           n8482, ZN => n1930);
   U351 : OAI22_X1 port map( A1 => n10511, A2 => n8484, B1 => n8530, B2 => 
                           n8483, ZN => n1929);
   U352 : OAI22_X1 port map( A1 => n10262, A2 => n8484, B1 => n8531, B2 => 
                           n8482, ZN => n1928);
   U353 : OAI22_X1 port map( A1 => n10263, A2 => n8484, B1 => n8532, B2 => 
                           n8483, ZN => n1927);
   U354 : OAI22_X1 port map( A1 => n10512, A2 => n8484, B1 => n8533, B2 => 
                           n8482, ZN => n1926);
   U355 : OAI22_X1 port map( A1 => n11048, A2 => n8484, B1 => n8534, B2 => 
                           n8482, ZN => n1925);
   U356 : OAI22_X1 port map( A1 => n10264, A2 => n8484, B1 => n8535, B2 => 
                           n8482, ZN => n1924);
   U357 : OAI22_X1 port map( A1 => n11049, A2 => n8484, B1 => n8536, B2 => 
                           n8482, ZN => n1923);
   U358 : OAI22_X1 port map( A1 => n10265, A2 => n8484, B1 => n8537, B2 => 
                           n8482, ZN => n1922);
   U359 : OAI22_X1 port map( A1 => n10784, A2 => n8484, B1 => n8538, B2 => 
                           n8482, ZN => n1921);
   U360 : OAI22_X1 port map( A1 => n10513, A2 => n8484, B1 => n8540, B2 => 
                           n8482, ZN => n1920);
   U361 : OAI22_X1 port map( A1 => n10514, A2 => n8484, B1 => n8541, B2 => 
                           n8483, ZN => n1919);
   U362 : OAI22_X1 port map( A1 => n10266, A2 => n8484, B1 => n8542, B2 => 
                           n8483, ZN => n1918);
   U363 : OAI22_X1 port map( A1 => n11050, A2 => n8484, B1 => n8543, B2 => 
                           n8483, ZN => n1917);
   U364 : OAI22_X1 port map( A1 => n10267, A2 => n8484, B1 => n8544, B2 => 
                           n8483, ZN => n1916);
   U365 : OAI22_X1 port map( A1 => n10515, A2 => n8484, B1 => n8545, B2 => 
                           n8483, ZN => n1915);
   U366 : OAI22_X1 port map( A1 => n10785, A2 => n8484, B1 => n8546, B2 => 
                           n8483, ZN => n1914);
   U367 : OAI22_X1 port map( A1 => n10268, A2 => n8484, B1 => n8547, B2 => 
                           n8483, ZN => n1913);
   U368 : OAI22_X1 port map( A1 => n10516, A2 => n8484, B1 => n8548, B2 => 
                           n8483, ZN => n1912);
   U369 : OAI22_X1 port map( A1 => n10269, A2 => n8484, B1 => n8550, B2 => 
                           n8483, ZN => n1911);
   U370 : NAND3_X1 port map( A1 => ENABLE, A2 => WR, A3 => ADD_WR(3), ZN => 
                           n8570);
   U371 : NAND2_X1 port map( A1 => n8572, A2 => n8507, ZN => n8485);
   U372 : CLKBUF_X1 port map( A => n8485, Z => n8486);
   U373 : OAI22_X1 port map( A1 => n10270, A2 => n8487, B1 => n8566, B2 => 
                           n8486, ZN => n1910);
   U374 : OAI22_X1 port map( A1 => n10517, A2 => n8487, B1 => n8518, B2 => 
                           n8485, ZN => n1909);
   U375 : OAI22_X1 port map( A1 => n10786, A2 => n8487, B1 => n8519, B2 => 
                           n8486, ZN => n1908);
   U376 : OAI22_X1 port map( A1 => n10518, A2 => n8487, B1 => n8520, B2 => 
                           n8485, ZN => n1907);
   U377 : OAI22_X1 port map( A1 => n10787, A2 => n8487, B1 => n8521, B2 => 
                           n8486, ZN => n1906);
   U378 : OAI22_X1 port map( A1 => n10271, A2 => n8487, B1 => n8522, B2 => 
                           n8485, ZN => n1905);
   U379 : OAI22_X1 port map( A1 => n10519, A2 => n8487, B1 => n8523, B2 => 
                           n8486, ZN => n1904);
   U380 : OAI22_X1 port map( A1 => n10520, A2 => n8487, B1 => n8524, B2 => 
                           n8485, ZN => n1903);
   U381 : OAI22_X1 port map( A1 => n10521, A2 => n8487, B1 => n8525, B2 => 
                           n8486, ZN => n1902);
   U382 : OAI22_X1 port map( A1 => n10272, A2 => n8487, B1 => n8526, B2 => 
                           n8485, ZN => n1901);
   U383 : OAI22_X1 port map( A1 => n10788, A2 => n8487, B1 => n8527, B2 => 
                           n8485, ZN => n1900);
   U384 : OAI22_X1 port map( A1 => n11051, A2 => n8487, B1 => n8528, B2 => 
                           n8486, ZN => n1899);
   U385 : OAI22_X1 port map( A1 => n10273, A2 => n8487, B1 => n8529, B2 => 
                           n8485, ZN => n1898);
   U386 : OAI22_X1 port map( A1 => n10522, A2 => n8487, B1 => n8530, B2 => 
                           n8486, ZN => n1897);
   U387 : OAI22_X1 port map( A1 => n10274, A2 => n8487, B1 => n8531, B2 => 
                           n8485, ZN => n1896);
   U388 : OAI22_X1 port map( A1 => n10523, A2 => n8487, B1 => n8532, B2 => 
                           n8486, ZN => n1895);
   U389 : OAI22_X1 port map( A1 => n10275, A2 => n8487, B1 => n8533, B2 => 
                           n8485, ZN => n1894);
   U390 : OAI22_X1 port map( A1 => n10276, A2 => n8487, B1 => n8534, B2 => 
                           n8485, ZN => n1893);
   U391 : OAI22_X1 port map( A1 => n10277, A2 => n8487, B1 => n8535, B2 => 
                           n8485, ZN => n1892);
   U392 : OAI22_X1 port map( A1 => n10278, A2 => n8487, B1 => n8536, B2 => 
                           n8485, ZN => n1891);
   U393 : OAI22_X1 port map( A1 => n10524, A2 => n8487, B1 => n8537, B2 => 
                           n8485, ZN => n1890);
   U394 : OAI22_X1 port map( A1 => n10279, A2 => n8487, B1 => n8538, B2 => 
                           n8485, ZN => n1889);
   U395 : OAI22_X1 port map( A1 => n10525, A2 => n8487, B1 => n8540, B2 => 
                           n8485, ZN => n1888);
   U396 : OAI22_X1 port map( A1 => n10526, A2 => n8487, B1 => n8541, B2 => 
                           n8486, ZN => n1887);
   U397 : OAI22_X1 port map( A1 => n11052, A2 => n8487, B1 => n8542, B2 => 
                           n8486, ZN => n1886);
   U398 : OAI22_X1 port map( A1 => n10280, A2 => n8487, B1 => n8543, B2 => 
                           n8486, ZN => n1885);
   U399 : OAI22_X1 port map( A1 => n10281, A2 => n8487, B1 => n8544, B2 => 
                           n8486, ZN => n1884);
   U400 : OAI22_X1 port map( A1 => n10282, A2 => n8487, B1 => n8545, B2 => 
                           n8486, ZN => n1883);
   U401 : OAI22_X1 port map( A1 => n10527, A2 => n8487, B1 => n8546, B2 => 
                           n8486, ZN => n1882);
   U402 : OAI22_X1 port map( A1 => n10528, A2 => n8487, B1 => n8547, B2 => 
                           n8486, ZN => n1881);
   U403 : OAI22_X1 port map( A1 => n10283, A2 => n8487, B1 => n8548, B2 => 
                           n8486, ZN => n1880);
   U404 : OAI22_X1 port map( A1 => n10284, A2 => n8487, B1 => n8550, B2 => 
                           n8486, ZN => n1879);
   U405 : NAND2_X1 port map( A1 => n8576, A2 => n8507, ZN => n8488);
   U406 : CLKBUF_X1 port map( A => n8488, Z => n8489);
   U407 : OAI22_X1 port map( A1 => n10529, A2 => n8490, B1 => n8603, B2 => 
                           n8489, ZN => n1878);
   U408 : OAI22_X1 port map( A1 => n10530, A2 => n8490, B1 => n8518, B2 => 
                           n8488, ZN => n1877);
   U409 : OAI22_X1 port map( A1 => n10285, A2 => n8490, B1 => n8519, B2 => 
                           n8489, ZN => n1876);
   U410 : OAI22_X1 port map( A1 => n10531, A2 => n8490, B1 => n8520, B2 => 
                           n8488, ZN => n1875);
   U411 : OAI22_X1 port map( A1 => n10532, A2 => n8490, B1 => n8521, B2 => 
                           n8489, ZN => n1874);
   U412 : OAI22_X1 port map( A1 => n10533, A2 => n8490, B1 => n8522, B2 => 
                           n8488, ZN => n1873);
   U413 : OAI22_X1 port map( A1 => n11053, A2 => n8490, B1 => n8523, B2 => 
                           n8489, ZN => n1872);
   U414 : OAI22_X1 port map( A1 => n10286, A2 => n8490, B1 => n8524, B2 => 
                           n8488, ZN => n1871);
   U415 : OAI22_X1 port map( A1 => n10789, A2 => n8490, B1 => n8525, B2 => 
                           n8489, ZN => n1870);
   U416 : OAI22_X1 port map( A1 => n10287, A2 => n8490, B1 => n8526, B2 => 
                           n8488, ZN => n1869);
   U417 : OAI22_X1 port map( A1 => n10288, A2 => n8490, B1 => n8527, B2 => 
                           n8488, ZN => n1868);
   U418 : OAI22_X1 port map( A1 => n10534, A2 => n8490, B1 => n8528, B2 => 
                           n8489, ZN => n1867);
   U419 : OAI22_X1 port map( A1 => n10535, A2 => n8490, B1 => n8529, B2 => 
                           n8488, ZN => n1866);
   U420 : OAI22_X1 port map( A1 => n10536, A2 => n8490, B1 => n8530, B2 => 
                           n8489, ZN => n1865);
   U421 : OAI22_X1 port map( A1 => n10289, A2 => n8490, B1 => n8531, B2 => 
                           n8488, ZN => n1864);
   U422 : OAI22_X1 port map( A1 => n10290, A2 => n8490, B1 => n8532, B2 => 
                           n8489, ZN => n1863);
   U423 : OAI22_X1 port map( A1 => n10537, A2 => n8490, B1 => n8533, B2 => 
                           n8488, ZN => n1862);
   U424 : OAI22_X1 port map( A1 => n10790, A2 => n8490, B1 => n8534, B2 => 
                           n8488, ZN => n1861);
   U425 : OAI22_X1 port map( A1 => n11054, A2 => n8490, B1 => n8535, B2 => 
                           n8488, ZN => n1860);
   U426 : OAI22_X1 port map( A1 => n10291, A2 => n8490, B1 => n8536, B2 => 
                           n8488, ZN => n1859);
   U427 : OAI22_X1 port map( A1 => n10292, A2 => n8490, B1 => n8537, B2 => 
                           n8488, ZN => n1858);
   U428 : OAI22_X1 port map( A1 => n10538, A2 => n8490, B1 => n8538, B2 => 
                           n8488, ZN => n1857);
   U429 : OAI22_X1 port map( A1 => n10791, A2 => n8490, B1 => n8540, B2 => 
                           n8488, ZN => n1856);
   U430 : OAI22_X1 port map( A1 => n10792, A2 => n8490, B1 => n8541, B2 => 
                           n8489, ZN => n1855);
   U431 : OAI22_X1 port map( A1 => n10293, A2 => n8490, B1 => n8542, B2 => 
                           n8489, ZN => n1854);
   U432 : OAI22_X1 port map( A1 => n10294, A2 => n8490, B1 => n8543, B2 => 
                           n8489, ZN => n1853);
   U433 : OAI22_X1 port map( A1 => n10539, A2 => n8490, B1 => n8544, B2 => 
                           n8489, ZN => n1852);
   U434 : OAI22_X1 port map( A1 => n11055, A2 => n8490, B1 => n8545, B2 => 
                           n8489, ZN => n1851);
   U435 : OAI22_X1 port map( A1 => n10540, A2 => n8490, B1 => n8546, B2 => 
                           n8489, ZN => n1850);
   U436 : OAI22_X1 port map( A1 => n10793, A2 => n8490, B1 => n8547, B2 => 
                           n8489, ZN => n1849);
   U437 : OAI22_X1 port map( A1 => n10794, A2 => n8490, B1 => n8548, B2 => 
                           n8489, ZN => n1848);
   U438 : OAI22_X1 port map( A1 => n10795, A2 => n8490, B1 => n8550, B2 => 
                           n8489, ZN => n1847);
   U439 : NAND2_X1 port map( A1 => n8581, A2 => n8507, ZN => n8491);
   U440 : CLKBUF_X1 port map( A => n8494, Z => n8492);
   U441 : CLKBUF_X1 port map( A => n8491, Z => n8493);
   U442 : OAI22_X1 port map( A1 => n10295, A2 => n8492, B1 => n8603, B2 => 
                           n8493, ZN => n1846);
   U443 : OAI22_X1 port map( A1 => n10296, A2 => n8494, B1 => n8518, B2 => 
                           n8491, ZN => n1845);
   U444 : OAI22_X1 port map( A1 => n10297, A2 => n8492, B1 => n8519, B2 => 
                           n8493, ZN => n1844);
   U445 : OAI22_X1 port map( A1 => n10541, A2 => n8494, B1 => n8520, B2 => 
                           n8491, ZN => n1843);
   U446 : OAI22_X1 port map( A1 => n10298, A2 => n8492, B1 => n8521, B2 => 
                           n8493, ZN => n1842);
   U447 : OAI22_X1 port map( A1 => n10542, A2 => n8494, B1 => n8522, B2 => 
                           n8491, ZN => n1841);
   U448 : OAI22_X1 port map( A1 => n10299, A2 => n8492, B1 => n8523, B2 => 
                           n8493, ZN => n1840);
   U449 : OAI22_X1 port map( A1 => n10300, A2 => n8494, B1 => n8524, B2 => 
                           n8491, ZN => n1839);
   U450 : OAI22_X1 port map( A1 => n10543, A2 => n8492, B1 => n8525, B2 => 
                           n8493, ZN => n1838);
   U451 : OAI22_X1 port map( A1 => n10544, A2 => n8494, B1 => n8526, B2 => 
                           n8491, ZN => n1837);
   U452 : OAI22_X1 port map( A1 => n10301, A2 => n8494, B1 => n8527, B2 => 
                           n8491, ZN => n1836);
   U453 : OAI22_X1 port map( A1 => n10545, A2 => n8494, B1 => n8528, B2 => 
                           n8493, ZN => n1835);
   U454 : OAI22_X1 port map( A1 => n10302, A2 => n8492, B1 => n8529, B2 => 
                           n8491, ZN => n1834);
   U455 : OAI22_X1 port map( A1 => n10303, A2 => n8492, B1 => n8530, B2 => 
                           n8493, ZN => n1833);
   U456 : OAI22_X1 port map( A1 => n10546, A2 => n8492, B1 => n8531, B2 => 
                           n8491, ZN => n1832);
   U457 : OAI22_X1 port map( A1 => n10547, A2 => n8492, B1 => n8532, B2 => 
                           n8493, ZN => n1831);
   U458 : OAI22_X1 port map( A1 => n10548, A2 => n8492, B1 => n8533, B2 => 
                           n8491, ZN => n1830);
   U459 : OAI22_X1 port map( A1 => n10549, A2 => n8492, B1 => n8534, B2 => 
                           n8491, ZN => n1829);
   U460 : OAI22_X1 port map( A1 => n10304, A2 => n8492, B1 => n8535, B2 => 
                           n8491, ZN => n1828);
   U461 : OAI22_X1 port map( A1 => n10550, A2 => n8492, B1 => n8536, B2 => 
                           n8491, ZN => n1827);
   U462 : OAI22_X1 port map( A1 => n10551, A2 => n8492, B1 => n8537, B2 => 
                           n8491, ZN => n1826);
   U463 : OAI22_X1 port map( A1 => n10552, A2 => n8492, B1 => n8538, B2 => 
                           n8491, ZN => n1825);
   U464 : OAI22_X1 port map( A1 => n10305, A2 => n8492, B1 => n8540, B2 => 
                           n8491, ZN => n1824);
   U465 : OAI22_X1 port map( A1 => n10553, A2 => n8492, B1 => n8541, B2 => 
                           n8493, ZN => n1823);
   U466 : OAI22_X1 port map( A1 => n10554, A2 => n8494, B1 => n8542, B2 => 
                           n8493, ZN => n1822);
   U467 : OAI22_X1 port map( A1 => n10555, A2 => n8494, B1 => n8543, B2 => 
                           n8493, ZN => n1821);
   U468 : OAI22_X1 port map( A1 => n10556, A2 => n8494, B1 => n8544, B2 => 
                           n8493, ZN => n1820);
   U469 : OAI22_X1 port map( A1 => n10306, A2 => n8494, B1 => n8545, B2 => 
                           n8493, ZN => n1819);
   U470 : OAI22_X1 port map( A1 => n10307, A2 => n8494, B1 => n8546, B2 => 
                           n8493, ZN => n1818);
   U471 : OAI22_X1 port map( A1 => n10557, A2 => n8494, B1 => n8547, B2 => 
                           n8493, ZN => n1817);
   U472 : OAI22_X1 port map( A1 => n10308, A2 => n8494, B1 => n8548, B2 => 
                           n8493, ZN => n1816);
   U473 : OAI22_X1 port map( A1 => n10558, A2 => n8494, B1 => n8550, B2 => 
                           n8493, ZN => n1815);
   U474 : NAND2_X1 port map( A1 => n8585, A2 => n8507, ZN => n8495);
   U475 : CLKBUF_X1 port map( A => n8495, Z => n8496);
   U476 : OAI22_X1 port map( A1 => n10796, A2 => n8497, B1 => n8603, B2 => 
                           n8496, ZN => n1814);
   U477 : CLKBUF_X1 port map( A => n8518, Z => n8604);
   U478 : OAI22_X1 port map( A1 => n10309, A2 => n8497, B1 => n8604, B2 => 
                           n8495, ZN => n1813);
   U479 : CLKBUF_X1 port map( A => n8519, Z => n8605);
   U480 : OAI22_X1 port map( A1 => n10310, A2 => n8497, B1 => n8605, B2 => 
                           n8496, ZN => n1812);
   U481 : CLKBUF_X1 port map( A => n8520, Z => n8606);
   U482 : OAI22_X1 port map( A1 => n10797, A2 => n8497, B1 => n8606, B2 => 
                           n8495, ZN => n1811);
   U483 : CLKBUF_X1 port map( A => n8521, Z => n8607);
   U484 : OAI22_X1 port map( A1 => n11056, A2 => n8497, B1 => n8607, B2 => 
                           n8496, ZN => n1810);
   U485 : CLKBUF_X1 port map( A => n8522, Z => n8608);
   U486 : OAI22_X1 port map( A1 => n10798, A2 => n8497, B1 => n8608, B2 => 
                           n8495, ZN => n1809);
   U487 : CLKBUF_X1 port map( A => n8523, Z => n8609);
   U488 : OAI22_X1 port map( A1 => n10311, A2 => n8497, B1 => n8609, B2 => 
                           n8496, ZN => n1808);
   U489 : CLKBUF_X1 port map( A => n8524, Z => n8610);
   U490 : OAI22_X1 port map( A1 => n10799, A2 => n8497, B1 => n8610, B2 => 
                           n8495, ZN => n1807);
   U491 : CLKBUF_X1 port map( A => n8525, Z => n8611);
   U492 : OAI22_X1 port map( A1 => n11057, A2 => n8497, B1 => n8611, B2 => 
                           n8496, ZN => n1806);
   U493 : CLKBUF_X1 port map( A => n8526, Z => n8612);
   U494 : OAI22_X1 port map( A1 => n10800, A2 => n8497, B1 => n8612, B2 => 
                           n8495, ZN => n1805);
   U495 : CLKBUF_X1 port map( A => n8527, Z => n8613);
   U496 : OAI22_X1 port map( A1 => n10801, A2 => n8497, B1 => n8613, B2 => 
                           n8495, ZN => n1804);
   U497 : OAI22_X1 port map( A1 => n10312, A2 => n8497, B1 => n8614, B2 => 
                           n8496, ZN => n1803);
   U498 : CLKBUF_X1 port map( A => n8529, Z => n8615);
   U499 : OAI22_X1 port map( A1 => n10802, A2 => n8497, B1 => n8615, B2 => 
                           n8495, ZN => n1802);
   U500 : CLKBUF_X1 port map( A => n8530, Z => n8616);
   U501 : OAI22_X1 port map( A1 => n10803, A2 => n8497, B1 => n8616, B2 => 
                           n8496, ZN => n1801);
   U502 : CLKBUF_X1 port map( A => n8531, Z => n8617);
   U503 : OAI22_X1 port map( A1 => n10559, A2 => n8497, B1 => n8617, B2 => 
                           n8495, ZN => n1800);
   U504 : CLKBUF_X1 port map( A => n8532, Z => n8618);
   U505 : OAI22_X1 port map( A1 => n10804, A2 => n8497, B1 => n8618, B2 => 
                           n8496, ZN => n1799);
   U506 : CLKBUF_X1 port map( A => n8533, Z => n8619);
   U507 : OAI22_X1 port map( A1 => n11058, A2 => n8497, B1 => n8619, B2 => 
                           n8495, ZN => n1798);
   U508 : CLKBUF_X1 port map( A => n8534, Z => n8620);
   U509 : OAI22_X1 port map( A1 => n10560, A2 => n8497, B1 => n8620, B2 => 
                           n8495, ZN => n1797);
   U510 : CLKBUF_X1 port map( A => n8535, Z => n8621);
   U511 : OAI22_X1 port map( A1 => n10561, A2 => n8497, B1 => n8621, B2 => 
                           n8495, ZN => n1796);
   U512 : CLKBUF_X1 port map( A => n8536, Z => n8622);
   U513 : OAI22_X1 port map( A1 => n10805, A2 => n8497, B1 => n8622, B2 => 
                           n8495, ZN => n1795);
   U514 : CLKBUF_X1 port map( A => n8537, Z => n8623);
   U515 : OAI22_X1 port map( A1 => n10313, A2 => n8497, B1 => n8623, B2 => 
                           n8495, ZN => n1794);
   U516 : CLKBUF_X1 port map( A => n8538, Z => n8624);
   U517 : OAI22_X1 port map( A1 => n11059, A2 => n8497, B1 => n8624, B2 => 
                           n8495, ZN => n1793);
   U518 : CLKBUF_X1 port map( A => n8540, Z => n8626);
   U519 : OAI22_X1 port map( A1 => n10562, A2 => n8497, B1 => n8626, B2 => 
                           n8495, ZN => n1792);
   U520 : CLKBUF_X1 port map( A => n8541, Z => n8627);
   U521 : OAI22_X1 port map( A1 => n11060, A2 => n8497, B1 => n8627, B2 => 
                           n8496, ZN => n1791);
   U522 : CLKBUF_X1 port map( A => n8542, Z => n8628);
   U523 : OAI22_X1 port map( A1 => n10563, A2 => n8497, B1 => n8628, B2 => 
                           n8496, ZN => n1790);
   U524 : CLKBUF_X1 port map( A => n8543, Z => n8629);
   U525 : OAI22_X1 port map( A1 => n11061, A2 => n8497, B1 => n8629, B2 => 
                           n8496, ZN => n1789);
   U526 : OAI22_X1 port map( A1 => n11062, A2 => n8497, B1 => n8630, B2 => 
                           n8496, ZN => n1788);
   U527 : CLKBUF_X1 port map( A => n8545, Z => n8631);
   U528 : OAI22_X1 port map( A1 => n10564, A2 => n8497, B1 => n8631, B2 => 
                           n8496, ZN => n1787);
   U529 : CLKBUF_X1 port map( A => n8546, Z => n8632);
   U530 : OAI22_X1 port map( A1 => n10806, A2 => n8497, B1 => n8632, B2 => 
                           n8496, ZN => n1786);
   U531 : CLKBUF_X1 port map( A => n8547, Z => n8633);
   U532 : OAI22_X1 port map( A1 => n11063, A2 => n8497, B1 => n8633, B2 => 
                           n8496, ZN => n1785);
   U533 : CLKBUF_X1 port map( A => n8548, Z => n8634);
   U534 : OAI22_X1 port map( A1 => n10565, A2 => n8497, B1 => n8634, B2 => 
                           n8496, ZN => n1784);
   U535 : CLKBUF_X1 port map( A => n8550, Z => n8636);
   U536 : OAI22_X1 port map( A1 => n10314, A2 => n8497, B1 => n8636, B2 => 
                           n8496, ZN => n1783);
   U537 : NAND2_X1 port map( A1 => n8589, A2 => n8507, ZN => n8498);
   U538 : CLKBUF_X1 port map( A => n8498, Z => n8499);
   U539 : OAI22_X1 port map( A1 => n11064, A2 => n8500, B1 => n8566, B2 => 
                           n8499, ZN => n1782);
   U540 : OAI22_X1 port map( A1 => n11065, A2 => n8500, B1 => n8518, B2 => 
                           n8498, ZN => n1781);
   U541 : OAI22_X1 port map( A1 => n11066, A2 => n8500, B1 => n8519, B2 => 
                           n8499, ZN => n1780);
   U542 : OAI22_X1 port map( A1 => n10807, A2 => n8500, B1 => n8520, B2 => 
                           n8498, ZN => n1779);
   U543 : OAI22_X1 port map( A1 => n11067, A2 => n8500, B1 => n8521, B2 => 
                           n8499, ZN => n1778);
   U544 : OAI22_X1 port map( A1 => n11068, A2 => n8500, B1 => n8522, B2 => 
                           n8498, ZN => n1777);
   U545 : OAI22_X1 port map( A1 => n11069, A2 => n8500, B1 => n8523, B2 => 
                           n8499, ZN => n1776);
   U546 : OAI22_X1 port map( A1 => n11070, A2 => n8500, B1 => n8524, B2 => 
                           n8498, ZN => n1775);
   U547 : OAI22_X1 port map( A1 => n10315, A2 => n8500, B1 => n8525, B2 => 
                           n8499, ZN => n1774);
   U548 : OAI22_X1 port map( A1 => n11071, A2 => n8500, B1 => n8526, B2 => 
                           n8498, ZN => n1773);
   U549 : OAI22_X1 port map( A1 => n10566, A2 => n8500, B1 => n8527, B2 => 
                           n8498, ZN => n1772);
   U550 : OAI22_X1 port map( A1 => n10808, A2 => n8500, B1 => n8528, B2 => 
                           n8499, ZN => n1771);
   U551 : OAI22_X1 port map( A1 => n11072, A2 => n8500, B1 => n8529, B2 => 
                           n8498, ZN => n1770);
   U552 : OAI22_X1 port map( A1 => n11073, A2 => n8500, B1 => n8530, B2 => 
                           n8499, ZN => n1769);
   U553 : OAI22_X1 port map( A1 => n11074, A2 => n8500, B1 => n8531, B2 => 
                           n8498, ZN => n1768);
   U554 : OAI22_X1 port map( A1 => n10809, A2 => n8500, B1 => n8532, B2 => 
                           n8499, ZN => n1767);
   U555 : OAI22_X1 port map( A1 => n10567, A2 => n8500, B1 => n8533, B2 => 
                           n8498, ZN => n1766);
   U556 : OAI22_X1 port map( A1 => n10810, A2 => n8500, B1 => n8534, B2 => 
                           n8498, ZN => n1765);
   U557 : OAI22_X1 port map( A1 => n10568, A2 => n8500, B1 => n8535, B2 => 
                           n8498, ZN => n1764);
   U558 : OAI22_X1 port map( A1 => n11075, A2 => n8500, B1 => n8536, B2 => 
                           n8498, ZN => n1763);
   U559 : OAI22_X1 port map( A1 => n11076, A2 => n8500, B1 => n8537, B2 => 
                           n8498, ZN => n1762);
   U560 : OAI22_X1 port map( A1 => n10811, A2 => n8500, B1 => n8538, B2 => 
                           n8498, ZN => n1761);
   U561 : OAI22_X1 port map( A1 => n10812, A2 => n8500, B1 => n8540, B2 => 
                           n8498, ZN => n1760);
   U562 : OAI22_X1 port map( A1 => n10316, A2 => n8500, B1 => n8541, B2 => 
                           n8499, ZN => n1759);
   U563 : OAI22_X1 port map( A1 => n10813, A2 => n8500, B1 => n8542, B2 => 
                           n8499, ZN => n1758);
   U564 : OAI22_X1 port map( A1 => n10814, A2 => n8500, B1 => n8543, B2 => 
                           n8499, ZN => n1757);
   U565 : OAI22_X1 port map( A1 => n10815, A2 => n8500, B1 => n8544, B2 => 
                           n8499, ZN => n1756);
   U566 : OAI22_X1 port map( A1 => n10816, A2 => n8500, B1 => n8545, B2 => 
                           n8499, ZN => n1755);
   U567 : OAI22_X1 port map( A1 => n11077, A2 => n8500, B1 => n8546, B2 => 
                           n8499, ZN => n1754);
   U568 : OAI22_X1 port map( A1 => n11078, A2 => n8500, B1 => n8547, B2 => 
                           n8499, ZN => n1753);
   U569 : OAI22_X1 port map( A1 => n11079, A2 => n8500, B1 => n8548, B2 => 
                           n8499, ZN => n1752);
   U570 : OAI22_X1 port map( A1 => n10569, A2 => n8500, B1 => n8550, B2 => 
                           n8499, ZN => n1751);
   U571 : NAND2_X1 port map( A1 => n8593, A2 => n8507, ZN => n8501);
   U572 : CLKBUF_X1 port map( A => n8501, Z => n8502);
   U573 : OAI22_X1 port map( A1 => n10817, A2 => n8503, B1 => n8566, B2 => 
                           n8502, ZN => n1750);
   U574 : OAI22_X1 port map( A1 => n10818, A2 => n8503, B1 => n8604, B2 => 
                           n8501, ZN => n1749);
   U575 : OAI22_X1 port map( A1 => n10570, A2 => n8503, B1 => n8605, B2 => 
                           n8502, ZN => n1748);
   U576 : OAI22_X1 port map( A1 => n11080, A2 => n8503, B1 => n8606, B2 => 
                           n8501, ZN => n1747);
   U577 : OAI22_X1 port map( A1 => n10317, A2 => n8503, B1 => n8607, B2 => 
                           n8502, ZN => n1746);
   U578 : OAI22_X1 port map( A1 => n10819, A2 => n8503, B1 => n8608, B2 => 
                           n8501, ZN => n1745);
   U579 : OAI22_X1 port map( A1 => n11081, A2 => n8503, B1 => n8609, B2 => 
                           n8502, ZN => n1744);
   U580 : OAI22_X1 port map( A1 => n11082, A2 => n8503, B1 => n8610, B2 => 
                           n8501, ZN => n1743);
   U581 : OAI22_X1 port map( A1 => n11083, A2 => n8503, B1 => n8611, B2 => 
                           n8502, ZN => n1742);
   U582 : OAI22_X1 port map( A1 => n10820, A2 => n8503, B1 => n8612, B2 => 
                           n8501, ZN => n1741);
   U583 : OAI22_X1 port map( A1 => n11084, A2 => n8503, B1 => n8613, B2 => 
                           n8501, ZN => n1740);
   U584 : OAI22_X1 port map( A1 => n11085, A2 => n8503, B1 => n8614, B2 => 
                           n8502, ZN => n1739);
   U585 : OAI22_X1 port map( A1 => n11086, A2 => n8503, B1 => n8615, B2 => 
                           n8501, ZN => n1738);
   U586 : OAI22_X1 port map( A1 => n10821, A2 => n8503, B1 => n8616, B2 => 
                           n8502, ZN => n1737);
   U587 : OAI22_X1 port map( A1 => n11087, A2 => n8503, B1 => n8617, B2 => 
                           n8501, ZN => n1736);
   U588 : OAI22_X1 port map( A1 => n10822, A2 => n8503, B1 => n8618, B2 => 
                           n8502, ZN => n1735);
   U589 : OAI22_X1 port map( A1 => n10823, A2 => n8503, B1 => n8619, B2 => 
                           n8501, ZN => n1734);
   U590 : OAI22_X1 port map( A1 => n10571, A2 => n8503, B1 => n8620, B2 => 
                           n8501, ZN => n1733);
   U591 : OAI22_X1 port map( A1 => n11088, A2 => n8503, B1 => n8621, B2 => 
                           n8501, ZN => n1732);
   U592 : OAI22_X1 port map( A1 => n10572, A2 => n8503, B1 => n8622, B2 => 
                           n8501, ZN => n1731);
   U593 : OAI22_X1 port map( A1 => n11089, A2 => n8503, B1 => n8623, B2 => 
                           n8501, ZN => n1730);
   U594 : OAI22_X1 port map( A1 => n10318, A2 => n8503, B1 => n8624, B2 => 
                           n8501, ZN => n1729);
   U595 : OAI22_X1 port map( A1 => n10319, A2 => n8503, B1 => n8626, B2 => 
                           n8501, ZN => n1728);
   U596 : OAI22_X1 port map( A1 => n10824, A2 => n8503, B1 => n8627, B2 => 
                           n8502, ZN => n1727);
   U597 : OAI22_X1 port map( A1 => n10825, A2 => n8503, B1 => n8628, B2 => 
                           n8502, ZN => n1726);
   U598 : OAI22_X1 port map( A1 => n10826, A2 => n8503, B1 => n8629, B2 => 
                           n8502, ZN => n1725);
   U599 : OAI22_X1 port map( A1 => n10827, A2 => n8503, B1 => n8630, B2 => 
                           n8502, ZN => n1724);
   U600 : OAI22_X1 port map( A1 => n10828, A2 => n8503, B1 => n8631, B2 => 
                           n8502, ZN => n1723);
   U601 : OAI22_X1 port map( A1 => n10573, A2 => n8503, B1 => n8632, B2 => 
                           n8502, ZN => n1722);
   U602 : OAI22_X1 port map( A1 => n10320, A2 => n8503, B1 => n8633, B2 => 
                           n8502, ZN => n1721);
   U603 : OAI22_X1 port map( A1 => n10574, A2 => n8503, B1 => n8634, B2 => 
                           n8502, ZN => n1720);
   U604 : OAI22_X1 port map( A1 => n11090, A2 => n8503, B1 => n8636, B2 => 
                           n8502, ZN => n1719);
   U605 : NAND2_X1 port map( A1 => n8597, A2 => n8507, ZN => n8504);
   U606 : OAI22_X1 port map( A1 => n11091, A2 => n8506, B1 => n8566, B2 => 
                           n8505, ZN => n1718);
   U607 : OAI22_X1 port map( A1 => n11092, A2 => n8506, B1 => n8518, B2 => 
                           n8504, ZN => n1717);
   U608 : OAI22_X1 port map( A1 => n11093, A2 => n8506, B1 => n8519, B2 => 
                           n8505, ZN => n1716);
   U609 : OAI22_X1 port map( A1 => n10829, A2 => n8506, B1 => n8520, B2 => 
                           n8504, ZN => n1715);
   U610 : OAI22_X1 port map( A1 => n10830, A2 => n8506, B1 => n8521, B2 => 
                           n8505, ZN => n1714);
   U611 : OAI22_X1 port map( A1 => n11094, A2 => n8506, B1 => n8522, B2 => 
                           n8504, ZN => n1713);
   U612 : OAI22_X1 port map( A1 => n10831, A2 => n8506, B1 => n8523, B2 => 
                           n8505, ZN => n1712);
   U613 : OAI22_X1 port map( A1 => n10832, A2 => n8506, B1 => n8524, B2 => 
                           n8504, ZN => n1711);
   U614 : OAI22_X1 port map( A1 => n10833, A2 => n8506, B1 => n8525, B2 => 
                           n8505, ZN => n1710);
   U615 : OAI22_X1 port map( A1 => n11095, A2 => n8506, B1 => n8526, B2 => 
                           n8504, ZN => n1709);
   U616 : OAI22_X1 port map( A1 => n11096, A2 => n8506, B1 => n8527, B2 => 
                           n8504, ZN => n1708);
   U617 : OAI22_X1 port map( A1 => n10834, A2 => n8506, B1 => n8528, B2 => 
                           n8505, ZN => n1707);
   U618 : OAI22_X1 port map( A1 => n10835, A2 => n8506, B1 => n8529, B2 => 
                           n8504, ZN => n1706);
   U619 : OAI22_X1 port map( A1 => n11097, A2 => n8506, B1 => n8530, B2 => 
                           n8505, ZN => n1705);
   U620 : OAI22_X1 port map( A1 => n10836, A2 => n8506, B1 => n8531, B2 => 
                           n8504, ZN => n1704);
   U621 : OAI22_X1 port map( A1 => n11098, A2 => n8506, B1 => n8532, B2 => 
                           n8505, ZN => n1703);
   U622 : OAI22_X1 port map( A1 => n10837, A2 => n8506, B1 => n8533, B2 => 
                           n8504, ZN => n1702);
   U623 : OAI22_X1 port map( A1 => n10838, A2 => n8506, B1 => n8534, B2 => 
                           n8504, ZN => n1701);
   U624 : OAI22_X1 port map( A1 => n10839, A2 => n8506, B1 => n8535, B2 => 
                           n8504, ZN => n1700);
   U625 : OAI22_X1 port map( A1 => n11099, A2 => n8506, B1 => n8536, B2 => 
                           n8504, ZN => n1699);
   U626 : OAI22_X1 port map( A1 => n10840, A2 => n8506, B1 => n8537, B2 => 
                           n8504, ZN => n1698);
   U627 : OAI22_X1 port map( A1 => n10841, A2 => n8506, B1 => n8538, B2 => 
                           n8504, ZN => n1697);
   U628 : OAI22_X1 port map( A1 => n11100, A2 => n8506, B1 => n8540, B2 => 
                           n8504, ZN => n1696);
   U629 : OAI22_X1 port map( A1 => n10842, A2 => n8506, B1 => n8541, B2 => 
                           n8505, ZN => n1695);
   U630 : OAI22_X1 port map( A1 => n11101, A2 => n8506, B1 => n8542, B2 => 
                           n8505, ZN => n1694);
   U631 : OAI22_X1 port map( A1 => n11102, A2 => n8506, B1 => n8543, B2 => 
                           n8505, ZN => n1693);
   U632 : OAI22_X1 port map( A1 => n11103, A2 => n8506, B1 => n8544, B2 => 
                           n8505, ZN => n1692);
   U633 : OAI22_X1 port map( A1 => n11104, A2 => n8506, B1 => n8545, B2 => 
                           n8505, ZN => n1691);
   U634 : OAI22_X1 port map( A1 => n10843, A2 => n8506, B1 => n8546, B2 => 
                           n8505, ZN => n1690);
   U635 : OAI22_X1 port map( A1 => n10844, A2 => n8506, B1 => n8547, B2 => 
                           n8505, ZN => n1689);
   U636 : OAI22_X1 port map( A1 => n11105, A2 => n8506, B1 => n8548, B2 => 
                           n8505, ZN => n1688);
   U637 : OAI22_X1 port map( A1 => n11106, A2 => n8506, B1 => n8550, B2 => 
                           n8505, ZN => n1687);
   U638 : NAND2_X1 port map( A1 => n8602, A2 => n8507, ZN => n8508);
   U639 : CLKBUF_X1 port map( A => n8508, Z => n8509);
   U640 : OAI22_X1 port map( A1 => n10575, A2 => n8510, B1 => n8566, B2 => 
                           n8509, ZN => n1686);
   U641 : OAI22_X1 port map( A1 => n10845, A2 => n8510, B1 => n8604, B2 => 
                           n8508, ZN => n1685);
   U642 : OAI22_X1 port map( A1 => n11107, A2 => n8510, B1 => n8605, B2 => 
                           n8509, ZN => n1684);
   U643 : OAI22_X1 port map( A1 => n10321, A2 => n8510, B1 => n8606, B2 => 
                           n8508, ZN => n1683);
   U644 : OAI22_X1 port map( A1 => n10576, A2 => n8510, B1 => n8607, B2 => 
                           n8509, ZN => n1682);
   U645 : OAI22_X1 port map( A1 => n10322, A2 => n8510, B1 => n8608, B2 => 
                           n8508, ZN => n1681);
   U646 : OAI22_X1 port map( A1 => n10323, A2 => n8510, B1 => n8609, B2 => 
                           n8509, ZN => n1680);
   U647 : OAI22_X1 port map( A1 => n10577, A2 => n8510, B1 => n8610, B2 => 
                           n8508, ZN => n1679);
   U648 : OAI22_X1 port map( A1 => n10324, A2 => n8510, B1 => n8611, B2 => 
                           n8509, ZN => n1678);
   U649 : OAI22_X1 port map( A1 => n10578, A2 => n8510, B1 => n8612, B2 => 
                           n8508, ZN => n1677);
   U650 : OAI22_X1 port map( A1 => n10579, A2 => n8510, B1 => n8613, B2 => 
                           n8508, ZN => n1676);
   U651 : OAI22_X1 port map( A1 => n10325, A2 => n8510, B1 => n8614, B2 => 
                           n8509, ZN => n1675);
   U652 : OAI22_X1 port map( A1 => n10580, A2 => n8510, B1 => n8615, B2 => 
                           n8508, ZN => n1674);
   U653 : OAI22_X1 port map( A1 => n10326, A2 => n8510, B1 => n8616, B2 => 
                           n8509, ZN => n1673);
   U654 : OAI22_X1 port map( A1 => n10846, A2 => n8510, B1 => n8617, B2 => 
                           n8508, ZN => n1672);
   U655 : OAI22_X1 port map( A1 => n10581, A2 => n8510, B1 => n8618, B2 => 
                           n8509, ZN => n1671);
   U656 : OAI22_X1 port map( A1 => n10847, A2 => n8510, B1 => n8619, B2 => 
                           n8508, ZN => n1670);
   U657 : OAI22_X1 port map( A1 => n11108, A2 => n8510, B1 => n8620, B2 => 
                           n8508, ZN => n1669);
   U658 : OAI22_X1 port map( A1 => n10848, A2 => n8510, B1 => n8621, B2 => 
                           n8508, ZN => n1668);
   U659 : OAI22_X1 port map( A1 => n10849, A2 => n8510, B1 => n8622, B2 => 
                           n8508, ZN => n1667);
   U660 : OAI22_X1 port map( A1 => n10850, A2 => n8510, B1 => n8623, B2 => 
                           n8508, ZN => n1666);
   U661 : OAI22_X1 port map( A1 => n11109, A2 => n8510, B1 => n8624, B2 => 
                           n8508, ZN => n1665);
   U662 : OAI22_X1 port map( A1 => n11110, A2 => n8510, B1 => n8626, B2 => 
                           n8508, ZN => n1664);
   U663 : OAI22_X1 port map( A1 => n10582, A2 => n8510, B1 => n8627, B2 => 
                           n8509, ZN => n1663);
   U664 : OAI22_X1 port map( A1 => n10327, A2 => n8510, B1 => n8628, B2 => 
                           n8509, ZN => n1662);
   U665 : OAI22_X1 port map( A1 => n10583, A2 => n8510, B1 => n8629, B2 => 
                           n8509, ZN => n1661);
   U666 : OAI22_X1 port map( A1 => n10328, A2 => n8510, B1 => n8630, B2 => 
                           n8509, ZN => n1660);
   U667 : OAI22_X1 port map( A1 => n10584, A2 => n8510, B1 => n8631, B2 => 
                           n8509, ZN => n1659);
   U668 : OAI22_X1 port map( A1 => n10851, A2 => n8510, B1 => n8632, B2 => 
                           n8509, ZN => n1658);
   U669 : OAI22_X1 port map( A1 => n10329, A2 => n8510, B1 => n8633, B2 => 
                           n8509, ZN => n1657);
   U670 : OAI22_X1 port map( A1 => n10852, A2 => n8510, B1 => n8634, B2 => 
                           n8509, ZN => n1656);
   U671 : OAI22_X1 port map( A1 => n10853, A2 => n8510, B1 => n8636, B2 => 
                           n8509, ZN => n1655);
   U672 : NOR2_X1 port map( A1 => n8571, A2 => n8511, ZN => n8565);
   U673 : NAND2_X1 port map( A1 => n8572, A2 => n8565, ZN => n8512);
   U674 : CLKBUF_X1 port map( A => n8512, Z => n8513);
   U675 : OAI22_X1 port map( A1 => n10445, A2 => n8514, B1 => n8566, B2 => 
                           n8513, ZN => n1654);
   U676 : OAI22_X1 port map( A1 => n10330, A2 => n8514, B1 => n8518, B2 => 
                           n8512, ZN => n1653);
   U677 : OAI22_X1 port map( A1 => n10585, A2 => n8514, B1 => n8519, B2 => 
                           n8513, ZN => n1652);
   U678 : OAI22_X1 port map( A1 => n10586, A2 => n8514, B1 => n8520, B2 => 
                           n8512, ZN => n1651);
   U679 : OAI22_X1 port map( A1 => n10587, A2 => n8514, B1 => n8521, B2 => 
                           n8513, ZN => n1650);
   U680 : OAI22_X1 port map( A1 => n10588, A2 => n8514, B1 => n8522, B2 => 
                           n8512, ZN => n1649);
   U681 : OAI22_X1 port map( A1 => n10854, A2 => n8514, B1 => n8523, B2 => 
                           n8513, ZN => n1648);
   U682 : OAI22_X1 port map( A1 => n10589, A2 => n8514, B1 => n8524, B2 => 
                           n8512, ZN => n1647);
   U683 : OAI22_X1 port map( A1 => n10590, A2 => n8514, B1 => n8525, B2 => 
                           n8513, ZN => n1646);
   U684 : OAI22_X1 port map( A1 => n10591, A2 => n8514, B1 => n8526, B2 => 
                           n8512, ZN => n1645);
   U685 : OAI22_X1 port map( A1 => n10592, A2 => n8514, B1 => n8527, B2 => 
                           n8512, ZN => n1644);
   U686 : OAI22_X1 port map( A1 => n10593, A2 => n8514, B1 => n8528, B2 => 
                           n8513, ZN => n1643);
   U687 : OAI22_X1 port map( A1 => n10594, A2 => n8514, B1 => n8529, B2 => 
                           n8512, ZN => n1642);
   U688 : OAI22_X1 port map( A1 => n10595, A2 => n8514, B1 => n8530, B2 => 
                           n8513, ZN => n1641);
   U689 : OAI22_X1 port map( A1 => n10855, A2 => n8514, B1 => n8531, B2 => 
                           n8512, ZN => n1640);
   U690 : OAI22_X1 port map( A1 => n10331, A2 => n8514, B1 => n8532, B2 => 
                           n8513, ZN => n1639);
   U691 : OAI22_X1 port map( A1 => n10332, A2 => n8514, B1 => n8533, B2 => 
                           n8512, ZN => n1638);
   U692 : OAI22_X1 port map( A1 => n10596, A2 => n8514, B1 => n8534, B2 => 
                           n8512, ZN => n1637);
   U693 : OAI22_X1 port map( A1 => n10597, A2 => n8514, B1 => n8535, B2 => 
                           n8512, ZN => n1636);
   U694 : OAI22_X1 port map( A1 => n11111, A2 => n8514, B1 => n8536, B2 => 
                           n8512, ZN => n1635);
   U695 : OAI22_X1 port map( A1 => n10333, A2 => n8514, B1 => n8537, B2 => 
                           n8512, ZN => n1634);
   U696 : OAI22_X1 port map( A1 => n10334, A2 => n8514, B1 => n8538, B2 => 
                           n8512, ZN => n1633);
   U697 : OAI22_X1 port map( A1 => n10598, A2 => n8514, B1 => n8540, B2 => 
                           n8512, ZN => n1632);
   U698 : OAI22_X1 port map( A1 => n10335, A2 => n8514, B1 => n8541, B2 => 
                           n8513, ZN => n1631);
   U699 : OAI22_X1 port map( A1 => n10599, A2 => n8514, B1 => n8542, B2 => 
                           n8513, ZN => n1630);
   U700 : OAI22_X1 port map( A1 => n11112, A2 => n8514, B1 => n8543, B2 => 
                           n8513, ZN => n1629);
   U701 : OAI22_X1 port map( A1 => n11113, A2 => n8514, B1 => n8544, B2 => 
                           n8513, ZN => n1628);
   U702 : OAI22_X1 port map( A1 => n10600, A2 => n8514, B1 => n8545, B2 => 
                           n8513, ZN => n1627);
   U703 : OAI22_X1 port map( A1 => n10336, A2 => n8514, B1 => n8546, B2 => 
                           n8513, ZN => n1626);
   U704 : OAI22_X1 port map( A1 => n11114, A2 => n8514, B1 => n8547, B2 => 
                           n8513, ZN => n1625);
   U705 : OAI22_X1 port map( A1 => n10601, A2 => n8514, B1 => n8548, B2 => 
                           n8513, ZN => n1624);
   U706 : OAI22_X1 port map( A1 => n10337, A2 => n8514, B1 => n8550, B2 => 
                           n8513, ZN => n1623);
   U707 : NAND2_X1 port map( A1 => n8576, A2 => n8565, ZN => n8515);
   U708 : CLKBUF_X1 port map( A => n8515, Z => n8516);
   U709 : OAI22_X1 port map( A1 => n10202, A2 => n8517, B1 => n8566, B2 => 
                           n8516, ZN => n1622);
   U710 : OAI22_X1 port map( A1 => n10338, A2 => n8517, B1 => n8604, B2 => 
                           n8515, ZN => n1621);
   U711 : OAI22_X1 port map( A1 => n10602, A2 => n8517, B1 => n8605, B2 => 
                           n8516, ZN => n1620);
   U712 : OAI22_X1 port map( A1 => n10339, A2 => n8517, B1 => n8606, B2 => 
                           n8515, ZN => n1619);
   U713 : OAI22_X1 port map( A1 => n10603, A2 => n8517, B1 => n8607, B2 => 
                           n8516, ZN => n1618);
   U714 : OAI22_X1 port map( A1 => n10604, A2 => n8517, B1 => n8608, B2 => 
                           n8515, ZN => n1617);
   U715 : OAI22_X1 port map( A1 => n10605, A2 => n8517, B1 => n8609, B2 => 
                           n8516, ZN => n1616);
   U716 : OAI22_X1 port map( A1 => n10340, A2 => n8517, B1 => n8610, B2 => 
                           n8515, ZN => n1615);
   U717 : OAI22_X1 port map( A1 => n10606, A2 => n8517, B1 => n8611, B2 => 
                           n8516, ZN => n1614);
   U718 : OAI22_X1 port map( A1 => n10607, A2 => n8517, B1 => n8612, B2 => 
                           n8515, ZN => n1613);
   U719 : OAI22_X1 port map( A1 => n10341, A2 => n8517, B1 => n8613, B2 => 
                           n8515, ZN => n1612);
   U720 : OAI22_X1 port map( A1 => n10608, A2 => n8517, B1 => n8614, B2 => 
                           n8516, ZN => n1611);
   U721 : OAI22_X1 port map( A1 => n10609, A2 => n8517, B1 => n8615, B2 => 
                           n8515, ZN => n1610);
   U722 : OAI22_X1 port map( A1 => n10610, A2 => n8517, B1 => n8616, B2 => 
                           n8516, ZN => n1609);
   U723 : OAI22_X1 port map( A1 => n10611, A2 => n8517, B1 => n8617, B2 => 
                           n8515, ZN => n1608);
   U724 : OAI22_X1 port map( A1 => n10342, A2 => n8517, B1 => n8618, B2 => 
                           n8516, ZN => n1607);
   U725 : OAI22_X1 port map( A1 => n10612, A2 => n8517, B1 => n8619, B2 => 
                           n8515, ZN => n1606);
   U726 : OAI22_X1 port map( A1 => n10343, A2 => n8517, B1 => n8620, B2 => 
                           n8515, ZN => n1605);
   U727 : OAI22_X1 port map( A1 => n10344, A2 => n8517, B1 => n8621, B2 => 
                           n8515, ZN => n1604);
   U728 : OAI22_X1 port map( A1 => n10345, A2 => n8517, B1 => n8622, B2 => 
                           n8515, ZN => n1603);
   U729 : OAI22_X1 port map( A1 => n10613, A2 => n8517, B1 => n8623, B2 => 
                           n8515, ZN => n1602);
   U730 : OAI22_X1 port map( A1 => n10614, A2 => n8517, B1 => n8624, B2 => 
                           n8515, ZN => n1601);
   U731 : OAI22_X1 port map( A1 => n10615, A2 => n8517, B1 => n8626, B2 => 
                           n8515, ZN => n1600);
   U732 : OAI22_X1 port map( A1 => n10616, A2 => n8517, B1 => n8627, B2 => 
                           n8516, ZN => n1599);
   U733 : OAI22_X1 port map( A1 => n10346, A2 => n8517, B1 => n8628, B2 => 
                           n8516, ZN => n1598);
   U734 : OAI22_X1 port map( A1 => n10347, A2 => n8517, B1 => n8629, B2 => 
                           n8516, ZN => n1597);
   U735 : OAI22_X1 port map( A1 => n10348, A2 => n8517, B1 => n8630, B2 => 
                           n8516, ZN => n1596);
   U736 : OAI22_X1 port map( A1 => n10617, A2 => n8517, B1 => n8631, B2 => 
                           n8516, ZN => n1595);
   U737 : OAI22_X1 port map( A1 => n10618, A2 => n8517, B1 => n8632, B2 => 
                           n8516, ZN => n1594);
   U738 : OAI22_X1 port map( A1 => n10619, A2 => n8517, B1 => n8633, B2 => 
                           n8516, ZN => n1593);
   U739 : OAI22_X1 port map( A1 => n10349, A2 => n8517, B1 => n8634, B2 => 
                           n8516, ZN => n1592);
   U740 : OAI22_X1 port map( A1 => n10620, A2 => n8517, B1 => n8636, B2 => 
                           n8516, ZN => n1591);
   U741 : NAND2_X1 port map( A1 => n8581, A2 => n8565, ZN => n8539);
   U742 : CLKBUF_X1 port map( A => n8539, Z => n8549);
   U743 : OAI22_X1 port map( A1 => n10446, A2 => n8551, B1 => n8566, B2 => 
                           n8549, ZN => n1590);
   U744 : OAI22_X1 port map( A1 => n10350, A2 => n8551, B1 => n8518, B2 => 
                           n8539, ZN => n1589);
   U745 : OAI22_X1 port map( A1 => n10621, A2 => n8551, B1 => n8519, B2 => 
                           n8549, ZN => n1588);
   U746 : OAI22_X1 port map( A1 => n10351, A2 => n8551, B1 => n8520, B2 => 
                           n8539, ZN => n1587);
   U747 : OAI22_X1 port map( A1 => n10352, A2 => n8551, B1 => n8521, B2 => 
                           n8549, ZN => n1586);
   U748 : OAI22_X1 port map( A1 => n10353, A2 => n8551, B1 => n8522, B2 => 
                           n8539, ZN => n1585);
   U749 : OAI22_X1 port map( A1 => n10354, A2 => n8551, B1 => n8523, B2 => 
                           n8549, ZN => n1584);
   U750 : OAI22_X1 port map( A1 => n10355, A2 => n8551, B1 => n8524, B2 => 
                           n8539, ZN => n1583);
   U751 : OAI22_X1 port map( A1 => n10356, A2 => n8551, B1 => n8525, B2 => 
                           n8549, ZN => n1582);
   U752 : OAI22_X1 port map( A1 => n10357, A2 => n8551, B1 => n8526, B2 => 
                           n8539, ZN => n1581);
   U753 : OAI22_X1 port map( A1 => n10358, A2 => n8551, B1 => n8527, B2 => 
                           n8539, ZN => n1580);
   U754 : OAI22_X1 port map( A1 => n10622, A2 => n8551, B1 => n8528, B2 => 
                           n8549, ZN => n1579);
   U755 : OAI22_X1 port map( A1 => n10359, A2 => n8551, B1 => n8529, B2 => 
                           n8539, ZN => n1578);
   U756 : OAI22_X1 port map( A1 => n10360, A2 => n8551, B1 => n8530, B2 => 
                           n8549, ZN => n1577);
   U757 : OAI22_X1 port map( A1 => n10623, A2 => n8551, B1 => n8531, B2 => 
                           n8539, ZN => n1576);
   U758 : OAI22_X1 port map( A1 => n10361, A2 => n8551, B1 => n8532, B2 => 
                           n8549, ZN => n1575);
   U759 : OAI22_X1 port map( A1 => n10362, A2 => n8551, B1 => n8533, B2 => 
                           n8539, ZN => n1574);
   U760 : OAI22_X1 port map( A1 => n10363, A2 => n8551, B1 => n8534, B2 => 
                           n8539, ZN => n1573);
   U761 : OAI22_X1 port map( A1 => n10624, A2 => n8551, B1 => n8535, B2 => 
                           n8539, ZN => n1572);
   U762 : OAI22_X1 port map( A1 => n10364, A2 => n8551, B1 => n8536, B2 => 
                           n8539, ZN => n1571);
   U763 : OAI22_X1 port map( A1 => n10365, A2 => n8551, B1 => n8537, B2 => 
                           n8539, ZN => n1570);
   U764 : OAI22_X1 port map( A1 => n10366, A2 => n8551, B1 => n8538, B2 => 
                           n8539, ZN => n1569);
   U765 : OAI22_X1 port map( A1 => n10367, A2 => n8551, B1 => n8540, B2 => 
                           n8539, ZN => n1568);
   U766 : OAI22_X1 port map( A1 => n10856, A2 => n8551, B1 => n8541, B2 => 
                           n8549, ZN => n1567);
   U767 : OAI22_X1 port map( A1 => n10625, A2 => n8551, B1 => n8542, B2 => 
                           n8549, ZN => n1566);
   U768 : OAI22_X1 port map( A1 => n10626, A2 => n8551, B1 => n8543, B2 => 
                           n8549, ZN => n1565);
   U769 : OAI22_X1 port map( A1 => n10627, A2 => n8551, B1 => n8544, B2 => 
                           n8549, ZN => n1564);
   U770 : OAI22_X1 port map( A1 => n10368, A2 => n8551, B1 => n8545, B2 => 
                           n8549, ZN => n1563);
   U771 : OAI22_X1 port map( A1 => n10628, A2 => n8551, B1 => n8546, B2 => 
                           n8549, ZN => n1562);
   U772 : OAI22_X1 port map( A1 => n10369, A2 => n8551, B1 => n8547, B2 => 
                           n8549, ZN => n1561);
   U773 : OAI22_X1 port map( A1 => n10629, A2 => n8551, B1 => n8548, B2 => 
                           n8549, ZN => n1560);
   U774 : OAI22_X1 port map( A1 => n11115, A2 => n8551, B1 => n8550, B2 => 
                           n8549, ZN => n1559);
   U775 : NAND2_X1 port map( A1 => n8585, A2 => n8565, ZN => n8552);
   U776 : CLKBUF_X1 port map( A => n8552, Z => n8553);
   U777 : OAI22_X1 port map( A1 => n10718, A2 => n8554, B1 => n8566, B2 => 
                           n8553, ZN => n1558);
   U778 : OAI22_X1 port map( A1 => n11116, A2 => n8554, B1 => n8604, B2 => 
                           n8552, ZN => n1557);
   U779 : OAI22_X1 port map( A1 => n10857, A2 => n8554, B1 => n8605, B2 => 
                           n8553, ZN => n1556);
   U780 : OAI22_X1 port map( A1 => n10630, A2 => n8554, B1 => n8606, B2 => 
                           n8552, ZN => n1555);
   U781 : OAI22_X1 port map( A1 => n10858, A2 => n8554, B1 => n8607, B2 => 
                           n8553, ZN => n1554);
   U782 : OAI22_X1 port map( A1 => n11117, A2 => n8554, B1 => n8608, B2 => 
                           n8552, ZN => n1553);
   U783 : OAI22_X1 port map( A1 => n10859, A2 => n8554, B1 => n8609, B2 => 
                           n8553, ZN => n1552);
   U784 : OAI22_X1 port map( A1 => n10860, A2 => n8554, B1 => n8610, B2 => 
                           n8552, ZN => n1551);
   U785 : OAI22_X1 port map( A1 => n11118, A2 => n8554, B1 => n8611, B2 => 
                           n8553, ZN => n1550);
   U786 : OAI22_X1 port map( A1 => n11119, A2 => n8554, B1 => n8612, B2 => 
                           n8552, ZN => n1549);
   U787 : OAI22_X1 port map( A1 => n11120, A2 => n8554, B1 => n8613, B2 => 
                           n8552, ZN => n1548);
   U788 : OAI22_X1 port map( A1 => n10861, A2 => n8554, B1 => n8614, B2 => 
                           n8553, ZN => n1547);
   U789 : OAI22_X1 port map( A1 => n10631, A2 => n8554, B1 => n8615, B2 => 
                           n8552, ZN => n1546);
   U790 : OAI22_X1 port map( A1 => n10862, A2 => n8554, B1 => n8616, B2 => 
                           n8553, ZN => n1545);
   U791 : OAI22_X1 port map( A1 => n10863, A2 => n8554, B1 => n8617, B2 => 
                           n8552, ZN => n1544);
   U792 : OAI22_X1 port map( A1 => n11121, A2 => n8554, B1 => n8618, B2 => 
                           n8553, ZN => n1543);
   U793 : OAI22_X1 port map( A1 => n10370, A2 => n8554, B1 => n8619, B2 => 
                           n8552, ZN => n1542);
   U794 : OAI22_X1 port map( A1 => n10864, A2 => n8554, B1 => n8620, B2 => 
                           n8552, ZN => n1541);
   U795 : OAI22_X1 port map( A1 => n10865, A2 => n8554, B1 => n8621, B2 => 
                           n8552, ZN => n1540);
   U796 : OAI22_X1 port map( A1 => n10371, A2 => n8554, B1 => n8622, B2 => 
                           n8552, ZN => n1539);
   U797 : OAI22_X1 port map( A1 => n11122, A2 => n8554, B1 => n8623, B2 => 
                           n8552, ZN => n1538);
   U798 : OAI22_X1 port map( A1 => n11123, A2 => n8554, B1 => n8624, B2 => 
                           n8552, ZN => n1537);
   U799 : OAI22_X1 port map( A1 => n11124, A2 => n8554, B1 => n8626, B2 => 
                           n8552, ZN => n1536);
   U800 : OAI22_X1 port map( A1 => n11125, A2 => n8554, B1 => n8627, B2 => 
                           n8553, ZN => n1535);
   U801 : OAI22_X1 port map( A1 => n10372, A2 => n8554, B1 => n8628, B2 => 
                           n8553, ZN => n1534);
   U802 : OAI22_X1 port map( A1 => n11126, A2 => n8554, B1 => n8629, B2 => 
                           n8553, ZN => n1533);
   U803 : OAI22_X1 port map( A1 => n10632, A2 => n8554, B1 => n8630, B2 => 
                           n8553, ZN => n1532);
   U804 : OAI22_X1 port map( A1 => n10866, A2 => n8554, B1 => n8631, B2 => 
                           n8553, ZN => n1531);
   U805 : OAI22_X1 port map( A1 => n10633, A2 => n8554, B1 => n8632, B2 => 
                           n8553, ZN => n1530);
   U806 : OAI22_X1 port map( A1 => n10867, A2 => n8554, B1 => n8633, B2 => 
                           n8553, ZN => n1529);
   U807 : OAI22_X1 port map( A1 => n10373, A2 => n8554, B1 => n8634, B2 => 
                           n8553, ZN => n1528);
   U808 : OAI22_X1 port map( A1 => n10868, A2 => n8554, B1 => n8636, B2 => 
                           n8553, ZN => n1527);
   U809 : NAND2_X1 port map( A1 => n8589, A2 => n8565, ZN => n8555);
   U810 : CLKBUF_X1 port map( A => n8555, Z => n8556);
   U811 : OAI22_X1 port map( A1 => n10447, A2 => n8557, B1 => n8566, B2 => 
                           n8556, ZN => n1526);
   U812 : OAI22_X1 port map( A1 => n11127, A2 => n8557, B1 => n8604, B2 => 
                           n8555, ZN => n1525);
   U813 : OAI22_X1 port map( A1 => n11128, A2 => n8557, B1 => n8605, B2 => 
                           n8556, ZN => n1524);
   U814 : OAI22_X1 port map( A1 => n10869, A2 => n8557, B1 => n8606, B2 => 
                           n8555, ZN => n1523);
   U815 : OAI22_X1 port map( A1 => n11129, A2 => n8557, B1 => n8607, B2 => 
                           n8556, ZN => n1522);
   U816 : OAI22_X1 port map( A1 => n11130, A2 => n8557, B1 => n8608, B2 => 
                           n8555, ZN => n1521);
   U817 : OAI22_X1 port map( A1 => n10634, A2 => n8557, B1 => n8609, B2 => 
                           n8556, ZN => n1520);
   U818 : OAI22_X1 port map( A1 => n10635, A2 => n8557, B1 => n8610, B2 => 
                           n8555, ZN => n1519);
   U819 : OAI22_X1 port map( A1 => n10870, A2 => n8557, B1 => n8611, B2 => 
                           n8556, ZN => n1518);
   U820 : OAI22_X1 port map( A1 => n10374, A2 => n8557, B1 => n8612, B2 => 
                           n8555, ZN => n1517);
   U821 : OAI22_X1 port map( A1 => n10636, A2 => n8557, B1 => n8613, B2 => 
                           n8555, ZN => n1516);
   U822 : OAI22_X1 port map( A1 => n10871, A2 => n8557, B1 => n8614, B2 => 
                           n8556, ZN => n1515);
   U823 : OAI22_X1 port map( A1 => n10872, A2 => n8557, B1 => n8615, B2 => 
                           n8555, ZN => n1514);
   U824 : OAI22_X1 port map( A1 => n11131, A2 => n8557, B1 => n8616, B2 => 
                           n8556, ZN => n1513);
   U825 : OAI22_X1 port map( A1 => n10637, A2 => n8557, B1 => n8617, B2 => 
                           n8555, ZN => n1512);
   U826 : OAI22_X1 port map( A1 => n11132, A2 => n8557, B1 => n8618, B2 => 
                           n8556, ZN => n1511);
   U827 : OAI22_X1 port map( A1 => n10638, A2 => n8557, B1 => n8619, B2 => 
                           n8555, ZN => n1510);
   U828 : OAI22_X1 port map( A1 => n10873, A2 => n8557, B1 => n8620, B2 => 
                           n8555, ZN => n1509);
   U829 : OAI22_X1 port map( A1 => n10874, A2 => n8557, B1 => n8621, B2 => 
                           n8555, ZN => n1508);
   U830 : OAI22_X1 port map( A1 => n11133, A2 => n8557, B1 => n8622, B2 => 
                           n8555, ZN => n1507);
   U831 : OAI22_X1 port map( A1 => n10875, A2 => n8557, B1 => n8623, B2 => 
                           n8555, ZN => n1506);
   U832 : OAI22_X1 port map( A1 => n10876, A2 => n8557, B1 => n8624, B2 => 
                           n8555, ZN => n1505);
   U833 : OAI22_X1 port map( A1 => n11134, A2 => n8557, B1 => n8626, B2 => 
                           n8555, ZN => n1504);
   U834 : OAI22_X1 port map( A1 => n11135, A2 => n8557, B1 => n8627, B2 => 
                           n8556, ZN => n1503);
   U835 : OAI22_X1 port map( A1 => n10877, A2 => n8557, B1 => n8628, B2 => 
                           n8556, ZN => n1502);
   U836 : OAI22_X1 port map( A1 => n10375, A2 => n8557, B1 => n8629, B2 => 
                           n8556, ZN => n1501);
   U837 : OAI22_X1 port map( A1 => n10878, A2 => n8557, B1 => n8630, B2 => 
                           n8556, ZN => n1500);
   U838 : OAI22_X1 port map( A1 => n10879, A2 => n8557, B1 => n8631, B2 => 
                           n8556, ZN => n1499);
   U839 : OAI22_X1 port map( A1 => n11136, A2 => n8557, B1 => n8632, B2 => 
                           n8556, ZN => n1498);
   U840 : OAI22_X1 port map( A1 => n10376, A2 => n8557, B1 => n8633, B2 => 
                           n8556, ZN => n1497);
   U841 : OAI22_X1 port map( A1 => n10880, A2 => n8557, B1 => n8634, B2 => 
                           n8556, ZN => n1496);
   U842 : OAI22_X1 port map( A1 => n10639, A2 => n8557, B1 => n8636, B2 => 
                           n8556, ZN => n1495);
   U843 : NAND2_X1 port map( A1 => n8593, A2 => n8565, ZN => n8558);
   U844 : CLKBUF_X1 port map( A => n8561, Z => n8559);
   U845 : CLKBUF_X1 port map( A => n8558, Z => n8560);
   U846 : OAI22_X1 port map( A1 => n10719, A2 => n8559, B1 => n8566, B2 => 
                           n8560, ZN => n1494);
   U847 : OAI22_X1 port map( A1 => n10881, A2 => n8561, B1 => n8604, B2 => 
                           n8558, ZN => n1493);
   U848 : OAI22_X1 port map( A1 => n10377, A2 => n8559, B1 => n8605, B2 => 
                           n8560, ZN => n1492);
   U849 : OAI22_X1 port map( A1 => n10882, A2 => n8561, B1 => n8606, B2 => 
                           n8558, ZN => n1491);
   U850 : OAI22_X1 port map( A1 => n10883, A2 => n8559, B1 => n8607, B2 => 
                           n8560, ZN => n1490);
   U851 : OAI22_X1 port map( A1 => n10884, A2 => n8561, B1 => n8608, B2 => 
                           n8558, ZN => n1489);
   U852 : OAI22_X1 port map( A1 => n11137, A2 => n8559, B1 => n8609, B2 => 
                           n8560, ZN => n1488);
   U853 : OAI22_X1 port map( A1 => n11138, A2 => n8561, B1 => n8610, B2 => 
                           n8558, ZN => n1487);
   U854 : OAI22_X1 port map( A1 => n11139, A2 => n8559, B1 => n8611, B2 => 
                           n8560, ZN => n1486);
   U855 : OAI22_X1 port map( A1 => n10885, A2 => n8561, B1 => n8612, B2 => 
                           n8558, ZN => n1485);
   U856 : OAI22_X1 port map( A1 => n10886, A2 => n8561, B1 => n8613, B2 => 
                           n8558, ZN => n1484);
   U857 : OAI22_X1 port map( A1 => n10887, A2 => n8561, B1 => n8614, B2 => 
                           n8560, ZN => n1483);
   U858 : OAI22_X1 port map( A1 => n10888, A2 => n8559, B1 => n8615, B2 => 
                           n8558, ZN => n1482);
   U859 : OAI22_X1 port map( A1 => n11140, A2 => n8559, B1 => n8616, B2 => 
                           n8560, ZN => n1481);
   U860 : OAI22_X1 port map( A1 => n11141, A2 => n8559, B1 => n8617, B2 => 
                           n8558, ZN => n1480);
   U861 : OAI22_X1 port map( A1 => n10378, A2 => n8559, B1 => n8618, B2 => 
                           n8560, ZN => n1479);
   U862 : OAI22_X1 port map( A1 => n11142, A2 => n8559, B1 => n8619, B2 => 
                           n8558, ZN => n1478);
   U863 : OAI22_X1 port map( A1 => n11143, A2 => n8559, B1 => n8620, B2 => 
                           n8558, ZN => n1477);
   U864 : OAI22_X1 port map( A1 => n11144, A2 => n8559, B1 => n8621, B2 => 
                           n8558, ZN => n1476);
   U865 : OAI22_X1 port map( A1 => n10640, A2 => n8559, B1 => n8622, B2 => 
                           n8558, ZN => n1475);
   U866 : OAI22_X1 port map( A1 => n10889, A2 => n8559, B1 => n8623, B2 => 
                           n8558, ZN => n1474);
   U867 : OAI22_X1 port map( A1 => n11145, A2 => n8559, B1 => n8624, B2 => 
                           n8558, ZN => n1473);
   U868 : OAI22_X1 port map( A1 => n11146, A2 => n8559, B1 => n8626, B2 => 
                           n8558, ZN => n1472);
   U869 : OAI22_X1 port map( A1 => n10890, A2 => n8559, B1 => n8627, B2 => 
                           n8560, ZN => n1471);
   U870 : OAI22_X1 port map( A1 => n11147, A2 => n8561, B1 => n8628, B2 => 
                           n8560, ZN => n1470);
   U871 : OAI22_X1 port map( A1 => n10891, A2 => n8561, B1 => n8629, B2 => 
                           n8560, ZN => n1469);
   U872 : OAI22_X1 port map( A1 => n10892, A2 => n8561, B1 => n8630, B2 => 
                           n8560, ZN => n1468);
   U873 : OAI22_X1 port map( A1 => n11148, A2 => n8561, B1 => n8631, B2 => 
                           n8560, ZN => n1467);
   U874 : OAI22_X1 port map( A1 => n10893, A2 => n8561, B1 => n8632, B2 => 
                           n8560, ZN => n1466);
   U875 : OAI22_X1 port map( A1 => n11149, A2 => n8561, B1 => n8633, B2 => 
                           n8560, ZN => n1465);
   U876 : OAI22_X1 port map( A1 => n11150, A2 => n8561, B1 => n8634, B2 => 
                           n8560, ZN => n1464);
   U877 : OAI22_X1 port map( A1 => n10379, A2 => n8561, B1 => n8636, B2 => 
                           n8560, ZN => n1463);
   U878 : NAND2_X1 port map( A1 => n8597, A2 => n8565, ZN => n8562);
   U879 : CLKBUF_X1 port map( A => n8562, Z => n8563);
   U880 : OAI22_X1 port map( A1 => n10448, A2 => n8564, B1 => n8566, B2 => 
                           n8563, ZN => n1462);
   U881 : OAI22_X1 port map( A1 => n11151, A2 => n8564, B1 => n8604, B2 => 
                           n8562, ZN => n1461);
   U882 : OAI22_X1 port map( A1 => n11152, A2 => n8564, B1 => n8605, B2 => 
                           n8563, ZN => n1460);
   U883 : OAI22_X1 port map( A1 => n10894, A2 => n8564, B1 => n8606, B2 => 
                           n8562, ZN => n1459);
   U884 : OAI22_X1 port map( A1 => n11153, A2 => n8564, B1 => n8607, B2 => 
                           n8563, ZN => n1458);
   U885 : OAI22_X1 port map( A1 => n10641, A2 => n8564, B1 => n8608, B2 => 
                           n8562, ZN => n1457);
   U886 : OAI22_X1 port map( A1 => n11154, A2 => n8564, B1 => n8609, B2 => 
                           n8563, ZN => n1456);
   U887 : OAI22_X1 port map( A1 => n11155, A2 => n8564, B1 => n8610, B2 => 
                           n8562, ZN => n1455);
   U888 : OAI22_X1 port map( A1 => n11156, A2 => n8564, B1 => n8611, B2 => 
                           n8563, ZN => n1454);
   U889 : OAI22_X1 port map( A1 => n10895, A2 => n8564, B1 => n8612, B2 => 
                           n8562, ZN => n1453);
   U890 : OAI22_X1 port map( A1 => n11157, A2 => n8564, B1 => n8613, B2 => 
                           n8562, ZN => n1452);
   U891 : OAI22_X1 port map( A1 => n10896, A2 => n8564, B1 => n8614, B2 => 
                           n8563, ZN => n1451);
   U892 : OAI22_X1 port map( A1 => n10897, A2 => n8564, B1 => n8615, B2 => 
                           n8562, ZN => n1450);
   U893 : OAI22_X1 port map( A1 => n11158, A2 => n8564, B1 => n8616, B2 => 
                           n8563, ZN => n1449);
   U894 : OAI22_X1 port map( A1 => n10898, A2 => n8564, B1 => n8617, B2 => 
                           n8562, ZN => n1448);
   U895 : OAI22_X1 port map( A1 => n11159, A2 => n8564, B1 => n8618, B2 => 
                           n8563, ZN => n1447);
   U896 : OAI22_X1 port map( A1 => n11160, A2 => n8564, B1 => n8619, B2 => 
                           n8562, ZN => n1446);
   U897 : OAI22_X1 port map( A1 => n11161, A2 => n8564, B1 => n8620, B2 => 
                           n8562, ZN => n1445);
   U898 : OAI22_X1 port map( A1 => n10899, A2 => n8564, B1 => n8621, B2 => 
                           n8562, ZN => n1444);
   U899 : OAI22_X1 port map( A1 => n10900, A2 => n8564, B1 => n8622, B2 => 
                           n8562, ZN => n1443);
   U900 : OAI22_X1 port map( A1 => n11162, A2 => n8564, B1 => n8623, B2 => 
                           n8562, ZN => n1442);
   U901 : OAI22_X1 port map( A1 => n10642, A2 => n8564, B1 => n8624, B2 => 
                           n8562, ZN => n1441);
   U902 : OAI22_X1 port map( A1 => n10901, A2 => n8564, B1 => n8626, B2 => 
                           n8562, ZN => n1440);
   U903 : OAI22_X1 port map( A1 => n10643, A2 => n8564, B1 => n8627, B2 => 
                           n8563, ZN => n1439);
   U904 : OAI22_X1 port map( A1 => n10902, A2 => n8564, B1 => n8628, B2 => 
                           n8563, ZN => n1438);
   U905 : OAI22_X1 port map( A1 => n10903, A2 => n8564, B1 => n8629, B2 => 
                           n8563, ZN => n1437);
   U906 : OAI22_X1 port map( A1 => n11163, A2 => n8564, B1 => n8630, B2 => 
                           n8563, ZN => n1436);
   U907 : OAI22_X1 port map( A1 => n10904, A2 => n8564, B1 => n8631, B2 => 
                           n8563, ZN => n1435);
   U908 : OAI22_X1 port map( A1 => n11164, A2 => n8564, B1 => n8632, B2 => 
                           n8563, ZN => n1434);
   U909 : OAI22_X1 port map( A1 => n10380, A2 => n8564, B1 => n8633, B2 => 
                           n8563, ZN => n1433);
   U910 : OAI22_X1 port map( A1 => n11165, A2 => n8564, B1 => n8634, B2 => 
                           n8563, ZN => n1432);
   U911 : OAI22_X1 port map( A1 => n10905, A2 => n8564, B1 => n8636, B2 => 
                           n8563, ZN => n1431);
   U912 : NAND2_X1 port map( A1 => n8602, A2 => n8565, ZN => n8567);
   U913 : CLKBUF_X1 port map( A => n8567, Z => n8568);
   U914 : OAI22_X1 port map( A1 => n10203, A2 => n8569, B1 => n8566, B2 => 
                           n8568, ZN => n1430);
   U915 : OAI22_X1 port map( A1 => n10906, A2 => n8569, B1 => n8604, B2 => 
                           n8567, ZN => n1429);
   U916 : OAI22_X1 port map( A1 => n11166, A2 => n8569, B1 => n8605, B2 => 
                           n8568, ZN => n1428);
   U917 : OAI22_X1 port map( A1 => n10381, A2 => n8569, B1 => n8606, B2 => 
                           n8567, ZN => n1427);
   U918 : OAI22_X1 port map( A1 => n11167, A2 => n8569, B1 => n8607, B2 => 
                           n8568, ZN => n1426);
   U919 : OAI22_X1 port map( A1 => n11168, A2 => n8569, B1 => n8608, B2 => 
                           n8567, ZN => n1425);
   U920 : OAI22_X1 port map( A1 => n10382, A2 => n8569, B1 => n8609, B2 => 
                           n8568, ZN => n1424);
   U921 : OAI22_X1 port map( A1 => n11169, A2 => n8569, B1 => n8610, B2 => 
                           n8567, ZN => n1423);
   U922 : OAI22_X1 port map( A1 => n10383, A2 => n8569, B1 => n8611, B2 => 
                           n8568, ZN => n1422);
   U923 : OAI22_X1 port map( A1 => n10644, A2 => n8569, B1 => n8612, B2 => 
                           n8567, ZN => n1421);
   U924 : OAI22_X1 port map( A1 => n10907, A2 => n8569, B1 => n8613, B2 => 
                           n8567, ZN => n1420);
   U925 : OAI22_X1 port map( A1 => n10645, A2 => n8569, B1 => n8614, B2 => 
                           n8568, ZN => n1419);
   U926 : OAI22_X1 port map( A1 => n10384, A2 => n8569, B1 => n8615, B2 => 
                           n8567, ZN => n1418);
   U927 : OAI22_X1 port map( A1 => n10646, A2 => n8569, B1 => n8616, B2 => 
                           n8568, ZN => n1417);
   U928 : OAI22_X1 port map( A1 => n10385, A2 => n8569, B1 => n8617, B2 => 
                           n8567, ZN => n1416);
   U929 : OAI22_X1 port map( A1 => n11170, A2 => n8569, B1 => n8618, B2 => 
                           n8568, ZN => n1415);
   U930 : OAI22_X1 port map( A1 => n10908, A2 => n8569, B1 => n8619, B2 => 
                           n8567, ZN => n1414);
   U931 : OAI22_X1 port map( A1 => n11171, A2 => n8569, B1 => n8620, B2 => 
                           n8567, ZN => n1413);
   U932 : OAI22_X1 port map( A1 => n10909, A2 => n8569, B1 => n8621, B2 => 
                           n8567, ZN => n1412);
   U933 : OAI22_X1 port map( A1 => n10647, A2 => n8569, B1 => n8622, B2 => 
                           n8567, ZN => n1411);
   U934 : OAI22_X1 port map( A1 => n10648, A2 => n8569, B1 => n8623, B2 => 
                           n8567, ZN => n1410);
   U935 : OAI22_X1 port map( A1 => n11172, A2 => n8569, B1 => n8624, B2 => 
                           n8567, ZN => n1409);
   U936 : OAI22_X1 port map( A1 => n10910, A2 => n8569, B1 => n8626, B2 => 
                           n8567, ZN => n1408);
   U937 : OAI22_X1 port map( A1 => n10649, A2 => n8569, B1 => n8627, B2 => 
                           n8568, ZN => n1407);
   U938 : OAI22_X1 port map( A1 => n10386, A2 => n8569, B1 => n8628, B2 => 
                           n8568, ZN => n1406);
   U939 : OAI22_X1 port map( A1 => n10650, A2 => n8569, B1 => n8629, B2 => 
                           n8568, ZN => n1405);
   U940 : OAI22_X1 port map( A1 => n10651, A2 => n8569, B1 => n8630, B2 => 
                           n8568, ZN => n1404);
   U941 : OAI22_X1 port map( A1 => n10911, A2 => n8569, B1 => n8631, B2 => 
                           n8568, ZN => n1403);
   U942 : OAI22_X1 port map( A1 => n10387, A2 => n8569, B1 => n8632, B2 => 
                           n8568, ZN => n1402);
   U943 : OAI22_X1 port map( A1 => n11173, A2 => n8569, B1 => n8633, B2 => 
                           n8568, ZN => n1401);
   U944 : OAI22_X1 port map( A1 => n10912, A2 => n8569, B1 => n8634, B2 => 
                           n8568, ZN => n1400);
   U945 : OAI22_X1 port map( A1 => n10388, A2 => n8569, B1 => n8636, B2 => 
                           n8568, ZN => n1399);
   U946 : NOR2_X1 port map( A1 => n8571, A2 => n8570, ZN => n8601);
   U947 : NAND2_X1 port map( A1 => n8572, A2 => n8601, ZN => n8573);
   U948 : CLKBUF_X1 port map( A => n8573, Z => n8574);
   U949 : OAI22_X1 port map( A1 => n10449, A2 => n8575, B1 => n8603, B2 => 
                           n8574, ZN => n1398);
   U950 : OAI22_X1 port map( A1 => n10389, A2 => n8575, B1 => n8604, B2 => 
                           n8573, ZN => n1397);
   U951 : OAI22_X1 port map( A1 => n10390, A2 => n8575, B1 => n8605, B2 => 
                           n8574, ZN => n1396);
   U952 : OAI22_X1 port map( A1 => n11174, A2 => n8575, B1 => n8606, B2 => 
                           n8573, ZN => n1395);
   U953 : OAI22_X1 port map( A1 => n10652, A2 => n8575, B1 => n8607, B2 => 
                           n8574, ZN => n1394);
   U954 : OAI22_X1 port map( A1 => n10913, A2 => n8575, B1 => n8608, B2 => 
                           n8573, ZN => n1393);
   U955 : OAI22_X1 port map( A1 => n11175, A2 => n8575, B1 => n8609, B2 => 
                           n8574, ZN => n1392);
   U956 : OAI22_X1 port map( A1 => n10653, A2 => n8575, B1 => n8610, B2 => 
                           n8573, ZN => n1391);
   U957 : OAI22_X1 port map( A1 => n10654, A2 => n8575, B1 => n8611, B2 => 
                           n8574, ZN => n1390);
   U958 : OAI22_X1 port map( A1 => n11176, A2 => n8575, B1 => n8612, B2 => 
                           n8573, ZN => n1389);
   U959 : OAI22_X1 port map( A1 => n10655, A2 => n8575, B1 => n8613, B2 => 
                           n8573, ZN => n1388);
   U960 : OAI22_X1 port map( A1 => n10391, A2 => n8575, B1 => n8614, B2 => 
                           n8574, ZN => n1387);
   U961 : OAI22_X1 port map( A1 => n11177, A2 => n8575, B1 => n8615, B2 => 
                           n8573, ZN => n1386);
   U962 : OAI22_X1 port map( A1 => n10914, A2 => n8575, B1 => n8616, B2 => 
                           n8574, ZN => n1385);
   U963 : OAI22_X1 port map( A1 => n11178, A2 => n8575, B1 => n8617, B2 => 
                           n8573, ZN => n1384);
   U964 : OAI22_X1 port map( A1 => n10656, A2 => n8575, B1 => n8618, B2 => 
                           n8574, ZN => n1383);
   U965 : OAI22_X1 port map( A1 => n10915, A2 => n8575, B1 => n8619, B2 => 
                           n8573, ZN => n1382);
   U966 : OAI22_X1 port map( A1 => n10392, A2 => n8575, B1 => n8620, B2 => 
                           n8573, ZN => n1381);
   U967 : OAI22_X1 port map( A1 => n10657, A2 => n8575, B1 => n8621, B2 => 
                           n8573, ZN => n1380);
   U968 : OAI22_X1 port map( A1 => n10916, A2 => n8575, B1 => n8622, B2 => 
                           n8573, ZN => n1379);
   U969 : OAI22_X1 port map( A1 => n11179, A2 => n8575, B1 => n8623, B2 => 
                           n8573, ZN => n1378);
   U970 : OAI22_X1 port map( A1 => n10658, A2 => n8575, B1 => n8624, B2 => 
                           n8573, ZN => n1377);
   U971 : OAI22_X1 port map( A1 => n10393, A2 => n8575, B1 => n8626, B2 => 
                           n8573, ZN => n1376);
   U972 : OAI22_X1 port map( A1 => n10394, A2 => n8575, B1 => n8627, B2 => 
                           n8574, ZN => n1375);
   U973 : OAI22_X1 port map( A1 => n10659, A2 => n8575, B1 => n8628, B2 => 
                           n8574, ZN => n1374);
   U974 : OAI22_X1 port map( A1 => n10395, A2 => n8575, B1 => n8629, B2 => 
                           n8574, ZN => n1373);
   U975 : OAI22_X1 port map( A1 => n10396, A2 => n8575, B1 => n8630, B2 => 
                           n8574, ZN => n1372);
   U976 : OAI22_X1 port map( A1 => n11180, A2 => n8575, B1 => n8631, B2 => 
                           n8574, ZN => n1371);
   U977 : OAI22_X1 port map( A1 => n11181, A2 => n8575, B1 => n8632, B2 => 
                           n8574, ZN => n1370);
   U978 : OAI22_X1 port map( A1 => n10397, A2 => n8575, B1 => n8633, B2 => 
                           n8574, ZN => n1369);
   U979 : OAI22_X1 port map( A1 => n10660, A2 => n8575, B1 => n8634, B2 => 
                           n8574, ZN => n1368);
   U980 : OAI22_X1 port map( A1 => n10398, A2 => n8575, B1 => n8636, B2 => 
                           n8574, ZN => n1367);
   U981 : NAND2_X1 port map( A1 => n8576, A2 => n8601, ZN => n8577);
   U982 : CLKBUF_X1 port map( A => n8580, Z => n8578);
   U983 : CLKBUF_X1 port map( A => n8577, Z => n8579);
   U984 : OAI22_X1 port map( A1 => n10450, A2 => n8578, B1 => n8603, B2 => 
                           n8579, ZN => n1366);
   U985 : OAI22_X1 port map( A1 => n10917, A2 => n8580, B1 => n8604, B2 => 
                           n8577, ZN => n1365);
   U986 : OAI22_X1 port map( A1 => n10918, A2 => n8578, B1 => n8605, B2 => 
                           n8579, ZN => n1364);
   U987 : OAI22_X1 port map( A1 => n10919, A2 => n8580, B1 => n8606, B2 => 
                           n8577, ZN => n1363);
   U988 : OAI22_X1 port map( A1 => n10399, A2 => n8578, B1 => n8607, B2 => 
                           n8579, ZN => n1362);
   U989 : OAI22_X1 port map( A1 => n10920, A2 => n8580, B1 => n8608, B2 => 
                           n8577, ZN => n1361);
   U990 : OAI22_X1 port map( A1 => n10661, A2 => n8578, B1 => n8609, B2 => 
                           n8579, ZN => n1360);
   U991 : OAI22_X1 port map( A1 => n10400, A2 => n8580, B1 => n8610, B2 => 
                           n8577, ZN => n1359);
   U992 : OAI22_X1 port map( A1 => n10401, A2 => n8578, B1 => n8611, B2 => 
                           n8579, ZN => n1358);
   U993 : OAI22_X1 port map( A1 => n10921, A2 => n8580, B1 => n8612, B2 => 
                           n8577, ZN => n1357);
   U994 : OAI22_X1 port map( A1 => n10922, A2 => n8580, B1 => n8613, B2 => 
                           n8577, ZN => n1356);
   U995 : OAI22_X1 port map( A1 => n10662, A2 => n8580, B1 => n8614, B2 => 
                           n8579, ZN => n1355);
   U996 : OAI22_X1 port map( A1 => n11182, A2 => n8578, B1 => n8615, B2 => 
                           n8577, ZN => n1354);
   U997 : OAI22_X1 port map( A1 => n10663, A2 => n8578, B1 => n8616, B2 => 
                           n8579, ZN => n1353);
   U998 : OAI22_X1 port map( A1 => n10402, A2 => n8578, B1 => n8617, B2 => 
                           n8577, ZN => n1352);
   U999 : OAI22_X1 port map( A1 => n10403, A2 => n8578, B1 => n8618, B2 => 
                           n8579, ZN => n1351);
   U1000 : OAI22_X1 port map( A1 => n11183, A2 => n8578, B1 => n8619, B2 => 
                           n8577, ZN => n1350);
   U1001 : OAI22_X1 port map( A1 => n10923, A2 => n8578, B1 => n8620, B2 => 
                           n8577, ZN => n1349);
   U1002 : OAI22_X1 port map( A1 => n10664, A2 => n8578, B1 => n8621, B2 => 
                           n8577, ZN => n1348);
   U1003 : OAI22_X1 port map( A1 => n10665, A2 => n8578, B1 => n8622, B2 => 
                           n8577, ZN => n1347);
   U1004 : OAI22_X1 port map( A1 => n10924, A2 => n8578, B1 => n8623, B2 => 
                           n8577, ZN => n1346);
   U1005 : OAI22_X1 port map( A1 => n10925, A2 => n8578, B1 => n8624, B2 => 
                           n8577, ZN => n1345);
   U1006 : OAI22_X1 port map( A1 => n10404, A2 => n8578, B1 => n8626, B2 => 
                           n8577, ZN => n1344);
   U1007 : OAI22_X1 port map( A1 => n11184, A2 => n8578, B1 => n8627, B2 => 
                           n8579, ZN => n1343);
   U1008 : OAI22_X1 port map( A1 => n11185, A2 => n8580, B1 => n8628, B2 => 
                           n8579, ZN => n1342);
   U1009 : OAI22_X1 port map( A1 => n11186, A2 => n8580, B1 => n8629, B2 => 
                           n8579, ZN => n1341);
   U1010 : OAI22_X1 port map( A1 => n10405, A2 => n8580, B1 => n8630, B2 => 
                           n8579, ZN => n1340);
   U1011 : OAI22_X1 port map( A1 => n10666, A2 => n8580, B1 => n8631, B2 => 
                           n8579, ZN => n1339);
   U1012 : OAI22_X1 port map( A1 => n10406, A2 => n8580, B1 => n8632, B2 => 
                           n8579, ZN => n1338);
   U1013 : OAI22_X1 port map( A1 => n10926, A2 => n8580, B1 => n8633, B2 => 
                           n8579, ZN => n1337);
   U1014 : OAI22_X1 port map( A1 => n11187, A2 => n8580, B1 => n8634, B2 => 
                           n8579, ZN => n1336);
   U1015 : OAI22_X1 port map( A1 => n10927, A2 => n8580, B1 => n8636, B2 => 
                           n8579, ZN => n1335);
   U1016 : NAND2_X1 port map( A1 => n8581, A2 => n8601, ZN => n8582);
   U1017 : CLKBUF_X1 port map( A => n8582, Z => n8583);
   U1018 : OAI22_X1 port map( A1 => n10720, A2 => n8584, B1 => n8603, B2 => 
                           n8583, ZN => n1334);
   U1019 : OAI22_X1 port map( A1 => n10667, A2 => n8584, B1 => n8604, B2 => 
                           n8582, ZN => n1333);
   U1020 : OAI22_X1 port map( A1 => n10668, A2 => n8584, B1 => n8605, B2 => 
                           n8583, ZN => n1332);
   U1021 : OAI22_X1 port map( A1 => n11188, A2 => n8584, B1 => n8606, B2 => 
                           n8582, ZN => n1331);
   U1022 : OAI22_X1 port map( A1 => n10407, A2 => n8584, B1 => n8607, B2 => 
                           n8583, ZN => n1330);
   U1023 : OAI22_X1 port map( A1 => n10669, A2 => n8584, B1 => n8608, B2 => 
                           n8582, ZN => n1329);
   U1024 : OAI22_X1 port map( A1 => n10408, A2 => n8584, B1 => n8609, B2 => 
                           n8583, ZN => n1328);
   U1025 : OAI22_X1 port map( A1 => n10670, A2 => n8584, B1 => n8610, B2 => 
                           n8582, ZN => n1327);
   U1026 : OAI22_X1 port map( A1 => n10671, A2 => n8584, B1 => n8611, B2 => 
                           n8583, ZN => n1326);
   U1027 : OAI22_X1 port map( A1 => n10409, A2 => n8584, B1 => n8612, B2 => 
                           n8582, ZN => n1325);
   U1028 : OAI22_X1 port map( A1 => n10672, A2 => n8584, B1 => n8613, B2 => 
                           n8582, ZN => n1324);
   U1029 : OAI22_X1 port map( A1 => n10410, A2 => n8584, B1 => n8614, B2 => 
                           n8583, ZN => n1323);
   U1030 : OAI22_X1 port map( A1 => n10673, A2 => n8584, B1 => n8615, B2 => 
                           n8582, ZN => n1322);
   U1031 : OAI22_X1 port map( A1 => n10674, A2 => n8584, B1 => n8616, B2 => 
                           n8583, ZN => n1321);
   U1032 : OAI22_X1 port map( A1 => n10411, A2 => n8584, B1 => n8617, B2 => 
                           n8582, ZN => n1320);
   U1033 : OAI22_X1 port map( A1 => n10675, A2 => n8584, B1 => n8618, B2 => 
                           n8583, ZN => n1319);
   U1034 : OAI22_X1 port map( A1 => n10412, A2 => n8584, B1 => n8619, B2 => 
                           n8582, ZN => n1318);
   U1035 : OAI22_X1 port map( A1 => n10676, A2 => n8584, B1 => n8620, B2 => 
                           n8582, ZN => n1317);
   U1036 : OAI22_X1 port map( A1 => n10677, A2 => n8584, B1 => n8621, B2 => 
                           n8582, ZN => n1316);
   U1037 : OAI22_X1 port map( A1 => n11189, A2 => n8584, B1 => n8622, B2 => 
                           n8582, ZN => n1315);
   U1038 : OAI22_X1 port map( A1 => n10413, A2 => n8584, B1 => n8623, B2 => 
                           n8582, ZN => n1314);
   U1039 : OAI22_X1 port map( A1 => n10928, A2 => n8584, B1 => n8624, B2 => 
                           n8582, ZN => n1313);
   U1040 : OAI22_X1 port map( A1 => n10414, A2 => n8584, B1 => n8626, B2 => 
                           n8582, ZN => n1312);
   U1041 : OAI22_X1 port map( A1 => n10415, A2 => n8584, B1 => n8627, B2 => 
                           n8583, ZN => n1311);
   U1042 : OAI22_X1 port map( A1 => n10678, A2 => n8584, B1 => n8628, B2 => 
                           n8583, ZN => n1310);
   U1043 : OAI22_X1 port map( A1 => n10416, A2 => n8584, B1 => n8629, B2 => 
                           n8583, ZN => n1309);
   U1044 : OAI22_X1 port map( A1 => n10679, A2 => n8584, B1 => n8630, B2 => 
                           n8583, ZN => n1308);
   U1045 : OAI22_X1 port map( A1 => n10680, A2 => n8584, B1 => n8631, B2 => 
                           n8583, ZN => n1307);
   U1046 : OAI22_X1 port map( A1 => n10929, A2 => n8584, B1 => n8632, B2 => 
                           n8583, ZN => n1306);
   U1047 : OAI22_X1 port map( A1 => n10417, A2 => n8584, B1 => n8633, B2 => 
                           n8583, ZN => n1305);
   U1048 : OAI22_X1 port map( A1 => n10418, A2 => n8584, B1 => n8634, B2 => 
                           n8583, ZN => n1304);
   U1049 : OAI22_X1 port map( A1 => n10681, A2 => n8584, B1 => n8636, B2 => 
                           n8583, ZN => n1303);
   U1050 : NAND2_X1 port map( A1 => n8585, A2 => n8601, ZN => n8586);
   U1051 : CLKBUF_X1 port map( A => n8586, Z => n8587);
   U1052 : OAI22_X1 port map( A1 => n10204, A2 => n8588, B1 => n8603, B2 => 
                           n8587, ZN => n1302);
   U1053 : OAI22_X1 port map( A1 => n10682, A2 => n8588, B1 => n8604, B2 => 
                           n8586, ZN => n1301);
   U1054 : OAI22_X1 port map( A1 => n10683, A2 => n8588, B1 => n8605, B2 => 
                           n8587, ZN => n1300);
   U1055 : OAI22_X1 port map( A1 => n10684, A2 => n8588, B1 => n8606, B2 => 
                           n8586, ZN => n1299);
   U1056 : OAI22_X1 port map( A1 => n10930, A2 => n8588, B1 => n8607, B2 => 
                           n8587, ZN => n1298);
   U1057 : OAI22_X1 port map( A1 => n10419, A2 => n8588, B1 => n8608, B2 => 
                           n8586, ZN => n1297);
   U1058 : OAI22_X1 port map( A1 => n10685, A2 => n8588, B1 => n8609, B2 => 
                           n8587, ZN => n1296);
   U1059 : OAI22_X1 port map( A1 => n10686, A2 => n8588, B1 => n8610, B2 => 
                           n8586, ZN => n1295);
   U1060 : OAI22_X1 port map( A1 => n10420, A2 => n8588, B1 => n8611, B2 => 
                           n8587, ZN => n1294);
   U1061 : OAI22_X1 port map( A1 => n10421, A2 => n8588, B1 => n8612, B2 => 
                           n8586, ZN => n1293);
   U1062 : OAI22_X1 port map( A1 => n10422, A2 => n8588, B1 => n8613, B2 => 
                           n8586, ZN => n1292);
   U1063 : OAI22_X1 port map( A1 => n10687, A2 => n8588, B1 => n8614, B2 => 
                           n8587, ZN => n1291);
   U1064 : OAI22_X1 port map( A1 => n10423, A2 => n8588, B1 => n8615, B2 => 
                           n8586, ZN => n1290);
   U1065 : OAI22_X1 port map( A1 => n10424, A2 => n8588, B1 => n8616, B2 => 
                           n8587, ZN => n1289);
   U1066 : OAI22_X1 port map( A1 => n10425, A2 => n8588, B1 => n8617, B2 => 
                           n8586, ZN => n1288);
   U1067 : OAI22_X1 port map( A1 => n10688, A2 => n8588, B1 => n8618, B2 => 
                           n8587, ZN => n1287);
   U1068 : OAI22_X1 port map( A1 => n10426, A2 => n8588, B1 => n8619, B2 => 
                           n8586, ZN => n1286);
   U1069 : OAI22_X1 port map( A1 => n10689, A2 => n8588, B1 => n8620, B2 => 
                           n8586, ZN => n1285);
   U1070 : OAI22_X1 port map( A1 => n10427, A2 => n8588, B1 => n8621, B2 => 
                           n8586, ZN => n1284);
   U1071 : OAI22_X1 port map( A1 => n10690, A2 => n8588, B1 => n8622, B2 => 
                           n8586, ZN => n1283);
   U1072 : OAI22_X1 port map( A1 => n10691, A2 => n8588, B1 => n8623, B2 => 
                           n8586, ZN => n1282);
   U1073 : OAI22_X1 port map( A1 => n10692, A2 => n8588, B1 => n8624, B2 => 
                           n8586, ZN => n1281);
   U1074 : OAI22_X1 port map( A1 => n10693, A2 => n8588, B1 => n8626, B2 => 
                           n8586, ZN => n1280);
   U1075 : OAI22_X1 port map( A1 => n10428, A2 => n8588, B1 => n8627, B2 => 
                           n8587, ZN => n1279);
   U1076 : OAI22_X1 port map( A1 => n10429, A2 => n8588, B1 => n8628, B2 => 
                           n8587, ZN => n1278);
   U1077 : OAI22_X1 port map( A1 => n10694, A2 => n8588, B1 => n8629, B2 => 
                           n8587, ZN => n1277);
   U1078 : OAI22_X1 port map( A1 => n10695, A2 => n8588, B1 => n8630, B2 => 
                           n8587, ZN => n1276);
   U1079 : OAI22_X1 port map( A1 => n10696, A2 => n8588, B1 => n8631, B2 => 
                           n8587, ZN => n1275);
   U1080 : OAI22_X1 port map( A1 => n10697, A2 => n8588, B1 => n8632, B2 => 
                           n8587, ZN => n1274);
   U1081 : OAI22_X1 port map( A1 => n10698, A2 => n8588, B1 => n8633, B2 => 
                           n8587, ZN => n1273);
   U1082 : OAI22_X1 port map( A1 => n10430, A2 => n8588, B1 => n8634, B2 => 
                           n8587, ZN => n1272);
   U1083 : OAI22_X1 port map( A1 => n10699, A2 => n8588, B1 => n8636, B2 => 
                           n8587, ZN => n1271);
   U1084 : NAND2_X1 port map( A1 => n8589, A2 => n8601, ZN => n8590);
   U1085 : CLKBUF_X1 port map( A => n8590, Z => n8591);
   U1086 : OAI22_X1 port map( A1 => n10451, A2 => n8592, B1 => n8603, B2 => 
                           n8591, ZN => n1270);
   U1087 : OAI22_X1 port map( A1 => n11190, A2 => n8592, B1 => n8604, B2 => 
                           n8590, ZN => n1269);
   U1088 : OAI22_X1 port map( A1 => n10931, A2 => n8592, B1 => n8605, B2 => 
                           n8591, ZN => n1268);
   U1089 : OAI22_X1 port map( A1 => n11191, A2 => n8592, B1 => n8606, B2 => 
                           n8590, ZN => n1267);
   U1090 : OAI22_X1 port map( A1 => n11192, A2 => n8592, B1 => n8607, B2 => 
                           n8591, ZN => n1266);
   U1091 : OAI22_X1 port map( A1 => n10932, A2 => n8592, B1 => n8608, B2 => 
                           n8590, ZN => n1265);
   U1092 : OAI22_X1 port map( A1 => n10933, A2 => n8592, B1 => n8609, B2 => 
                           n8591, ZN => n1264);
   U1093 : OAI22_X1 port map( A1 => n10934, A2 => n8592, B1 => n8610, B2 => 
                           n8590, ZN => n1263);
   U1094 : OAI22_X1 port map( A1 => n10935, A2 => n8592, B1 => n8611, B2 => 
                           n8591, ZN => n1262);
   U1095 : OAI22_X1 port map( A1 => n11193, A2 => n8592, B1 => n8612, B2 => 
                           n8590, ZN => n1261);
   U1096 : OAI22_X1 port map( A1 => n10936, A2 => n8592, B1 => n8613, B2 => 
                           n8590, ZN => n1260);
   U1097 : OAI22_X1 port map( A1 => n10937, A2 => n8592, B1 => n8614, B2 => 
                           n8591, ZN => n1259);
   U1098 : OAI22_X1 port map( A1 => n11194, A2 => n8592, B1 => n8615, B2 => 
                           n8590, ZN => n1258);
   U1099 : OAI22_X1 port map( A1 => n10938, A2 => n8592, B1 => n8616, B2 => 
                           n8591, ZN => n1257);
   U1100 : OAI22_X1 port map( A1 => n10700, A2 => n8592, B1 => n8617, B2 => 
                           n8590, ZN => n1256);
   U1101 : OAI22_X1 port map( A1 => n10939, A2 => n8592, B1 => n8618, B2 => 
                           n8591, ZN => n1255);
   U1102 : OAI22_X1 port map( A1 => n10940, A2 => n8592, B1 => n8619, B2 => 
                           n8590, ZN => n1254);
   U1103 : OAI22_X1 port map( A1 => n11195, A2 => n8592, B1 => n8620, B2 => 
                           n8590, ZN => n1253);
   U1104 : OAI22_X1 port map( A1 => n10941, A2 => n8592, B1 => n8621, B2 => 
                           n8590, ZN => n1252);
   U1105 : OAI22_X1 port map( A1 => n10942, A2 => n8592, B1 => n8622, B2 => 
                           n8590, ZN => n1251);
   U1106 : OAI22_X1 port map( A1 => n10943, A2 => n8592, B1 => n8623, B2 => 
                           n8590, ZN => n1250);
   U1107 : OAI22_X1 port map( A1 => n10944, A2 => n8592, B1 => n8624, B2 => 
                           n8590, ZN => n1249);
   U1108 : OAI22_X1 port map( A1 => n10945, A2 => n8592, B1 => n8626, B2 => 
                           n8590, ZN => n1248);
   U1109 : OAI22_X1 port map( A1 => n10946, A2 => n8592, B1 => n8627, B2 => 
                           n8591, ZN => n1247);
   U1110 : OAI22_X1 port map( A1 => n10947, A2 => n8592, B1 => n8628, B2 => 
                           n8591, ZN => n1246);
   U1111 : OAI22_X1 port map( A1 => n10948, A2 => n8592, B1 => n8629, B2 => 
                           n8591, ZN => n1245);
   U1112 : OAI22_X1 port map( A1 => n11196, A2 => n8592, B1 => n8630, B2 => 
                           n8591, ZN => n1244);
   U1113 : OAI22_X1 port map( A1 => n10949, A2 => n8592, B1 => n8631, B2 => 
                           n8591, ZN => n1243);
   U1114 : OAI22_X1 port map( A1 => n10950, A2 => n8592, B1 => n8632, B2 => 
                           n8591, ZN => n1242);
   U1115 : OAI22_X1 port map( A1 => n10951, A2 => n8592, B1 => n8633, B2 => 
                           n8591, ZN => n1241);
   U1116 : OAI22_X1 port map( A1 => n10952, A2 => n8592, B1 => n8634, B2 => 
                           n8591, ZN => n1240);
   U1117 : OAI22_X1 port map( A1 => n11197, A2 => n8592, B1 => n8636, B2 => 
                           n8591, ZN => n1239);
   U1118 : NAND2_X1 port map( A1 => n8593, A2 => n8601, ZN => n8594);
   U1119 : OAI22_X1 port map( A1 => n10452, A2 => n8596, B1 => n8603, B2 => 
                           n8595, ZN => n1238);
   U1120 : OAI22_X1 port map( A1 => n10701, A2 => n8596, B1 => n8604, B2 => 
                           n8594, ZN => n1237);
   U1121 : OAI22_X1 port map( A1 => n10431, A2 => n8596, B1 => n8605, B2 => 
                           n8595, ZN => n1236);
   U1122 : OAI22_X1 port map( A1 => n10702, A2 => n8596, B1 => n8606, B2 => 
                           n8594, ZN => n1235);
   U1123 : OAI22_X1 port map( A1 => n10432, A2 => n8596, B1 => n8607, B2 => 
                           n8595, ZN => n1234);
   U1124 : OAI22_X1 port map( A1 => n10433, A2 => n8596, B1 => n8608, B2 => 
                           n8594, ZN => n1233);
   U1125 : OAI22_X1 port map( A1 => n11198, A2 => n8596, B1 => n8609, B2 => 
                           n8595, ZN => n1232);
   U1126 : OAI22_X1 port map( A1 => n10953, A2 => n8596, B1 => n8610, B2 => 
                           n8594, ZN => n1231);
   U1127 : OAI22_X1 port map( A1 => n10954, A2 => n8596, B1 => n8611, B2 => 
                           n8595, ZN => n1230);
   U1128 : OAI22_X1 port map( A1 => n10955, A2 => n8596, B1 => n8612, B2 => 
                           n8594, ZN => n1229);
   U1129 : OAI22_X1 port map( A1 => n10956, A2 => n8596, B1 => n8613, B2 => 
                           n8594, ZN => n1228);
   U1130 : OAI22_X1 port map( A1 => n11199, A2 => n8596, B1 => n8614, B2 => 
                           n8595, ZN => n1227);
   U1131 : OAI22_X1 port map( A1 => n10957, A2 => n8596, B1 => n8615, B2 => 
                           n8594, ZN => n1226);
   U1132 : OAI22_X1 port map( A1 => n10958, A2 => n8596, B1 => n8616, B2 => 
                           n8595, ZN => n1225);
   U1133 : OAI22_X1 port map( A1 => n10959, A2 => n8596, B1 => n8617, B2 => 
                           n8594, ZN => n1224);
   U1134 : OAI22_X1 port map( A1 => n10960, A2 => n8596, B1 => n8618, B2 => 
                           n8595, ZN => n1223);
   U1135 : OAI22_X1 port map( A1 => n11200, A2 => n8596, B1 => n8619, B2 => 
                           n8594, ZN => n1222);
   U1136 : OAI22_X1 port map( A1 => n10703, A2 => n8596, B1 => n8620, B2 => 
                           n8594, ZN => n1221);
   U1137 : OAI22_X1 port map( A1 => n11201, A2 => n8596, B1 => n8621, B2 => 
                           n8594, ZN => n1220);
   U1138 : OAI22_X1 port map( A1 => n10961, A2 => n8596, B1 => n8622, B2 => 
                           n8594, ZN => n1219);
   U1139 : OAI22_X1 port map( A1 => n10434, A2 => n8596, B1 => n8623, B2 => 
                           n8594, ZN => n1218);
   U1140 : OAI22_X1 port map( A1 => n10435, A2 => n8596, B1 => n8624, B2 => 
                           n8594, ZN => n1217);
   U1141 : OAI22_X1 port map( A1 => n11202, A2 => n8596, B1 => n8626, B2 => 
                           n8594, ZN => n1216);
   U1142 : OAI22_X1 port map( A1 => n10704, A2 => n8596, B1 => n8627, B2 => 
                           n8595, ZN => n1215);
   U1143 : OAI22_X1 port map( A1 => n10962, A2 => n8596, B1 => n8628, B2 => 
                           n8595, ZN => n1214);
   U1144 : OAI22_X1 port map( A1 => n11203, A2 => n8596, B1 => n8629, B2 => 
                           n8595, ZN => n1213);
   U1145 : OAI22_X1 port map( A1 => n10963, A2 => n8596, B1 => n8630, B2 => 
                           n8595, ZN => n1212);
   U1146 : OAI22_X1 port map( A1 => n10436, A2 => n8596, B1 => n8631, B2 => 
                           n8595, ZN => n1211);
   U1147 : OAI22_X1 port map( A1 => n10964, A2 => n8596, B1 => n8632, B2 => 
                           n8595, ZN => n1210);
   U1148 : OAI22_X1 port map( A1 => n11204, A2 => n8596, B1 => n8633, B2 => 
                           n8595, ZN => n1209);
   U1149 : OAI22_X1 port map( A1 => n10705, A2 => n8596, B1 => n8634, B2 => 
                           n8595, ZN => n1208);
   U1150 : OAI22_X1 port map( A1 => n10965, A2 => n8596, B1 => n8636, B2 => 
                           n8595, ZN => n1207);
   U1151 : NAND2_X1 port map( A1 => n8597, A2 => n8601, ZN => n8598);
   U1152 : CLKBUF_X1 port map( A => n8598, Z => n8599);
   U1153 : OAI22_X1 port map( A1 => n10721, A2 => n8600, B1 => n8603, B2 => 
                           n8599, ZN => n1206);
   U1154 : OAI22_X1 port map( A1 => n11205, A2 => n8600, B1 => n8604, B2 => 
                           n8598, ZN => n1205);
   U1155 : OAI22_X1 port map( A1 => n10966, A2 => n8600, B1 => n8605, B2 => 
                           n8599, ZN => n1204);
   U1156 : OAI22_X1 port map( A1 => n10967, A2 => n8600, B1 => n8606, B2 => 
                           n8598, ZN => n1203);
   U1157 : OAI22_X1 port map( A1 => n10968, A2 => n8600, B1 => n8607, B2 => 
                           n8599, ZN => n1202);
   U1158 : OAI22_X1 port map( A1 => n11206, A2 => n8600, B1 => n8608, B2 => 
                           n8598, ZN => n1201);
   U1159 : OAI22_X1 port map( A1 => n10969, A2 => n8600, B1 => n8609, B2 => 
                           n8599, ZN => n1200);
   U1160 : OAI22_X1 port map( A1 => n10970, A2 => n8600, B1 => n8610, B2 => 
                           n8598, ZN => n1199);
   U1161 : OAI22_X1 port map( A1 => n10971, A2 => n8600, B1 => n8611, B2 => 
                           n8599, ZN => n1198);
   U1162 : OAI22_X1 port map( A1 => n11207, A2 => n8600, B1 => n8612, B2 => 
                           n8598, ZN => n1197);
   U1163 : OAI22_X1 port map( A1 => n11208, A2 => n8600, B1 => n8613, B2 => 
                           n8598, ZN => n1196);
   U1164 : OAI22_X1 port map( A1 => n11209, A2 => n8600, B1 => n8614, B2 => 
                           n8599, ZN => n1195);
   U1165 : OAI22_X1 port map( A1 => n11210, A2 => n8600, B1 => n8615, B2 => 
                           n8598, ZN => n1194);
   U1166 : OAI22_X1 port map( A1 => n10972, A2 => n8600, B1 => n8616, B2 => 
                           n8599, ZN => n1193);
   U1167 : OAI22_X1 port map( A1 => n11211, A2 => n8600, B1 => n8617, B2 => 
                           n8598, ZN => n1192);
   U1168 : OAI22_X1 port map( A1 => n10973, A2 => n8600, B1 => n8618, B2 => 
                           n8599, ZN => n1191);
   U1169 : OAI22_X1 port map( A1 => n11212, A2 => n8600, B1 => n8619, B2 => 
                           n8598, ZN => n1190);
   U1170 : OAI22_X1 port map( A1 => n10974, A2 => n8600, B1 => n8620, B2 => 
                           n8598, ZN => n1189);
   U1171 : OAI22_X1 port map( A1 => n10975, A2 => n8600, B1 => n8621, B2 => 
                           n8598, ZN => n1188);
   U1172 : OAI22_X1 port map( A1 => n11213, A2 => n8600, B1 => n8622, B2 => 
                           n8598, ZN => n1187);
   U1173 : OAI22_X1 port map( A1 => n11214, A2 => n8600, B1 => n8623, B2 => 
                           n8598, ZN => n1186);
   U1174 : OAI22_X1 port map( A1 => n10976, A2 => n8600, B1 => n8624, B2 => 
                           n8598, ZN => n1185);
   U1175 : OAI22_X1 port map( A1 => n10977, A2 => n8600, B1 => n8626, B2 => 
                           n8598, ZN => n1184);
   U1176 : OAI22_X1 port map( A1 => n11215, A2 => n8600, B1 => n8627, B2 => 
                           n8599, ZN => n1183);
   U1177 : OAI22_X1 port map( A1 => n11216, A2 => n8600, B1 => n8628, B2 => 
                           n8599, ZN => n1182);
   U1178 : OAI22_X1 port map( A1 => n10978, A2 => n8600, B1 => n8629, B2 => 
                           n8599, ZN => n1181);
   U1179 : OAI22_X1 port map( A1 => n10979, A2 => n8600, B1 => n8630, B2 => 
                           n8599, ZN => n1180);
   U1180 : OAI22_X1 port map( A1 => n10980, A2 => n8600, B1 => n8631, B2 => 
                           n8599, ZN => n1179);
   U1181 : OAI22_X1 port map( A1 => n11217, A2 => n8600, B1 => n8632, B2 => 
                           n8599, ZN => n1178);
   U1182 : OAI22_X1 port map( A1 => n11218, A2 => n8600, B1 => n8633, B2 => 
                           n8599, ZN => n1177);
   U1183 : OAI22_X1 port map( A1 => n10981, A2 => n8600, B1 => n8634, B2 => 
                           n8599, ZN => n1176);
   U1184 : OAI22_X1 port map( A1 => n11219, A2 => n8600, B1 => n8636, B2 => 
                           n8599, ZN => n1175);
   U1185 : NAND2_X1 port map( A1 => n8602, A2 => n8601, ZN => n8625);
   U1186 : CLKBUF_X1 port map( A => n8625, Z => n8635);
   U1187 : OAI22_X1 port map( A1 => n10205, A2 => n8637, B1 => n8603, B2 => 
                           n8635, ZN => n1174);
   U1188 : OAI22_X1 port map( A1 => n10437, A2 => n8637, B1 => n8604, B2 => 
                           n8625, ZN => n1173);
   U1189 : OAI22_X1 port map( A1 => n10982, A2 => n8637, B1 => n8605, B2 => 
                           n8635, ZN => n1172);
   U1190 : OAI22_X1 port map( A1 => n10706, A2 => n8637, B1 => n8606, B2 => 
                           n8625, ZN => n1171);
   U1191 : OAI22_X1 port map( A1 => n10707, A2 => n8637, B1 => n8607, B2 => 
                           n8635, ZN => n1170);
   U1192 : OAI22_X1 port map( A1 => n10438, A2 => n8637, B1 => n8608, B2 => 
                           n8625, ZN => n1169);
   U1193 : OAI22_X1 port map( A1 => n10439, A2 => n8637, B1 => n8609, B2 => 
                           n8635, ZN => n1168);
   U1194 : OAI22_X1 port map( A1 => n10983, A2 => n8637, B1 => n8610, B2 => 
                           n8625, ZN => n1167);
   U1195 : OAI22_X1 port map( A1 => n11220, A2 => n8637, B1 => n8611, B2 => 
                           n8635, ZN => n1166);
   U1196 : OAI22_X1 port map( A1 => n10708, A2 => n8637, B1 => n8612, B2 => 
                           n8625, ZN => n1165);
   U1197 : OAI22_X1 port map( A1 => n10709, A2 => n8637, B1 => n8613, B2 => 
                           n8625, ZN => n1164);
   U1198 : OAI22_X1 port map( A1 => n10984, A2 => n8637, B1 => n8614, B2 => 
                           n8635, ZN => n1163);
   U1199 : OAI22_X1 port map( A1 => n10440, A2 => n8637, B1 => n8615, B2 => 
                           n8625, ZN => n1162);
   U1200 : OAI22_X1 port map( A1 => n10441, A2 => n8637, B1 => n8616, B2 => 
                           n8635, ZN => n1161);
   U1201 : OAI22_X1 port map( A1 => n11221, A2 => n8637, B1 => n8617, B2 => 
                           n8625, ZN => n1160);
   U1202 : OAI22_X1 port map( A1 => n11222, A2 => n8637, B1 => n8618, B2 => 
                           n8635, ZN => n1159);
   U1203 : OAI22_X1 port map( A1 => n10710, A2 => n8637, B1 => n8619, B2 => 
                           n8625, ZN => n1158);
   U1204 : OAI22_X1 port map( A1 => n10442, A2 => n8637, B1 => n8620, B2 => 
                           n8625, ZN => n1157);
   U1205 : OAI22_X1 port map( A1 => n10711, A2 => n8637, B1 => n8621, B2 => 
                           n8625, ZN => n1156);
   U1206 : OAI22_X1 port map( A1 => n10443, A2 => n8637, B1 => n8622, B2 => 
                           n8625, ZN => n1155);
   U1207 : OAI22_X1 port map( A1 => n10712, A2 => n8637, B1 => n8623, B2 => 
                           n8625, ZN => n1154);
   U1208 : OAI22_X1 port map( A1 => n10713, A2 => n8637, B1 => n8624, B2 => 
                           n8625, ZN => n1153);
   U1209 : OAI22_X1 port map( A1 => n10714, A2 => n8637, B1 => n8626, B2 => 
                           n8625, ZN => n1152);
   U1210 : OAI22_X1 port map( A1 => n10985, A2 => n8637, B1 => n8627, B2 => 
                           n8635, ZN => n1151);
   U1211 : OAI22_X1 port map( A1 => n11223, A2 => n8637, B1 => n8628, B2 => 
                           n8635, ZN => n1150);
   U1212 : OAI22_X1 port map( A1 => n10715, A2 => n8637, B1 => n8629, B2 => 
                           n8635, ZN => n1149);
   U1213 : OAI22_X1 port map( A1 => n10986, A2 => n8637, B1 => n8630, B2 => 
                           n8635, ZN => n1148);
   U1214 : OAI22_X1 port map( A1 => n10716, A2 => n8637, B1 => n8631, B2 => 
                           n8635, ZN => n1147);
   U1215 : OAI22_X1 port map( A1 => n10444, A2 => n8637, B1 => n8632, B2 => 
                           n8635, ZN => n1146);
   U1216 : OAI22_X1 port map( A1 => n10717, A2 => n8637, B1 => n8633, B2 => 
                           n8635, ZN => n1145);
   U1217 : OAI22_X1 port map( A1 => n11224, A2 => n8637, B1 => n8634, B2 => 
                           n8635, ZN => n1144);
   U1218 : OAI22_X1 port map( A1 => n11225, A2 => n8637, B1 => n8636, B2 => 
                           n8635, ZN => n1143);
   U1219 : NAND3_X1 port map( A1 => n8451, A2 => ENABLE, A3 => RD2, ZN => n9419
                           );
   U1220 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n8646);
   U1221 : INV_X1 port map( A => ADD_RD2(0), ZN => n8645);
   U1222 : INV_X1 port map( A => ADD_RD2(2), ZN => n8639);
   U1223 : NAND3_X1 port map( A1 => ADD_RD2(1), A2 => n8645, A3 => n8639, ZN =>
                           n8655);
   U1224 : NOR2_X1 port map( A1 => n8646, A2 => n8655, ZN => n9120);
   U1225 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(1), ZN => n8659);
   U1226 : NOR2_X1 port map( A1 => n8646, A2 => n8659, ZN => n9307);
   U1227 : CLKBUF_X1 port map( A => n9307, Z => n9381);
   U1228 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n9120, B1 => 
                           REGISTERS_31_31_port, B2 => n9381, ZN => n8643);
   U1229 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), ZN => n8638);
   U1230 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n8638, ZN => n8661);
   U1231 : NOR2_X1 port map( A1 => n8646, A2 => n8661, ZN => n9077);
   U1232 : NAND2_X1 port map( A1 => n8638, A2 => n8645, ZN => n8657);
   U1233 : NOR2_X1 port map( A1 => n8646, A2 => n8657, ZN => n9071);
   U1234 : CLKBUF_X1 port map( A => n9071, Z => n9372);
   U1235 : AOI22_X1 port map( A1 => REGISTERS_25_31_port, A2 => n9077, B1 => 
                           REGISTERS_24_31_port, B2 => n9372, ZN => n8642);
   U1236 : INV_X1 port map( A => ADD_RD2(3), ZN => n8666);
   U1237 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => n8666, ZN => n8647);
   U1238 : NOR2_X1 port map( A1 => n8647, A2 => n8655, ZN => n9379);
   U1239 : NOR2_X1 port map( A1 => n8647, A2 => n8661, ZN => n9378);
   U1240 : AOI22_X1 port map( A1 => REGISTERS_18_31_port, A2 => n9379, B1 => 
                           REGISTERS_17_31_port, B2 => n9378, ZN => n8641);
   U1241 : NOR2_X1 port map( A1 => n8647, A2 => n8657, ZN => n9076);
   U1242 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), A3 => n8639, 
                           ZN => n8658);
   U1243 : NOR2_X1 port map( A1 => n8646, A2 => n8658, ZN => n9144);
   U1244 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n9076, B1 => 
                           REGISTERS_27_31_port, B2 => n9144, ZN => n8640);
   U1245 : NAND4_X1 port map( A1 => n8643, A2 => n8642, A3 => n8641, A4 => 
                           n8640, ZN => n8653);
   U1246 : INV_X1 port map( A => ADD_RD2(1), ZN => n8644);
   U1247 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(0), A3 => n8644, 
                           ZN => n8656);
   U1248 : NOR2_X1 port map( A1 => n8647, A2 => n8656, ZN => n9368);
   U1249 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(1), A3 => n8645, 
                           ZN => n8660);
   U1250 : NOR2_X1 port map( A1 => n8660, A2 => n8647, ZN => n9312);
   U1251 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n9368, B1 => 
                           REGISTERS_22_31_port, B2 => n9312, ZN => n8651);
   U1252 : NOR2_X1 port map( A1 => n8646, A2 => n8660, ZN => n9369);
   U1253 : NAND3_X1 port map( A1 => ADD_RD2(2), A2 => n8645, A3 => n8644, ZN =>
                           n8654);
   U1254 : NOR2_X1 port map( A1 => n8646, A2 => n8654, ZN => n9121);
   U1255 : AOI22_X1 port map( A1 => REGISTERS_30_31_port, A2 => n9369, B1 => 
                           REGISTERS_28_31_port, B2 => n9121, ZN => n8650);
   U1256 : NOR2_X1 port map( A1 => n8646, A2 => n8656, ZN => n9342);
   U1257 : NOR2_X1 port map( A1 => n8647, A2 => n8659, ZN => n9261);
   U1258 : CLKBUF_X1 port map( A => n9261, Z => n9370);
   U1259 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n9342, B1 => 
                           REGISTERS_23_31_port, B2 => n9370, ZN => n8649);
   U1260 : NOR2_X1 port map( A1 => n8647, A2 => n8658, ZN => n9343);
   U1261 : NOR2_X1 port map( A1 => n8654, A2 => n8647, ZN => n9382);
   U1262 : CLKBUF_X1 port map( A => n9382, Z => n9337);
   U1263 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n9343, B1 => 
                           REGISTERS_20_31_port, B2 => n9337, ZN => n8648);
   U1264 : NAND4_X1 port map( A1 => n8651, A2 => n8650, A3 => n8649, A4 => 
                           n8648, ZN => n8652);
   U1265 : NOR2_X1 port map( A1 => n8653, A2 => n8652, ZN => n8674);
   U1266 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n9365, 
                           ZN => n9416);
   U1267 : CLKBUF_X1 port map( A => n9416, Z => n9234);
   U1268 : INV_X1 port map( A => n8654, ZN => n9201);
   U1269 : INV_X1 port map( A => n8655, ZN => n9322);
   U1270 : CLKBUF_X1 port map( A => n9322, Z => n9110);
   U1271 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_31_port, B1 => 
                           n9110, B2 => REGISTERS_2_31_port, ZN => n8665);
   U1272 : INV_X1 port map( A => n8656, ZN => n9319);
   U1273 : CLKBUF_X1 port map( A => n9319, Z => n9404);
   U1274 : INV_X1 port map( A => n8657, ZN => n9407);
   U1275 : CLKBUF_X1 port map( A => n9407, Z => n9327);
   U1276 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_31_port, B1 => 
                           n9327, B2 => REGISTERS_0_31_port, ZN => n8664);
   U1277 : INV_X1 port map( A => n8658, ZN => n9294);
   U1278 : INV_X1 port map( A => n8659, ZN => n9395);
   U1279 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_3_31_port, B1 => 
                           n9395, B2 => REGISTERS_7_31_port, ZN => n8663);
   U1280 : INV_X1 port map( A => n8660, ZN => n9321);
   U1281 : CLKBUF_X1 port map( A => n9321, Z => n9111);
   U1282 : INV_X1 port map( A => n8661, ZN => n9394);
   U1283 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_31_port, B1 => 
                           n9394, B2 => REGISTERS_1_31_port, ZN => n8662);
   U1284 : NAND4_X1 port map( A1 => n8665, A2 => n8664, A3 => n8663, A4 => 
                           n8662, ZN => n8672);
   U1285 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => n8666, A3 => n9365, ZN => 
                           n9414);
   U1286 : CLKBUF_X1 port map( A => n9414, Z => n9256);
   U1287 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_31_port, B1 => 
                           n9394, B2 => REGISTERS_9_31_port, ZN => n8670);
   U1288 : CLKBUF_X1 port map( A => n9395, Z => n9351);
   U1289 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_31_port, B1 => 
                           n9351, B2 => REGISTERS_15_31_port, ZN => n8669);
   U1290 : CLKBUF_X1 port map( A => n9201, Z => n9401);
   U1291 : CLKBUF_X1 port map( A => n9407, Z => n9392);
   U1292 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_31_port, B1 => 
                           n9392, B2 => REGISTERS_8_31_port, ZN => n8668);
   U1293 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_11_31_port, B1 => 
                           n9110, B2 => REGISTERS_10_31_port, ZN => n8667);
   U1294 : NAND4_X1 port map( A1 => n8670, A2 => n8669, A3 => n8668, A4 => 
                           n8667, ZN => n8671);
   U1295 : AOI22_X1 port map( A1 => n9234, A2 => n8672, B1 => n9256, B2 => 
                           n8671, ZN => n8673);
   U1296 : OAI21_X1 port map( B1 => n9365, B2 => n8674, A => n8673, ZN => N448)
                           ;
   U1297 : CLKBUF_X1 port map( A => n9379, Z => n9336);
   U1298 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_30_port, B1 => 
                           n9336, B2 => REGISTERS_18_30_port, ZN => n8678);
   U1299 : CLKBUF_X1 port map( A => n9369, Z => n9167);
   U1300 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_30_port, B1 => 
                           n9307, B2 => REGISTERS_31_30_port, ZN => n8677);
   U1301 : CLKBUF_X1 port map( A => n9368, Z => n9344);
   U1302 : CLKBUF_X1 port map( A => n9076, Z => n9366);
   U1303 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_30_port, B1 => 
                           n9366, B2 => REGISTERS_16_30_port, ZN => n8676);
   U1304 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_30_port, B1 => 
                           n9372, B2 => REGISTERS_24_30_port, ZN => n8675);
   U1305 : NAND4_X1 port map( A1 => n8678, A2 => n8677, A3 => n8676, A4 => 
                           n8675, ZN => n8684);
   U1306 : CLKBUF_X1 port map( A => n9343, Z => n9383);
   U1307 : CLKBUF_X1 port map( A => n9120, Z => n9384);
   U1308 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_30_port, B1 => 
                           n9384, B2 => REGISTERS_26_30_port, ZN => n8682);
   U1309 : AOI22_X1 port map( A1 => n9312, A2 => REGISTERS_22_30_port, B1 => 
                           n9342, B2 => REGISTERS_29_30_port, ZN => n8681);
   U1310 : CLKBUF_X1 port map( A => n9077, Z => n9373);
   U1311 : CLKBUF_X1 port map( A => n9144, Z => n9380);
   U1312 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_30_port, B1 => 
                           n9380, B2 => REGISTERS_27_30_port, ZN => n8680);
   U1313 : CLKBUF_X1 port map( A => n9378, Z => n9172);
   U1314 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_30_port, B1 => 
                           n9172, B2 => REGISTERS_17_30_port, ZN => n8679);
   U1315 : NAND4_X1 port map( A1 => n8682, A2 => n8681, A3 => n8680, A4 => 
                           n8679, ZN => n8683);
   U1316 : NOR2_X1 port map( A1 => n8684, A2 => n8683, ZN => n8696);
   U1317 : CLKBUF_X1 port map( A => n9319, Z => n9356);
   U1318 : CLKBUF_X1 port map( A => n9394, Z => n9320);
   U1319 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_5_30_port, B1 => 
                           n9320, B2 => REGISTERS_1_30_port, ZN => n8688);
   U1320 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_3_30_port, B1 => 
                           n9392, B2 => REGISTERS_0_30_port, ZN => n8687);
   U1321 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_30_port, B1 => 
                           n9110, B2 => REGISTERS_2_30_port, ZN => n8686);
   U1322 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_30_port, B1 => 
                           n9351, B2 => REGISTERS_7_30_port, ZN => n8685);
   U1323 : NAND4_X1 port map( A1 => n8688, A2 => n8687, A3 => n8686, A4 => 
                           n8685, ZN => n8694);
   U1324 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_30_port, B1 => 
                           n9320, B2 => REGISTERS_9_30_port, ZN => n8692);
   U1325 : CLKBUF_X1 port map( A => n9395, Z => n9408);
   U1326 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_30_port, B1 => 
                           n9392, B2 => REGISTERS_8_30_port, ZN => n8691);
   U1327 : CLKBUF_X1 port map( A => n9294, Z => n9403);
   U1328 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_12_30_port, B1 => 
                           n9403, B2 => REGISTERS_11_30_port, ZN => n8690);
   U1329 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_30_port, B1 => 
                           n9110, B2 => REGISTERS_10_30_port, ZN => n8689);
   U1330 : NAND4_X1 port map( A1 => n8692, A2 => n8691, A3 => n8690, A4 => 
                           n8689, ZN => n8693);
   U1331 : AOI22_X1 port map( A1 => n9234, A2 => n8694, B1 => n9256, B2 => 
                           n8693, ZN => n8695);
   U1332 : OAI21_X1 port map( B1 => n9365, B2 => n8696, A => n8695, ZN => N447)
                           ;
   U1333 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_29_port, B1 => 
                           n9120, B2 => REGISTERS_26_29_port, ZN => n8700);
   U1334 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_29_port, B1 => 
                           n9368, B2 => REGISTERS_21_29_port, ZN => n8699);
   U1335 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_29_port, B1 => 
                           n9342, B2 => REGISTERS_29_29_port, ZN => n8698);
   U1336 : AOI22_X1 port map( A1 => n9312, A2 => REGISTERS_22_29_port, B1 => 
                           n9071, B2 => REGISTERS_24_29_port, ZN => n8697);
   U1337 : NAND4_X1 port map( A1 => n8700, A2 => n8699, A3 => n8698, A4 => 
                           n8697, ZN => n8706);
   U1338 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_29_port, B1 => 
                           n9076, B2 => REGISTERS_16_29_port, ZN => n8704);
   U1339 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_29_port, B1 => 
                           n9144, B2 => REGISTERS_27_29_port, ZN => n8703);
   U1340 : AOI22_X1 port map( A1 => n9307, A2 => REGISTERS_31_29_port, B1 => 
                           n9172, B2 => REGISTERS_17_29_port, ZN => n8702);
   U1341 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_29_port, B1 => 
                           n9379, B2 => REGISTERS_18_29_port, ZN => n8701);
   U1342 : NAND4_X1 port map( A1 => n8704, A2 => n8703, A3 => n8702, A4 => 
                           n8701, ZN => n8705);
   U1343 : NOR2_X1 port map( A1 => n8706, A2 => n8705, ZN => n8718);
   U1344 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_3_29_port, B1 => 
                           n9351, B2 => REGISTERS_7_29_port, ZN => n8710);
   U1345 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_4_29_port, B1 => 
                           n9320, B2 => REGISTERS_1_29_port, ZN => n8709);
   U1346 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_0_29_port, B1 => 
                           n9110, B2 => REGISTERS_2_29_port, ZN => n8708);
   U1347 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_29_port, B1 => 
                           n9356, B2 => REGISTERS_5_29_port, ZN => n8707);
   U1348 : NAND4_X1 port map( A1 => n8710, A2 => n8709, A3 => n8708, A4 => 
                           n8707, ZN => n8716);
   U1349 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_29_port, B1 => 
                           n9356, B2 => REGISTERS_13_29_port, ZN => n8714);
   U1350 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_29_port, B1 => 
                           n9403, B2 => REGISTERS_11_29_port, ZN => n8713);
   U1351 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_29_port, B1 => 
                           n9320, B2 => REGISTERS_9_29_port, ZN => n8712);
   U1352 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_8_29_port, B1 => 
                           n9110, B2 => REGISTERS_10_29_port, ZN => n8711);
   U1353 : NAND4_X1 port map( A1 => n8714, A2 => n8713, A3 => n8712, A4 => 
                           n8711, ZN => n8715);
   U1354 : AOI22_X1 port map( A1 => n9234, A2 => n8716, B1 => n9256, B2 => 
                           n8715, ZN => n8717);
   U1355 : OAI21_X1 port map( B1 => n9365, B2 => n8718, A => n8717, ZN => N446)
                           ;
   U1356 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_28_port, B1 => 
                           n9144, B2 => REGISTERS_27_28_port, ZN => n8722);
   U1357 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_28_port, B1 => 
                           n9379, B2 => REGISTERS_18_28_port, ZN => n8721);
   U1358 : AOI22_X1 port map( A1 => n9312, A2 => REGISTERS_22_28_port, B1 => 
                           n9370, B2 => REGISTERS_23_28_port, ZN => n8720);
   U1359 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_28_port, B1 => 
                           n9172, B2 => REGISTERS_17_28_port, ZN => n8719);
   U1360 : NAND4_X1 port map( A1 => n8722, A2 => n8721, A3 => n8720, A4 => 
                           n8719, ZN => n8728);
   U1361 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_28_port, B1 => 
                           n9343, B2 => REGISTERS_19_28_port, ZN => n8726);
   U1362 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_28_port, B1 => 
                           n9076, B2 => REGISTERS_16_28_port, ZN => n8725);
   U1363 : AOI22_X1 port map( A1 => n9384, A2 => REGISTERS_26_28_port, B1 => 
                           n9307, B2 => REGISTERS_31_28_port, ZN => n8724);
   U1364 : AOI22_X1 port map( A1 => n9368, A2 => REGISTERS_21_28_port, B1 => 
                           n9342, B2 => REGISTERS_29_28_port, ZN => n8723);
   U1365 : NAND4_X1 port map( A1 => n8726, A2 => n8725, A3 => n8724, A4 => 
                           n8723, ZN => n8727);
   U1366 : NOR2_X1 port map( A1 => n8728, A2 => n8727, ZN => n8740);
   U1367 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_28_port, B1 => 
                           n9356, B2 => REGISTERS_5_28_port, ZN => n8732);
   U1368 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_4_28_port, B1 => 
                           n9351, B2 => REGISTERS_7_28_port, ZN => n8731);
   U1369 : AOI22_X1 port map( A1 => n9403, A2 => REGISTERS_3_28_port, B1 => 
                           n9320, B2 => REGISTERS_1_28_port, ZN => n8730);
   U1370 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_0_28_port, B1 => 
                           n9110, B2 => REGISTERS_2_28_port, ZN => n8729);
   U1371 : NAND4_X1 port map( A1 => n8732, A2 => n8731, A3 => n8730, A4 => 
                           n8729, ZN => n8738);
   U1372 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_28_port, B1 => 
                           n9394, B2 => REGISTERS_9_28_port, ZN => n8736);
   U1373 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_12_28_port, B1 => 
                           n9392, B2 => REGISTERS_8_28_port, ZN => n8735);
   U1374 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_28_port, B1 => 
                           n9110, B2 => REGISTERS_10_28_port, ZN => n8734);
   U1375 : AOI22_X1 port map( A1 => n9403, A2 => REGISTERS_11_28_port, B1 => 
                           n9351, B2 => REGISTERS_15_28_port, ZN => n8733);
   U1376 : NAND4_X1 port map( A1 => n8736, A2 => n8735, A3 => n8734, A4 => 
                           n8733, ZN => n8737);
   U1377 : AOI22_X1 port map( A1 => n9234, A2 => n8738, B1 => n9256, B2 => 
                           n8737, ZN => n8739);
   U1378 : OAI21_X1 port map( B1 => n9365, B2 => n8740, A => n8739, ZN => N445)
                           ;
   U1379 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_27_port, B1 => 
                           n9120, B2 => REGISTERS_26_27_port, ZN => n8744);
   U1380 : AOI22_X1 port map( A1 => n9144, A2 => REGISTERS_27_27_port, B1 => 
                           n9379, B2 => REGISTERS_18_27_port, ZN => n8743);
   U1381 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_27_port, B1 => 
                           n9076, B2 => REGISTERS_16_27_port, ZN => n8742);
   U1382 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_27_port, B1 => 
                           n9342, B2 => REGISTERS_29_27_port, ZN => n8741);
   U1383 : NAND4_X1 port map( A1 => n8744, A2 => n8743, A3 => n8742, A4 => 
                           n8741, ZN => n8750);
   U1384 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_27_port, B1 => 
                           n9307, B2 => REGISTERS_31_27_port, ZN => n8748);
   U1385 : AOI22_X1 port map( A1 => n9312, A2 => REGISTERS_22_27_port, B1 => 
                           n9172, B2 => REGISTERS_17_27_port, ZN => n8747);
   U1386 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_27_port, B1 => 
                           n9373, B2 => REGISTERS_25_27_port, ZN => n8746);
   U1387 : AOI22_X1 port map( A1 => n9368, A2 => REGISTERS_21_27_port, B1 => 
                           n9071, B2 => REGISTERS_24_27_port, ZN => n8745);
   U1388 : NAND4_X1 port map( A1 => n8748, A2 => n8747, A3 => n8746, A4 => 
                           n8745, ZN => n8749);
   U1389 : NOR2_X1 port map( A1 => n8750, A2 => n8749, ZN => n8762);
   U1390 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_5_27_port, B1 => 
                           n9392, B2 => REGISTERS_0_27_port, ZN => n8754);
   U1391 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_27_port, B1 => 
                           n9320, B2 => REGISTERS_1_27_port, ZN => n8753);
   U1392 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_27_port, B1 => 
                           n9294, B2 => REGISTERS_3_27_port, ZN => n8752);
   U1393 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_7_27_port, B1 => 
                           n9110, B2 => REGISTERS_2_27_port, ZN => n8751);
   U1394 : NAND4_X1 port map( A1 => n8754, A2 => n8753, A3 => n8752, A4 => 
                           n8751, ZN => n8760);
   U1395 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_27_port, B1 => 
                           n9395, B2 => REGISTERS_15_27_port, ZN => n8758);
   U1396 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_8_27_port, B1 => 
                           n9110, B2 => REGISTERS_10_27_port, ZN => n8757);
   U1397 : CLKBUF_X1 port map( A => n9294, Z => n9396);
   U1398 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_27_port, B1 => 
                           n9394, B2 => REGISTERS_9_27_port, ZN => n8756);
   U1399 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_27_port, B1 => 
                           n9319, B2 => REGISTERS_13_27_port, ZN => n8755);
   U1400 : NAND4_X1 port map( A1 => n8758, A2 => n8757, A3 => n8756, A4 => 
                           n8755, ZN => n8759);
   U1401 : AOI22_X1 port map( A1 => n9234, A2 => n8760, B1 => n9256, B2 => 
                           n8759, ZN => n8761);
   U1402 : OAI21_X1 port map( B1 => n9365, B2 => n8762, A => n8761, ZN => N444)
                           ;
   U1403 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_26_port, B1 => 
                           n9381, B2 => REGISTERS_31_26_port, ZN => n8766);
   U1404 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_26_port, B1 => 
                           n9144, B2 => REGISTERS_27_26_port, ZN => n8765);
   U1405 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_26_port, B1 => 
                           n9342, B2 => REGISTERS_29_26_port, ZN => n8764);
   U1406 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_26_port, B1 => 
                           n9312, B2 => REGISTERS_22_26_port, ZN => n8763);
   U1407 : NAND4_X1 port map( A1 => n8766, A2 => n8765, A3 => n8764, A4 => 
                           n8763, ZN => n8772);
   U1408 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_26_port, B1 => 
                           n9076, B2 => REGISTERS_16_26_port, ZN => n8770);
   U1409 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_26_port, B1 => 
                           n9172, B2 => REGISTERS_17_26_port, ZN => n8769);
   U1410 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_26_port, B1 => 
                           n9120, B2 => REGISTERS_26_26_port, ZN => n8768);
   U1411 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_26_port, B1 => 
                           n9379, B2 => REGISTERS_18_26_port, ZN => n8767);
   U1412 : NAND4_X1 port map( A1 => n8770, A2 => n8769, A3 => n8768, A4 => 
                           n8767, ZN => n8771);
   U1413 : NOR2_X1 port map( A1 => n8772, A2 => n8771, ZN => n8784);
   U1414 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_4_26_port, B1 => 
                           n9351, B2 => REGISTERS_7_26_port, ZN => n8776);
   U1415 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_26_port, B1 => 
                           n9403, B2 => REGISTERS_3_26_port, ZN => n8775);
   U1416 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_5_26_port, B1 => 
                           n9320, B2 => REGISTERS_1_26_port, ZN => n8774);
   U1417 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_0_26_port, B1 => 
                           n9110, B2 => REGISTERS_2_26_port, ZN => n8773);
   U1418 : NAND4_X1 port map( A1 => n8776, A2 => n8775, A3 => n8774, A4 => 
                           n8773, ZN => n8782);
   U1419 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_26_port, B1 => 
                           n9110, B2 => REGISTERS_10_26_port, ZN => n8780);
   U1420 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_26_port, B1 => 
                           n9394, B2 => REGISTERS_9_26_port, ZN => n8779);
   U1421 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_12_26_port, B1 => 
                           n9407, B2 => REGISTERS_8_26_port, ZN => n8778);
   U1422 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_26_port, B1 => 
                           n9395, B2 => REGISTERS_15_26_port, ZN => n8777);
   U1423 : NAND4_X1 port map( A1 => n8780, A2 => n8779, A3 => n8778, A4 => 
                           n8777, ZN => n8781);
   U1424 : AOI22_X1 port map( A1 => n9234, A2 => n8782, B1 => n9256, B2 => 
                           n8781, ZN => n8783);
   U1425 : OAI21_X1 port map( B1 => n9365, B2 => n8784, A => n8783, ZN => N443)
                           ;
   U1426 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_25_port, B1 => 
                           n9120, B2 => REGISTERS_26_25_port, ZN => n8788);
   U1427 : AOI22_X1 port map( A1 => n9312, A2 => REGISTERS_22_25_port, B1 => 
                           n9382, B2 => REGISTERS_20_25_port, ZN => n8787);
   U1428 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_25_port, B1 => 
                           n9261, B2 => REGISTERS_23_25_port, ZN => n8786);
   U1429 : AOI22_X1 port map( A1 => n9366, A2 => REGISTERS_16_25_port, B1 => 
                           n9379, B2 => REGISTERS_18_25_port, ZN => n8785);
   U1430 : NAND4_X1 port map( A1 => n8788, A2 => n8787, A3 => n8786, A4 => 
                           n8785, ZN => n8794);
   U1431 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_25_port, B1 => 
                           n9172, B2 => REGISTERS_17_25_port, ZN => n8792);
   U1432 : AOI22_X1 port map( A1 => n9368, A2 => REGISTERS_21_25_port, B1 => 
                           n9077, B2 => REGISTERS_25_25_port, ZN => n8791);
   U1433 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_25_port, B1 => 
                           n9144, B2 => REGISTERS_27_25_port, ZN => n8790);
   U1434 : CLKBUF_X1 port map( A => n9342, Z => n9371);
   U1435 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_25_port, B1 => 
                           n9381, B2 => REGISTERS_31_25_port, ZN => n8789);
   U1436 : NAND4_X1 port map( A1 => n8792, A2 => n8791, A3 => n8790, A4 => 
                           n8789, ZN => n8793);
   U1437 : NOR2_X1 port map( A1 => n8794, A2 => n8793, ZN => n8806);
   U1438 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_25_port, B1 => 
                           n9392, B2 => REGISTERS_0_25_port, ZN => n8798);
   U1439 : CLKBUF_X1 port map( A => n9201, Z => n9393);
   U1440 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_25_port, B1 => 
                           n9351, B2 => REGISTERS_7_25_port, ZN => n8797);
   U1441 : CLKBUF_X1 port map( A => n9394, Z => n9406);
   U1442 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_25_port, B1 => 
                           n9110, B2 => REGISTERS_2_25_port, ZN => n8796);
   U1443 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_25_port, B1 => 
                           n9294, B2 => REGISTERS_3_25_port, ZN => n8795);
   U1444 : NAND4_X1 port map( A1 => n8798, A2 => n8797, A3 => n8796, A4 => 
                           n8795, ZN => n8804);
   U1445 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_9_25_port, B1 => 
                           n9407, B2 => REGISTERS_8_25_port, ZN => n8802);
   U1446 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_12_25_port, B1 => 
                           n9403, B2 => REGISTERS_11_25_port, ZN => n8801);
   U1447 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_13_25_port, B1 => 
                           n9395, B2 => REGISTERS_15_25_port, ZN => n8800);
   U1448 : CLKBUF_X1 port map( A => n9321, Z => n9402);
   U1449 : CLKBUF_X1 port map( A => n9322, Z => n9405);
   U1450 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_25_port, B1 => 
                           n9405, B2 => REGISTERS_10_25_port, ZN => n8799);
   U1451 : NAND4_X1 port map( A1 => n8802, A2 => n8801, A3 => n8800, A4 => 
                           n8799, ZN => n8803);
   U1452 : AOI22_X1 port map( A1 => n9234, A2 => n8804, B1 => n9256, B2 => 
                           n8803, ZN => n8805);
   U1453 : OAI21_X1 port map( B1 => n9365, B2 => n8806, A => n8805, ZN => N442)
                           ;
   U1454 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_24_port, B1 => 
                           n9379, B2 => REGISTERS_18_24_port, ZN => n8810);
   U1455 : AOI22_X1 port map( A1 => n9368, A2 => REGISTERS_21_24_port, B1 => 
                           n9144, B2 => REGISTERS_27_24_port, ZN => n8809);
   U1456 : CLKBUF_X1 port map( A => n9121, Z => n9385);
   U1457 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_24_port, B1 => 
                           n9172, B2 => REGISTERS_17_24_port, ZN => n8808);
   U1458 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_24_port, B1 => 
                           n9382, B2 => REGISTERS_20_24_port, ZN => n8807);
   U1459 : NAND4_X1 port map( A1 => n8810, A2 => n8809, A3 => n8808, A4 => 
                           n8807, ZN => n8816);
   U1460 : AOI22_X1 port map( A1 => n9307, A2 => REGISTERS_31_24_port, B1 => 
                           n9076, B2 => REGISTERS_16_24_port, ZN => n8814);
   U1461 : AOI22_X1 port map( A1 => n9312, A2 => REGISTERS_22_24_port, B1 => 
                           n9120, B2 => REGISTERS_26_24_port, ZN => n8813);
   U1462 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_24_port, B1 => 
                           n9071, B2 => REGISTERS_24_24_port, ZN => n8812);
   U1463 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_24_port, B1 => 
                           n9077, B2 => REGISTERS_25_24_port, ZN => n8811);
   U1464 : NAND4_X1 port map( A1 => n8814, A2 => n8813, A3 => n8812, A4 => 
                           n8811, ZN => n8815);
   U1465 : NOR2_X1 port map( A1 => n8816, A2 => n8815, ZN => n8828);
   U1466 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_7_24_port, B1 => 
                           n9322, B2 => REGISTERS_2_24_port, ZN => n8820);
   U1467 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_24_port, B1 => 
                           n9392, B2 => REGISTERS_0_24_port, ZN => n8819);
   U1468 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_24_port, B1 => 
                           n9403, B2 => REGISTERS_3_24_port, ZN => n8818);
   U1469 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_24_port, B1 => 
                           n9319, B2 => REGISTERS_5_24_port, ZN => n8817);
   U1470 : NAND4_X1 port map( A1 => n8820, A2 => n8819, A3 => n8818, A4 => 
                           n8817, ZN => n8826);
   U1471 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_13_24_port, B1 => 
                           n9407, B2 => REGISTERS_8_24_port, ZN => n8824);
   U1472 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_24_port, B1 => 
                           n9351, B2 => REGISTERS_15_24_port, ZN => n8823);
   U1473 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_24_port, B1 => 
                           n9320, B2 => REGISTERS_9_24_port, ZN => n8822);
   U1474 : AOI22_X1 port map( A1 => n9403, A2 => REGISTERS_11_24_port, B1 => 
                           n9110, B2 => REGISTERS_10_24_port, ZN => n8821);
   U1475 : NAND4_X1 port map( A1 => n8824, A2 => n8823, A3 => n8822, A4 => 
                           n8821, ZN => n8825);
   U1476 : AOI22_X1 port map( A1 => n9234, A2 => n8826, B1 => n9256, B2 => 
                           n8825, ZN => n8827);
   U1477 : OAI21_X1 port map( B1 => n9365, B2 => n8828, A => n8827, ZN => N441)
                           ;
   U1478 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_23_port, B1 => 
                           n9261, B2 => REGISTERS_23_23_port, ZN => n8832);
   U1479 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_23_port, B1 => 
                           n9373, B2 => REGISTERS_25_23_port, ZN => n8831);
   U1480 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_23_port, B1 => 
                           n9144, B2 => REGISTERS_27_23_port, ZN => n8830);
   U1481 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_23_port, B1 => 
                           n9336, B2 => REGISTERS_18_23_port, ZN => n8829);
   U1482 : NAND4_X1 port map( A1 => n8832, A2 => n8831, A3 => n8830, A4 => 
                           n8829, ZN => n8838);
   U1483 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_23_port, B1 => 
                           n9120, B2 => REGISTERS_26_23_port, ZN => n8836);
   U1484 : CLKBUF_X1 port map( A => n9312, Z => n9367);
   U1485 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_23_port, B1 => 
                           n9172, B2 => REGISTERS_17_23_port, ZN => n8835);
   U1486 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_23_port, B1 => 
                           n9076, B2 => REGISTERS_16_23_port, ZN => n8834);
   U1487 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_23_port, B1 => 
                           n9071, B2 => REGISTERS_24_23_port, ZN => n8833);
   U1488 : NAND4_X1 port map( A1 => n8836, A2 => n8835, A3 => n8834, A4 => 
                           n8833, ZN => n8837);
   U1489 : NOR2_X1 port map( A1 => n8838, A2 => n8837, ZN => n8850);
   U1490 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_23_port, B1 => 
                           n9392, B2 => REGISTERS_0_23_port, ZN => n8842);
   U1491 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_6_23_port, B1 => 
                           n9395, B2 => REGISTERS_7_23_port, ZN => n8841);
   U1492 : AOI22_X1 port map( A1 => n9394, A2 => REGISTERS_1_23_port, B1 => 
                           n9405, B2 => REGISTERS_2_23_port, ZN => n8840);
   U1493 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_23_port, B1 => 
                           n9319, B2 => REGISTERS_5_23_port, ZN => n8839);
   U1494 : NAND4_X1 port map( A1 => n8842, A2 => n8841, A3 => n8840, A4 => 
                           n8839, ZN => n8848);
   U1495 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_11_23_port, B1 => 
                           n9322, B2 => REGISTERS_10_23_port, ZN => n8846);
   U1496 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_9_23_port, B1 => 
                           n9407, B2 => REGISTERS_8_23_port, ZN => n8845);
   U1497 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_23_port, B1 => 
                           n9351, B2 => REGISTERS_15_23_port, ZN => n8844);
   U1498 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_14_23_port, B1 => 
                           n9401, B2 => REGISTERS_12_23_port, ZN => n8843);
   U1499 : NAND4_X1 port map( A1 => n8846, A2 => n8845, A3 => n8844, A4 => 
                           n8843, ZN => n8847);
   U1500 : AOI22_X1 port map( A1 => n9234, A2 => n8848, B1 => n9256, B2 => 
                           n8847, ZN => n8849);
   U1501 : OAI21_X1 port map( B1 => n9419, B2 => n8850, A => n8849, ZN => N440)
                           ;
   U1502 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_22_port, B1 => 
                           n9379, B2 => REGISTERS_18_22_port, ZN => n8854);
   U1503 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_22_port, B1 => 
                           n9382, B2 => REGISTERS_20_22_port, ZN => n8853);
   U1504 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_22_port, B1 => 
                           n9144, B2 => REGISTERS_27_22_port, ZN => n8852);
   U1505 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_22_port, B1 => 
                           n9120, B2 => REGISTERS_26_22_port, ZN => n8851);
   U1506 : NAND4_X1 port map( A1 => n8854, A2 => n8853, A3 => n8852, A4 => 
                           n8851, ZN => n8860);
   U1507 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_22_port, B1 => 
                           n9076, B2 => REGISTERS_16_22_port, ZN => n8858);
   U1508 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_22_port, B1 => 
                           n9172, B2 => REGISTERS_17_22_port, ZN => n8857);
   U1509 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_22_port, B1 => 
                           n9381, B2 => REGISTERS_31_22_port, ZN => n8856);
   U1510 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_22_port, B1 => 
                           n9261, B2 => REGISTERS_23_22_port, ZN => n8855);
   U1511 : NAND4_X1 port map( A1 => n8858, A2 => n8857, A3 => n8856, A4 => 
                           n8855, ZN => n8859);
   U1512 : NOR2_X1 port map( A1 => n8860, A2 => n8859, ZN => n8872);
   U1513 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_22_port, B1 => 
                           n9294, B2 => REGISTERS_3_22_port, ZN => n8864);
   U1514 : AOI22_X1 port map( A1 => n9395, A2 => REGISTERS_7_22_port, B1 => 
                           n9394, B2 => REGISTERS_1_22_port, ZN => n8863);
   U1515 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_4_22_port, B1 => 
                           n9392, B2 => REGISTERS_0_22_port, ZN => n8862);
   U1516 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_5_22_port, B1 => 
                           n9110, B2 => REGISTERS_2_22_port, ZN => n8861);
   U1517 : NAND4_X1 port map( A1 => n8864, A2 => n8863, A3 => n8862, A4 => 
                           n8861, ZN => n8870);
   U1518 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_12_22_port, B1 => 
                           n9405, B2 => REGISTERS_10_22_port, ZN => n8868);
   U1519 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_22_port, B1 => 
                           n9407, B2 => REGISTERS_8_22_port, ZN => n8867);
   U1520 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_22_port, B1 => 
                           n9395, B2 => REGISTERS_15_22_port, ZN => n8866);
   U1521 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_13_22_port, B1 => 
                           n9320, B2 => REGISTERS_9_22_port, ZN => n8865);
   U1522 : NAND4_X1 port map( A1 => n8868, A2 => n8867, A3 => n8866, A4 => 
                           n8865, ZN => n8869);
   U1523 : AOI22_X1 port map( A1 => n9234, A2 => n8870, B1 => n9256, B2 => 
                           n8869, ZN => n8871);
   U1524 : OAI21_X1 port map( B1 => n9419, B2 => n8872, A => n8871, ZN => N439)
                           ;
   U1525 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_21_port, B1 => 
                           n9381, B2 => REGISTERS_31_21_port, ZN => n8876);
   U1526 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_21_port, B1 => 
                           n9382, B2 => REGISTERS_20_21_port, ZN => n8875);
   U1527 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_21_port, B1 => 
                           n9144, B2 => REGISTERS_27_21_port, ZN => n8874);
   U1528 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_21_port, B1 => 
                           n9379, B2 => REGISTERS_18_21_port, ZN => n8873);
   U1529 : NAND4_X1 port map( A1 => n8876, A2 => n8875, A3 => n8874, A4 => 
                           n8873, ZN => n8882);
   U1530 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_21_port, B1 => 
                           n9071, B2 => REGISTERS_24_21_port, ZN => n8880);
   U1531 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_21_port, B1 => 
                           n9378, B2 => REGISTERS_17_21_port, ZN => n8879);
   U1532 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_21_port, B1 => 
                           n9076, B2 => REGISTERS_16_21_port, ZN => n8878);
   U1533 : AOI22_X1 port map( A1 => n9261, A2 => REGISTERS_23_21_port, B1 => 
                           n9120, B2 => REGISTERS_26_21_port, ZN => n8877);
   U1534 : NAND4_X1 port map( A1 => n8880, A2 => n8879, A3 => n8878, A4 => 
                           n8877, ZN => n8881);
   U1535 : NOR2_X1 port map( A1 => n8882, A2 => n8881, ZN => n8894);
   U1536 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_21_port, B1 => 
                           n9392, B2 => REGISTERS_0_21_port, ZN => n8886);
   U1537 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_21_port, B1 => 
                           n9394, B2 => REGISTERS_1_21_port, ZN => n8885);
   U1538 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_21_port, B1 => 
                           n9294, B2 => REGISTERS_3_21_port, ZN => n8884);
   U1539 : AOI22_X1 port map( A1 => n9351, A2 => REGISTERS_7_21_port, B1 => 
                           n9322, B2 => REGISTERS_2_21_port, ZN => n8883);
   U1540 : NAND4_X1 port map( A1 => n8886, A2 => n8885, A3 => n8884, A4 => 
                           n8883, ZN => n8892);
   U1541 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_21_port, B1 => 
                           n9201, B2 => REGISTERS_12_21_port, ZN => n8890);
   U1542 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_21_port, B1 => 
                           n9351, B2 => REGISTERS_15_21_port, ZN => n8889);
   U1543 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_8_21_port, B1 => 
                           n9110, B2 => REGISTERS_10_21_port, ZN => n8888);
   U1544 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_11_21_port, B1 => 
                           n9320, B2 => REGISTERS_9_21_port, ZN => n8887);
   U1545 : NAND4_X1 port map( A1 => n8890, A2 => n8889, A3 => n8888, A4 => 
                           n8887, ZN => n8891);
   U1546 : AOI22_X1 port map( A1 => n9234, A2 => n8892, B1 => n9256, B2 => 
                           n8891, ZN => n8893);
   U1547 : OAI21_X1 port map( B1 => n9419, B2 => n8894, A => n8893, ZN => N438)
                           ;
   U1548 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_20_port, B1 => 
                           n9261, B2 => REGISTERS_23_20_port, ZN => n8898);
   U1549 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_20_port, B1 => 
                           n9380, B2 => REGISTERS_27_20_port, ZN => n8897);
   U1550 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_20_port, B1 => 
                           n9077, B2 => REGISTERS_25_20_port, ZN => n8896);
   U1551 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_20_port, B1 => 
                           n9384, B2 => REGISTERS_26_20_port, ZN => n8895);
   U1552 : NAND4_X1 port map( A1 => n8898, A2 => n8897, A3 => n8896, A4 => 
                           n8895, ZN => n8904);
   U1553 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_20_port, B1 => 
                           n9366, B2 => REGISTERS_16_20_port, ZN => n8902);
   U1554 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_20_port, B1 => 
                           n9378, B2 => REGISTERS_17_20_port, ZN => n8901);
   U1555 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_20_port, B1 => 
                           n9071, B2 => REGISTERS_24_20_port, ZN => n8900);
   U1556 : AOI22_X1 port map( A1 => n9307, A2 => REGISTERS_31_20_port, B1 => 
                           n9336, B2 => REGISTERS_18_20_port, ZN => n8899);
   U1557 : NAND4_X1 port map( A1 => n8902, A2 => n8901, A3 => n8900, A4 => 
                           n8899, ZN => n8903);
   U1558 : NOR2_X1 port map( A1 => n8904, A2 => n8903, ZN => n8916);
   U1559 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_20_port, B1 => 
                           n9405, B2 => REGISTERS_2_20_port, ZN => n8908);
   U1560 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_5_20_port, B1 => 
                           n9395, B2 => REGISTERS_7_20_port, ZN => n8907);
   U1561 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_6_20_port, B1 => 
                           n9407, B2 => REGISTERS_0_20_port, ZN => n8906);
   U1562 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_20_port, B1 => 
                           n9394, B2 => REGISTERS_1_20_port, ZN => n8905);
   U1563 : NAND4_X1 port map( A1 => n8908, A2 => n8907, A3 => n8906, A4 => 
                           n8905, ZN => n8914);
   U1564 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_8_20_port, B1 => 
                           n9322, B2 => REGISTERS_10_20_port, ZN => n8912);
   U1565 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_20_port, B1 => 
                           n9395, B2 => REGISTERS_15_20_port, ZN => n8911);
   U1566 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_14_20_port, B1 => 
                           n9394, B2 => REGISTERS_9_20_port, ZN => n8910);
   U1567 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_20_port, B1 => 
                           n9403, B2 => REGISTERS_11_20_port, ZN => n8909);
   U1568 : NAND4_X1 port map( A1 => n8912, A2 => n8911, A3 => n8910, A4 => 
                           n8909, ZN => n8913);
   U1569 : AOI22_X1 port map( A1 => n9234, A2 => n8914, B1 => n9414, B2 => 
                           n8913, ZN => n8915);
   U1570 : OAI21_X1 port map( B1 => n9419, B2 => n8916, A => n8915, ZN => N437)
                           ;
   U1571 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_19_port, B1 => 
                           n9261, B2 => REGISTERS_23_19_port, ZN => n8920);
   U1572 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_19_port, B1 => 
                           n9384, B2 => REGISTERS_26_19_port, ZN => n8919);
   U1573 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_19_port, B1 => 
                           n9380, B2 => REGISTERS_27_19_port, ZN => n8918);
   U1574 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_19_port, B1 => 
                           n9336, B2 => REGISTERS_18_19_port, ZN => n8917);
   U1575 : NAND4_X1 port map( A1 => n8920, A2 => n8919, A3 => n8918, A4 => 
                           n8917, ZN => n8926);
   U1576 : AOI22_X1 port map( A1 => n9077, A2 => REGISTERS_25_19_port, B1 => 
                           n9366, B2 => REGISTERS_16_19_port, ZN => n8924);
   U1577 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_19_port, B1 => 
                           n9343, B2 => REGISTERS_19_19_port, ZN => n8923);
   U1578 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_19_port, B1 => 
                           n9381, B2 => REGISTERS_31_19_port, ZN => n8922);
   U1579 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_19_port, B1 => 
                           n9172, B2 => REGISTERS_17_19_port, ZN => n8921);
   U1580 : NAND4_X1 port map( A1 => n8924, A2 => n8923, A3 => n8922, A4 => 
                           n8921, ZN => n8925);
   U1581 : NOR2_X1 port map( A1 => n8926, A2 => n8925, ZN => n8938);
   U1582 : CLKBUF_X1 port map( A => n9416, Z => n9258);
   U1583 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_19_port, B1 => 
                           n9407, B2 => REGISTERS_0_19_port, ZN => n8930);
   U1584 : AOI22_X1 port map( A1 => n9395, A2 => REGISTERS_7_19_port, B1 => 
                           n9110, B2 => REGISTERS_2_19_port, ZN => n8929);
   U1585 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_19_port, B1 => 
                           n9403, B2 => REGISTERS_3_19_port, ZN => n8928);
   U1586 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_19_port, B1 => 
                           n9320, B2 => REGISTERS_1_19_port, ZN => n8927);
   U1587 : NAND4_X1 port map( A1 => n8930, A2 => n8929, A3 => n8928, A4 => 
                           n8927, ZN => n8936);
   U1588 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_13_19_port, B1 => 
                           n9351, B2 => REGISTERS_15_19_port, ZN => n8934);
   U1589 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_19_port, B1 => 
                           n9394, B2 => REGISTERS_9_19_port, ZN => n8933);
   U1590 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_12_19_port, B1 => 
                           n9405, B2 => REGISTERS_10_19_port, ZN => n8932);
   U1591 : AOI22_X1 port map( A1 => n9403, A2 => REGISTERS_11_19_port, B1 => 
                           n9392, B2 => REGISTERS_8_19_port, ZN => n8931);
   U1592 : NAND4_X1 port map( A1 => n8934, A2 => n8933, A3 => n8932, A4 => 
                           n8931, ZN => n8935);
   U1593 : AOI22_X1 port map( A1 => n9258, A2 => n8936, B1 => n9256, B2 => 
                           n8935, ZN => n8937);
   U1594 : OAI21_X1 port map( B1 => n9419, B2 => n8938, A => n8937, ZN => N436)
                           ;
   U1595 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_18_port, B1 => 
                           n9380, B2 => REGISTERS_27_18_port, ZN => n8942);
   U1596 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_18_port, B1 => 
                           n9336, B2 => REGISTERS_18_18_port, ZN => n8941);
   U1597 : AOI22_X1 port map( A1 => n9071, A2 => REGISTERS_24_18_port, B1 => 
                           n9172, B2 => REGISTERS_17_18_port, ZN => n8940);
   U1598 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_18_port, B1 => 
                           n9381, B2 => REGISTERS_31_18_port, ZN => n8939);
   U1599 : NAND4_X1 port map( A1 => n8942, A2 => n8941, A3 => n8940, A4 => 
                           n8939, ZN => n8948);
   U1600 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_18_port, B1 => 
                           n9077, B2 => REGISTERS_25_18_port, ZN => n8946);
   U1601 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_18_port, B1 => 
                           n9261, B2 => REGISTERS_23_18_port, ZN => n8945);
   U1602 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_18_port, B1 => 
                           n9366, B2 => REGISTERS_16_18_port, ZN => n8944);
   U1603 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_18_port, B1 => 
                           n9384, B2 => REGISTERS_26_18_port, ZN => n8943);
   U1604 : NAND4_X1 port map( A1 => n8946, A2 => n8945, A3 => n8944, A4 => 
                           n8943, ZN => n8947);
   U1605 : NOR2_X1 port map( A1 => n8948, A2 => n8947, ZN => n8960);
   U1606 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_5_18_port, B1 => 
                           n9395, B2 => REGISTERS_7_18_port, ZN => n8952);
   U1607 : AOI22_X1 port map( A1 => n9320, A2 => REGISTERS_1_18_port, B1 => 
                           n9322, B2 => REGISTERS_2_18_port, ZN => n8951);
   U1608 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_18_port, B1 => 
                           n9294, B2 => REGISTERS_3_18_port, ZN => n8950);
   U1609 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_4_18_port, B1 => 
                           n9407, B2 => REGISTERS_0_18_port, ZN => n8949);
   U1610 : NAND4_X1 port map( A1 => n8952, A2 => n8951, A3 => n8950, A4 => 
                           n8949, ZN => n8958);
   U1611 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_18_port, B1 => 
                           n9392, B2 => REGISTERS_8_18_port, ZN => n8956);
   U1612 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_18_port, B1 => 
                           n9320, B2 => REGISTERS_9_18_port, ZN => n8955);
   U1613 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_18_port, B1 => 
                           n9351, B2 => REGISTERS_15_18_port, ZN => n8954);
   U1614 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_11_18_port, B1 => 
                           n9110, B2 => REGISTERS_10_18_port, ZN => n8953);
   U1615 : NAND4_X1 port map( A1 => n8956, A2 => n8955, A3 => n8954, A4 => 
                           n8953, ZN => n8957);
   U1616 : AOI22_X1 port map( A1 => n9258, A2 => n8958, B1 => n9256, B2 => 
                           n8957, ZN => n8959);
   U1617 : OAI21_X1 port map( B1 => n9419, B2 => n8960, A => n8959, ZN => N435)
                           ;
   U1618 : AOI22_X1 port map( A1 => n9076, A2 => REGISTERS_16_17_port, B1 => 
                           n9380, B2 => REGISTERS_27_17_port, ZN => n8964);
   U1619 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_17_port, B1 => 
                           n9077, B2 => REGISTERS_25_17_port, ZN => n8963);
   U1620 : AOI22_X1 port map( A1 => n9342, A2 => REGISTERS_29_17_port, B1 => 
                           n9261, B2 => REGISTERS_23_17_port, ZN => n8962);
   U1621 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_17_port, B1 => 
                           n9384, B2 => REGISTERS_26_17_port, ZN => n8961);
   U1622 : NAND4_X1 port map( A1 => n8964, A2 => n8963, A3 => n8962, A4 => 
                           n8961, ZN => n8970);
   U1623 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_17_port, B1 => 
                           n9121, B2 => REGISTERS_28_17_port, ZN => n8968);
   U1624 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_17_port, B1 => 
                           n9336, B2 => REGISTERS_18_17_port, ZN => n8967);
   U1625 : AOI22_X1 port map( A1 => n9071, A2 => REGISTERS_24_17_port, B1 => 
                           n9172, B2 => REGISTERS_17_17_port, ZN => n8966);
   U1626 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_17_port, B1 => 
                           n9337, B2 => REGISTERS_20_17_port, ZN => n8965);
   U1627 : NAND4_X1 port map( A1 => n8968, A2 => n8967, A3 => n8966, A4 => 
                           n8965, ZN => n8969);
   U1628 : NOR2_X1 port map( A1 => n8970, A2 => n8969, ZN => n8982);
   U1629 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_17_port, B1 => 
                           n9401, B2 => REGISTERS_4_17_port, ZN => n8974);
   U1630 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_17_port, B1 => 
                           n9407, B2 => REGISTERS_0_17_port, ZN => n8973);
   U1631 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_17_port, B1 => 
                           n9395, B2 => REGISTERS_7_17_port, ZN => n8972);
   U1632 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_17_port, B1 => 
                           n9110, B2 => REGISTERS_2_17_port, ZN => n8971);
   U1633 : NAND4_X1 port map( A1 => n8974, A2 => n8973, A3 => n8972, A4 => 
                           n8971, ZN => n8980);
   U1634 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_13_17_port, B1 => 
                           n9405, B2 => REGISTERS_10_17_port, ZN => n8978);
   U1635 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_17_port, B1 => 
                           n9392, B2 => REGISTERS_8_17_port, ZN => n8977);
   U1636 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_17_port, B1 => 
                           n9403, B2 => REGISTERS_11_17_port, ZN => n8976);
   U1637 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_17_port, B1 => 
                           n9394, B2 => REGISTERS_9_17_port, ZN => n8975);
   U1638 : NAND4_X1 port map( A1 => n8978, A2 => n8977, A3 => n8976, A4 => 
                           n8975, ZN => n8979);
   U1639 : AOI22_X1 port map( A1 => n9258, A2 => n8980, B1 => n9256, B2 => 
                           n8979, ZN => n8981);
   U1640 : OAI21_X1 port map( B1 => n9419, B2 => n8982, A => n8981, ZN => N434)
                           ;
   U1641 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_16_port, B1 => 
                           n9366, B2 => REGISTERS_16_16_port, ZN => n8986);
   U1642 : AOI22_X1 port map( A1 => n9261, A2 => REGISTERS_23_16_port, B1 => 
                           n9384, B2 => REGISTERS_26_16_port, ZN => n8985);
   U1643 : AOI22_X1 port map( A1 => n9342, A2 => REGISTERS_29_16_port, B1 => 
                           n9077, B2 => REGISTERS_25_16_port, ZN => n8984);
   U1644 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_16_port, B1 => 
                           n9368, B2 => REGISTERS_21_16_port, ZN => n8983);
   U1645 : NAND4_X1 port map( A1 => n8986, A2 => n8985, A3 => n8984, A4 => 
                           n8983, ZN => n8992);
   U1646 : AOI22_X1 port map( A1 => n9343, A2 => REGISTERS_19_16_port, B1 => 
                           n9071, B2 => REGISTERS_24_16_port, ZN => n8990);
   U1647 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_16_port, B1 => 
                           n9380, B2 => REGISTERS_27_16_port, ZN => n8989);
   U1648 : AOI22_X1 port map( A1 => n9382, A2 => REGISTERS_20_16_port, B1 => 
                           n9172, B2 => REGISTERS_17_16_port, ZN => n8988);
   U1649 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_16_port, B1 => 
                           n9336, B2 => REGISTERS_18_16_port, ZN => n8987);
   U1650 : NAND4_X1 port map( A1 => n8990, A2 => n8989, A3 => n8988, A4 => 
                           n8987, ZN => n8991);
   U1651 : NOR2_X1 port map( A1 => n8992, A2 => n8991, ZN => n9004);
   U1652 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_5_16_port, B1 => 
                           n9294, B2 => REGISTERS_3_16_port, ZN => n8996);
   U1653 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_16_port, B1 => 
                           n9351, B2 => REGISTERS_7_16_port, ZN => n8995);
   U1654 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_0_16_port, B1 => 
                           n9322, B2 => REGISTERS_2_16_port, ZN => n8994);
   U1655 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_16_port, B1 => 
                           n9320, B2 => REGISTERS_1_16_port, ZN => n8993);
   U1656 : NAND4_X1 port map( A1 => n8996, A2 => n8995, A3 => n8994, A4 => 
                           n8993, ZN => n9002);
   U1657 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_16_port, B1 => 
                           n9407, B2 => REGISTERS_8_16_port, ZN => n9000);
   U1658 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_16_port, B1 => 
                           n9405, B2 => REGISTERS_10_16_port, ZN => n8999);
   U1659 : AOI22_X1 port map( A1 => n9403, A2 => REGISTERS_11_16_port, B1 => 
                           n9395, B2 => REGISTERS_15_16_port, ZN => n8998);
   U1660 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_13_16_port, B1 => 
                           n9394, B2 => REGISTERS_9_16_port, ZN => n8997);
   U1661 : NAND4_X1 port map( A1 => n9000, A2 => n8999, A3 => n8998, A4 => 
                           n8997, ZN => n9001);
   U1662 : AOI22_X1 port map( A1 => n9258, A2 => n9002, B1 => n9256, B2 => 
                           n9001, ZN => n9003);
   U1663 : OAI21_X1 port map( B1 => n9419, B2 => n9004, A => n9003, ZN => N433)
                           ;
   U1664 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_15_port, B1 => 
                           n9384, B2 => REGISTERS_26_15_port, ZN => n9008);
   U1665 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_15_port, B1 => 
                           n9172, B2 => REGISTERS_17_15_port, ZN => n9007);
   U1666 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_15_port, B1 => 
                           n9366, B2 => REGISTERS_16_15_port, ZN => n9006);
   U1667 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_15_port, B1 => 
                           n9343, B2 => REGISTERS_19_15_port, ZN => n9005);
   U1668 : NAND4_X1 port map( A1 => n9008, A2 => n9007, A3 => n9006, A4 => 
                           n9005, ZN => n9014);
   U1669 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_15_port, B1 => 
                           n9381, B2 => REGISTERS_31_15_port, ZN => n9012);
   U1670 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_15_port, B1 => 
                           n9382, B2 => REGISTERS_20_15_port, ZN => n9011);
   U1671 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_15_port, B1 => 
                           n9380, B2 => REGISTERS_27_15_port, ZN => n9010);
   U1672 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_15_port, B1 => 
                           n9336, B2 => REGISTERS_18_15_port, ZN => n9009);
   U1673 : NAND4_X1 port map( A1 => n9012, A2 => n9011, A3 => n9010, A4 => 
                           n9009, ZN => n9013);
   U1674 : NOR2_X1 port map( A1 => n9014, A2 => n9013, ZN => n9026);
   U1675 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_15_port, B1 => 
                           n9407, B2 => REGISTERS_0_15_port, ZN => n9018);
   U1676 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_3_15_port, B1 => 
                           n9110, B2 => REGISTERS_2_15_port, ZN => n9017);
   U1677 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_5_15_port, B1 => 
                           n9351, B2 => REGISTERS_7_15_port, ZN => n9016);
   U1678 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_15_port, B1 => 
                           n9320, B2 => REGISTERS_1_15_port, ZN => n9015);
   U1679 : NAND4_X1 port map( A1 => n9018, A2 => n9017, A3 => n9016, A4 => 
                           n9015, ZN => n9024);
   U1680 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_15_port, B1 => 
                           n9406, B2 => REGISTERS_9_15_port, ZN => n9022);
   U1681 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_15_port, B1 => 
                           n9405, B2 => REGISTERS_10_15_port, ZN => n9021);
   U1682 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_15_port, B1 => 
                           n9201, B2 => REGISTERS_12_15_port, ZN => n9020);
   U1683 : AOI22_X1 port map( A1 => n9351, A2 => REGISTERS_15_15_port, B1 => 
                           n9327, B2 => REGISTERS_8_15_port, ZN => n9019);
   U1684 : NAND4_X1 port map( A1 => n9022, A2 => n9021, A3 => n9020, A4 => 
                           n9019, ZN => n9023);
   U1685 : AOI22_X1 port map( A1 => n9258, A2 => n9024, B1 => n9256, B2 => 
                           n9023, ZN => n9025);
   U1686 : OAI21_X1 port map( B1 => n9365, B2 => n9026, A => n9025, ZN => N432)
                           ;
   U1687 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_14_port, B1 => 
                           n9381, B2 => REGISTERS_31_14_port, ZN => n9030);
   U1688 : AOI22_X1 port map( A1 => n9343, A2 => REGISTERS_19_14_port, B1 => 
                           n9371, B2 => REGISTERS_29_14_port, ZN => n9029);
   U1689 : AOI22_X1 port map( A1 => n9077, A2 => REGISTERS_25_14_port, B1 => 
                           n9071, B2 => REGISTERS_24_14_port, ZN => n9028);
   U1690 : AOI22_X1 port map( A1 => n9382, A2 => REGISTERS_20_14_port, B1 => 
                           n9172, B2 => REGISTERS_17_14_port, ZN => n9027);
   U1691 : NAND4_X1 port map( A1 => n9030, A2 => n9029, A3 => n9028, A4 => 
                           n9027, ZN => n9036);
   U1692 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_14_port, B1 => 
                           n9384, B2 => REGISTERS_26_14_port, ZN => n9034);
   U1693 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_14_port, B1 => 
                           n9366, B2 => REGISTERS_16_14_port, ZN => n9033);
   U1694 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_14_port, B1 => 
                           n9380, B2 => REGISTERS_27_14_port, ZN => n9032);
   U1695 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_14_port, B1 => 
                           n9336, B2 => REGISTERS_18_14_port, ZN => n9031);
   U1696 : NAND4_X1 port map( A1 => n9034, A2 => n9033, A3 => n9032, A4 => 
                           n9031, ZN => n9035);
   U1697 : NOR2_X1 port map( A1 => n9036, A2 => n9035, ZN => n9048);
   U1698 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_5_14_port, B1 => 
                           n9407, B2 => REGISTERS_0_14_port, ZN => n9040);
   U1699 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_7_14_port, B1 => 
                           n9394, B2 => REGISTERS_1_14_port, ZN => n9039);
   U1700 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_14_port, B1 => 
                           n9322, B2 => REGISTERS_2_14_port, ZN => n9038);
   U1701 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_14_port, B1 => 
                           n9294, B2 => REGISTERS_3_14_port, ZN => n9037);
   U1702 : NAND4_X1 port map( A1 => n9040, A2 => n9039, A3 => n9038, A4 => 
                           n9037, ZN => n9046);
   U1703 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_14_port, B1 => 
                           n9322, B2 => REGISTERS_10_14_port, ZN => n9044);
   U1704 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_14_14_port, B1 => 
                           n9319, B2 => REGISTERS_13_14_port, ZN => n9043);
   U1705 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_14_port, B1 => 
                           n9294, B2 => REGISTERS_11_14_port, ZN => n9042);
   U1706 : AOI22_X1 port map( A1 => n9320, A2 => REGISTERS_9_14_port, B1 => 
                           n9392, B2 => REGISTERS_8_14_port, ZN => n9041);
   U1707 : NAND4_X1 port map( A1 => n9044, A2 => n9043, A3 => n9042, A4 => 
                           n9041, ZN => n9045);
   U1708 : AOI22_X1 port map( A1 => n9258, A2 => n9046, B1 => n9256, B2 => 
                           n9045, ZN => n9047);
   U1709 : OAI21_X1 port map( B1 => n9419, B2 => n9048, A => n9047, ZN => N431)
                           ;
   U1710 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_13_port, B1 => 
                           n9384, B2 => REGISTERS_26_13_port, ZN => n9052);
   U1711 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_13_port, B1 => 
                           n9372, B2 => REGISTERS_24_13_port, ZN => n9051);
   U1712 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_13_port, B1 => 
                           n9380, B2 => REGISTERS_27_13_port, ZN => n9050);
   U1713 : AOI22_X1 port map( A1 => n9382, A2 => REGISTERS_20_13_port, B1 => 
                           n9172, B2 => REGISTERS_17_13_port, ZN => n9049);
   U1714 : NAND4_X1 port map( A1 => n9052, A2 => n9051, A3 => n9050, A4 => 
                           n9049, ZN => n9058);
   U1715 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_13_port, B1 => 
                           n9077, B2 => REGISTERS_25_13_port, ZN => n9056);
   U1716 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_13_port, B1 => 
                           n9366, B2 => REGISTERS_16_13_port, ZN => n9055);
   U1717 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_13_port, B1 => 
                           n9381, B2 => REGISTERS_31_13_port, ZN => n9054);
   U1718 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_13_port, B1 => 
                           n9336, B2 => REGISTERS_18_13_port, ZN => n9053);
   U1719 : NAND4_X1 port map( A1 => n9056, A2 => n9055, A3 => n9054, A4 => 
                           n9053, ZN => n9057);
   U1720 : NOR2_X1 port map( A1 => n9058, A2 => n9057, ZN => n9070);
   U1721 : AOI22_X1 port map( A1 => n9403, A2 => REGISTERS_3_13_port, B1 => 
                           n9110, B2 => REGISTERS_2_13_port, ZN => n9062);
   U1722 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_13_port, B1 => 
                           n9320, B2 => REGISTERS_1_13_port, ZN => n9061);
   U1723 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_6_13_port, B1 => 
                           n9407, B2 => REGISTERS_0_13_port, ZN => n9060);
   U1724 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_5_13_port, B1 => 
                           n9408, B2 => REGISTERS_7_13_port, ZN => n9059);
   U1725 : NAND4_X1 port map( A1 => n9062, A2 => n9061, A3 => n9060, A4 => 
                           n9059, ZN => n9068);
   U1726 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_13_port, B1 => 
                           n9396, B2 => REGISTERS_11_13_port, ZN => n9066);
   U1727 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_13_port, B1 => 
                           n9401, B2 => REGISTERS_12_13_port, ZN => n9065);
   U1728 : AOI22_X1 port map( A1 => n9394, A2 => REGISTERS_9_13_port, B1 => 
                           n9327, B2 => REGISTERS_8_13_port, ZN => n9064);
   U1729 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_13_port, B1 => 
                           n9405, B2 => REGISTERS_10_13_port, ZN => n9063);
   U1730 : NAND4_X1 port map( A1 => n9066, A2 => n9065, A3 => n9064, A4 => 
                           n9063, ZN => n9067);
   U1731 : AOI22_X1 port map( A1 => n9258, A2 => n9068, B1 => n9256, B2 => 
                           n9067, ZN => n9069);
   U1732 : OAI21_X1 port map( B1 => n9365, B2 => n9070, A => n9069, ZN => N430)
                           ;
   U1733 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_12_port, B1 => 
                           n9343, B2 => REGISTERS_19_12_port, ZN => n9075);
   U1734 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_12_port, B1 => 
                           n9261, B2 => REGISTERS_23_12_port, ZN => n9074);
   U1735 : AOI22_X1 port map( A1 => n9071, A2 => REGISTERS_24_12_port, B1 => 
                           n9381, B2 => REGISTERS_31_12_port, ZN => n9073);
   U1736 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_12_port, B1 => 
                           n9172, B2 => REGISTERS_17_12_port, ZN => n9072);
   U1737 : NAND4_X1 port map( A1 => n9075, A2 => n9074, A3 => n9073, A4 => 
                           n9072, ZN => n9083);
   U1738 : AOI22_X1 port map( A1 => n9120, A2 => REGISTERS_26_12_port, B1 => 
                           n9336, B2 => REGISTERS_18_12_port, ZN => n9081);
   U1739 : AOI22_X1 port map( A1 => n9076, A2 => REGISTERS_16_12_port, B1 => 
                           n9380, B2 => REGISTERS_27_12_port, ZN => n9080);
   U1740 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_12_port, B1 => 
                           n9077, B2 => REGISTERS_25_12_port, ZN => n9079);
   U1741 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_12_port, B1 => 
                           n9368, B2 => REGISTERS_21_12_port, ZN => n9078);
   U1742 : NAND4_X1 port map( A1 => n9081, A2 => n9080, A3 => n9079, A4 => 
                           n9078, ZN => n9082);
   U1743 : NOR2_X1 port map( A1 => n9083, A2 => n9082, ZN => n9095);
   U1744 : AOI22_X1 port map( A1 => n9395, A2 => REGISTERS_7_12_port, B1 => 
                           n9322, B2 => REGISTERS_2_12_port, ZN => n9087);
   U1745 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_12_port, B1 => 
                           n9406, B2 => REGISTERS_1_12_port, ZN => n9086);
   U1746 : AOI22_X1 port map( A1 => n9294, A2 => REGISTERS_3_12_port, B1 => 
                           n9392, B2 => REGISTERS_0_12_port, ZN => n9085);
   U1747 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_12_port, B1 => 
                           n9319, B2 => REGISTERS_5_12_port, ZN => n9084);
   U1748 : NAND4_X1 port map( A1 => n9087, A2 => n9086, A3 => n9085, A4 => 
                           n9084, ZN => n9093);
   U1749 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_14_12_port, B1 => 
                           n9356, B2 => REGISTERS_13_12_port, ZN => n9091);
   U1750 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_12_port, B1 => 
                           n9322, B2 => REGISTERS_10_12_port, ZN => n9090);
   U1751 : AOI22_X1 port map( A1 => n9395, A2 => REGISTERS_15_12_port, B1 => 
                           n9320, B2 => REGISTERS_9_12_port, ZN => n9089);
   U1752 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_12_port, B1 => 
                           n9327, B2 => REGISTERS_8_12_port, ZN => n9088);
   U1753 : NAND4_X1 port map( A1 => n9091, A2 => n9090, A3 => n9089, A4 => 
                           n9088, ZN => n9092);
   U1754 : AOI22_X1 port map( A1 => n9258, A2 => n9093, B1 => n9256, B2 => 
                           n9092, ZN => n9094);
   U1755 : OAI21_X1 port map( B1 => n9419, B2 => n9095, A => n9094, ZN => N429)
                           ;
   U1756 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_11_port, B1 => 
                           n9371, B2 => REGISTERS_29_11_port, ZN => n9099);
   U1757 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_11_port, B1 => 
                           n9172, B2 => REGISTERS_17_11_port, ZN => n9098);
   U1758 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_11_port, B1 => 
                           n9366, B2 => REGISTERS_16_11_port, ZN => n9097);
   U1759 : AOI22_X1 port map( A1 => n9368, A2 => REGISTERS_21_11_port, B1 => 
                           n9336, B2 => REGISTERS_18_11_port, ZN => n9096);
   U1760 : NAND4_X1 port map( A1 => n9099, A2 => n9098, A3 => n9097, A4 => 
                           n9096, ZN => n9105);
   U1761 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_11_port, B1 => 
                           n9380, B2 => REGISTERS_27_11_port, ZN => n9103);
   U1762 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_11_port, B1 => 
                           n9381, B2 => REGISTERS_31_11_port, ZN => n9102);
   U1763 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_11_port, B1 => 
                           n9370, B2 => REGISTERS_23_11_port, ZN => n9101);
   U1764 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_11_port, B1 => 
                           n9384, B2 => REGISTERS_26_11_port, ZN => n9100);
   U1765 : NAND4_X1 port map( A1 => n9103, A2 => n9102, A3 => n9101, A4 => 
                           n9100, ZN => n9104);
   U1766 : NOR2_X1 port map( A1 => n9105, A2 => n9104, ZN => n9119);
   U1767 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_11_port, B1 => 
                           n9394, B2 => REGISTERS_1_11_port, ZN => n9109);
   U1768 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_5_11_port, B1 => 
                           n9322, B2 => REGISTERS_2_11_port, ZN => n9108);
   U1769 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_11_port, B1 => 
                           n9395, B2 => REGISTERS_7_11_port, ZN => n9107);
   U1770 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_11_port, B1 => 
                           n9407, B2 => REGISTERS_0_11_port, ZN => n9106);
   U1771 : NAND4_X1 port map( A1 => n9109, A2 => n9108, A3 => n9107, A4 => 
                           n9106, ZN => n9117);
   U1772 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_13_11_port, B1 => 
                           n9110, B2 => REGISTERS_10_11_port, ZN => n9115);
   U1773 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_12_11_port, B1 => 
                           n9327, B2 => REGISTERS_8_11_port, ZN => n9114);
   U1774 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_11_port, B1 => 
                           n9406, B2 => REGISTERS_9_11_port, ZN => n9113);
   U1775 : AOI22_X1 port map( A1 => n9111, A2 => REGISTERS_14_11_port, B1 => 
                           n9403, B2 => REGISTERS_11_11_port, ZN => n9112);
   U1776 : NAND4_X1 port map( A1 => n9115, A2 => n9114, A3 => n9113, A4 => 
                           n9112, ZN => n9116);
   U1777 : AOI22_X1 port map( A1 => n9258, A2 => n9117, B1 => n9256, B2 => 
                           n9116, ZN => n9118);
   U1778 : OAI21_X1 port map( B1 => n9419, B2 => n9119, A => n9118, ZN => N428)
                           ;
   U1779 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_10_port, B1 => 
                           n9372, B2 => REGISTERS_24_10_port, ZN => n9125);
   U1780 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_10_port, B1 => 
                           n9366, B2 => REGISTERS_16_10_port, ZN => n9124);
   U1781 : AOI22_X1 port map( A1 => n9120, A2 => REGISTERS_26_10_port, B1 => 
                           n9336, B2 => REGISTERS_18_10_port, ZN => n9123);
   U1782 : AOI22_X1 port map( A1 => n9121, A2 => REGISTERS_28_10_port, B1 => 
                           n9312, B2 => REGISTERS_22_10_port, ZN => n9122);
   U1783 : NAND4_X1 port map( A1 => n9125, A2 => n9124, A3 => n9123, A4 => 
                           n9122, ZN => n9131);
   U1784 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_10_port, B1 => 
                           n9371, B2 => REGISTERS_29_10_port, ZN => n9129);
   U1785 : AOI22_X1 port map( A1 => n9368, A2 => REGISTERS_21_10_port, B1 => 
                           n9172, B2 => REGISTERS_17_10_port, ZN => n9128);
   U1786 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_10_port, B1 => 
                           n9307, B2 => REGISTERS_31_10_port, ZN => n9127);
   U1787 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_10_port, B1 => 
                           n9380, B2 => REGISTERS_27_10_port, ZN => n9126);
   U1788 : NAND4_X1 port map( A1 => n9129, A2 => n9128, A3 => n9127, A4 => 
                           n9126, ZN => n9130);
   U1789 : NOR2_X1 port map( A1 => n9131, A2 => n9130, ZN => n9143);
   U1790 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_10_port, B1 => 
                           n9392, B2 => REGISTERS_0_10_port, ZN => n9135);
   U1791 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_7_10_port, B1 => 
                           n9406, B2 => REGISTERS_1_10_port, ZN => n9134);
   U1792 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_10_port, B1 => 
                           n9405, B2 => REGISTERS_2_10_port, ZN => n9133);
   U1793 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_6_10_port, B1 => 
                           n9401, B2 => REGISTERS_4_10_port, ZN => n9132);
   U1794 : NAND4_X1 port map( A1 => n9135, A2 => n9134, A3 => n9133, A4 => 
                           n9132, ZN => n9141);
   U1795 : AOI22_X1 port map( A1 => n9351, A2 => REGISTERS_15_10_port, B1 => 
                           n9320, B2 => REGISTERS_9_10_port, ZN => n9139);
   U1796 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_10_port, B1 => 
                           n9322, B2 => REGISTERS_10_10_port, ZN => n9138);
   U1797 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_14_10_port, B1 => 
                           n9392, B2 => REGISTERS_8_10_port, ZN => n9137);
   U1798 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_10_port, B1 => 
                           n9356, B2 => REGISTERS_13_10_port, ZN => n9136);
   U1799 : NAND4_X1 port map( A1 => n9139, A2 => n9138, A3 => n9137, A4 => 
                           n9136, ZN => n9140);
   U1800 : AOI22_X1 port map( A1 => n9258, A2 => n9141, B1 => n9256, B2 => 
                           n9140, ZN => n9142);
   U1801 : OAI21_X1 port map( B1 => n9419, B2 => n9143, A => n9142, ZN => N427)
                           ;
   U1802 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_9_port, B1 => 
                           n9373, B2 => REGISTERS_25_9_port, ZN => n9148);
   U1803 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_9_port, B1 => 
                           n9144, B2 => REGISTERS_27_9_port, ZN => n9147);
   U1804 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_9_port, B1 => 
                           n9336, B2 => REGISTERS_18_9_port, ZN => n9146);
   U1805 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_9_port, B1 => 
                           n9372, B2 => REGISTERS_24_9_port, ZN => n9145);
   U1806 : NAND4_X1 port map( A1 => n9148, A2 => n9147, A3 => n9146, A4 => 
                           n9145, ZN => n9154);
   U1807 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_9_port, B1 => 
                           n9172, B2 => REGISTERS_17_9_port, ZN => n9152);
   U1808 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_9_port, B1 => 
                           n9381, B2 => REGISTERS_31_9_port, ZN => n9151);
   U1809 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_9_port, B1 => 
                           n9366, B2 => REGISTERS_16_9_port, ZN => n9150);
   U1810 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_9_port, B1 => 
                           n9384, B2 => REGISTERS_26_9_port, ZN => n9149);
   U1811 : NAND4_X1 port map( A1 => n9152, A2 => n9151, A3 => n9150, A4 => 
                           n9149, ZN => n9153);
   U1812 : NOR2_X1 port map( A1 => n9154, A2 => n9153, ZN => n9166);
   U1813 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_9_port, B1 => 
                           n9395, B2 => REGISTERS_7_9_port, ZN => n9158);
   U1814 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_9_port, B1 => 
                           n9405, B2 => REGISTERS_2_9_port, ZN => n9157);
   U1815 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_6_9_port, B1 => 
                           n9201, B2 => REGISTERS_4_9_port, ZN => n9156);
   U1816 : AOI22_X1 port map( A1 => n9319, A2 => REGISTERS_5_9_port, B1 => 
                           n9407, B2 => REGISTERS_0_9_port, ZN => n9155);
   U1817 : NAND4_X1 port map( A1 => n9158, A2 => n9157, A3 => n9156, A4 => 
                           n9155, ZN => n9164);
   U1818 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_14_9_port, B1 => 
                           n9403, B2 => REGISTERS_11_9_port, ZN => n9162);
   U1819 : AOI22_X1 port map( A1 => n9394, A2 => REGISTERS_9_9_port, B1 => 
                           n9322, B2 => REGISTERS_10_9_port, ZN => n9161);
   U1820 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_9_port, B1 => 
                           n9327, B2 => REGISTERS_8_9_port, ZN => n9160);
   U1821 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_9_port, B1 => 
                           n9356, B2 => REGISTERS_13_9_port, ZN => n9159);
   U1822 : NAND4_X1 port map( A1 => n9162, A2 => n9161, A3 => n9160, A4 => 
                           n9159, ZN => n9163);
   U1823 : AOI22_X1 port map( A1 => n9258, A2 => n9164, B1 => n9256, B2 => 
                           n9163, ZN => n9165);
   U1824 : OAI21_X1 port map( B1 => n9365, B2 => n9166, A => n9165, ZN => N426)
                           ;
   U1825 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_8_port, B1 => 
                           n9384, B2 => REGISTERS_26_8_port, ZN => n9171);
   U1826 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_8_port, B1 => 
                           n9366, B2 => REGISTERS_16_8_port, ZN => n9170);
   U1827 : AOI22_X1 port map( A1 => n9167, A2 => REGISTERS_30_8_port, B1 => 
                           n9372, B2 => REGISTERS_24_8_port, ZN => n9169);
   U1828 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_8_port, B1 => 
                           n9380, B2 => REGISTERS_27_8_port, ZN => n9168);
   U1829 : NAND4_X1 port map( A1 => n9171, A2 => n9170, A3 => n9169, A4 => 
                           n9168, ZN => n9178);
   U1830 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_8_port, B1 => 
                           n9312, B2 => REGISTERS_22_8_port, ZN => n9176);
   U1831 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_8_port, B1 => 
                           n9370, B2 => REGISTERS_23_8_port, ZN => n9175);
   U1832 : AOI22_X1 port map( A1 => n9379, A2 => REGISTERS_18_8_port, B1 => 
                           n9172, B2 => REGISTERS_17_8_port, ZN => n9174);
   U1833 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_8_port, B1 => 
                           n9342, B2 => REGISTERS_29_8_port, ZN => n9173);
   U1834 : NAND4_X1 port map( A1 => n9176, A2 => n9175, A3 => n9174, A4 => 
                           n9173, ZN => n9177);
   U1835 : NOR2_X1 port map( A1 => n9178, A2 => n9177, ZN => n9190);
   U1836 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_8_port, B1 => 
                           n9392, B2 => REGISTERS_0_8_port, ZN => n9182);
   U1837 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_6_8_port, B1 => 
                           n9401, B2 => REGISTERS_4_8_port, ZN => n9181);
   U1838 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_8_port, B1 => 
                           n9405, B2 => REGISTERS_2_8_port, ZN => n9180);
   U1839 : AOI22_X1 port map( A1 => n9356, A2 => REGISTERS_5_8_port, B1 => 
                           n9408, B2 => REGISTERS_7_8_port, ZN => n9179);
   U1840 : NAND4_X1 port map( A1 => n9182, A2 => n9181, A3 => n9180, A4 => 
                           n9179, ZN => n9188);
   U1841 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_8_port, B1 => 
                           n9322, B2 => REGISTERS_10_8_port, ZN => n9186);
   U1842 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_14_8_port, B1 => 
                           n9401, B2 => REGISTERS_12_8_port, ZN => n9185);
   U1843 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_8_port, B1 => 
                           n9395, B2 => REGISTERS_15_8_port, ZN => n9184);
   U1844 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_9_8_port, B1 => 
                           n9327, B2 => REGISTERS_8_8_port, ZN => n9183);
   U1845 : NAND4_X1 port map( A1 => n9186, A2 => n9185, A3 => n9184, A4 => 
                           n9183, ZN => n9187);
   U1846 : AOI22_X1 port map( A1 => n9258, A2 => n9188, B1 => n9256, B2 => 
                           n9187, ZN => n9189);
   U1847 : OAI21_X1 port map( B1 => n9419, B2 => n9190, A => n9189, ZN => N425)
                           ;
   U1848 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_7_port, B1 => 
                           n9378, B2 => REGISTERS_17_7_port, ZN => n9194);
   U1849 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_7_port, B1 => 
                           n9336, B2 => REGISTERS_18_7_port, ZN => n9193);
   U1850 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_7_port, B1 => 
                           n9370, B2 => REGISTERS_23_7_port, ZN => n9192);
   U1851 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_7_port, B1 => 
                           n9343, B2 => REGISTERS_19_7_port, ZN => n9191);
   U1852 : NAND4_X1 port map( A1 => n9194, A2 => n9193, A3 => n9192, A4 => 
                           n9191, ZN => n9200);
   U1853 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_7_port, B1 => 
                           n9366, B2 => REGISTERS_16_7_port, ZN => n9198);
   U1854 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_7_port, B1 => 
                           n9372, B2 => REGISTERS_24_7_port, ZN => n9197);
   U1855 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_7_port, B1 => 
                           n9384, B2 => REGISTERS_26_7_port, ZN => n9196);
   U1856 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_7_port, B1 => 
                           n9380, B2 => REGISTERS_27_7_port, ZN => n9195);
   U1857 : NAND4_X1 port map( A1 => n9198, A2 => n9197, A3 => n9196, A4 => 
                           n9195, ZN => n9199);
   U1858 : NOR2_X1 port map( A1 => n9200, A2 => n9199, ZN => n9213);
   U1859 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_0_7_port, B1 => 
                           n9322, B2 => REGISTERS_2_7_port, ZN => n9205);
   U1860 : AOI22_X1 port map( A1 => n9201, A2 => REGISTERS_4_7_port, B1 => 
                           n9351, B2 => REGISTERS_7_7_port, ZN => n9204);
   U1861 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_7_port, B1 => 
                           n9320, B2 => REGISTERS_1_7_port, ZN => n9203);
   U1862 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_7_port, B1 => 
                           n9294, B2 => REGISTERS_3_7_port, ZN => n9202);
   U1863 : NAND4_X1 port map( A1 => n9205, A2 => n9204, A3 => n9203, A4 => 
                           n9202, ZN => n9211);
   U1864 : AOI22_X1 port map( A1 => n9401, A2 => REGISTERS_12_7_port, B1 => 
                           n9403, B2 => REGISTERS_11_7_port, ZN => n9209);
   U1865 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_7_port, B1 => 
                           n9394, B2 => REGISTERS_9_7_port, ZN => n9208);
   U1866 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_8_7_port, B1 => 
                           n9405, B2 => REGISTERS_10_7_port, ZN => n9207);
   U1867 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_7_port, B1 => 
                           n9395, B2 => REGISTERS_15_7_port, ZN => n9206);
   U1868 : NAND4_X1 port map( A1 => n9209, A2 => n9208, A3 => n9207, A4 => 
                           n9206, ZN => n9210);
   U1869 : AOI22_X1 port map( A1 => n9258, A2 => n9211, B1 => n9256, B2 => 
                           n9210, ZN => n9212);
   U1870 : OAI21_X1 port map( B1 => n9365, B2 => n9213, A => n9212, ZN => N424)
                           ;
   U1871 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_6_port, B1 => 
                           n9382, B2 => REGISTERS_20_6_port, ZN => n9217);
   U1872 : AOI22_X1 port map( A1 => n9366, A2 => REGISTERS_16_6_port, B1 => 
                           n9380, B2 => REGISTERS_27_6_port, ZN => n9216);
   U1873 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_6_port, B1 => 
                           n9370, B2 => REGISTERS_23_6_port, ZN => n9215);
   U1874 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_6_port, B1 => 
                           n9372, B2 => REGISTERS_24_6_port, ZN => n9214);
   U1875 : NAND4_X1 port map( A1 => n9217, A2 => n9216, A3 => n9215, A4 => 
                           n9214, ZN => n9223);
   U1876 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_6_port, B1 => 
                           n9384, B2 => REGISTERS_26_6_port, ZN => n9221);
   U1877 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_6_port, B1 => 
                           n9307, B2 => REGISTERS_31_6_port, ZN => n9220);
   U1878 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_6_port, B1 => 
                           n9378, B2 => REGISTERS_17_6_port, ZN => n9219);
   U1879 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_6_port, B1 => 
                           n9336, B2 => REGISTERS_18_6_port, ZN => n9218);
   U1880 : NAND4_X1 port map( A1 => n9221, A2 => n9220, A3 => n9219, A4 => 
                           n9218, ZN => n9222);
   U1881 : NOR2_X1 port map( A1 => n9223, A2 => n9222, ZN => n9236);
   U1882 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_7_6_port, B1 => 
                           n9406, B2 => REGISTERS_1_6_port, ZN => n9227);
   U1883 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_6_port, B1 => 
                           n9327, B2 => REGISTERS_0_6_port, ZN => n9226);
   U1884 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_6_port, B1 => 
                           n9294, B2 => REGISTERS_3_6_port, ZN => n9225);
   U1885 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_6_port, B1 => 
                           n9322, B2 => REGISTERS_2_6_port, ZN => n9224);
   U1886 : NAND4_X1 port map( A1 => n9227, A2 => n9226, A3 => n9225, A4 => 
                           n9224, ZN => n9233);
   U1887 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_6_port, B1 => 
                           n9408, B2 => REGISTERS_15_6_port, ZN => n9231);
   U1888 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_6_port, B1 => 
                           n9407, B2 => REGISTERS_8_6_port, ZN => n9230);
   U1889 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_6_port, B1 => 
                           n9394, B2 => REGISTERS_9_6_port, ZN => n9229);
   U1890 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_6_port, B1 => 
                           n9405, B2 => REGISTERS_10_6_port, ZN => n9228);
   U1891 : NAND4_X1 port map( A1 => n9231, A2 => n9230, A3 => n9229, A4 => 
                           n9228, ZN => n9232);
   U1892 : AOI22_X1 port map( A1 => n9234, A2 => n9233, B1 => n9256, B2 => 
                           n9232, ZN => n9235);
   U1893 : OAI21_X1 port map( B1 => n9419, B2 => n9236, A => n9235, ZN => N423)
                           ;
   U1894 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_5_port, B1 => 
                           n9380, B2 => REGISTERS_27_5_port, ZN => n9240);
   U1895 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_5_port, B1 => 
                           n9384, B2 => REGISTERS_26_5_port, ZN => n9239);
   U1896 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_5_port, B1 => 
                           n9378, B2 => REGISTERS_17_5_port, ZN => n9238);
   U1897 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_5_port, B1 => 
                           n9373, B2 => REGISTERS_25_5_port, ZN => n9237);
   U1898 : NAND4_X1 port map( A1 => n9240, A2 => n9239, A3 => n9238, A4 => 
                           n9237, ZN => n9246);
   U1899 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_5_port, B1 => 
                           n9343, B2 => REGISTERS_19_5_port, ZN => n9244);
   U1900 : AOI22_X1 port map( A1 => n9366, A2 => REGISTERS_16_5_port, B1 => 
                           n9336, B2 => REGISTERS_18_5_port, ZN => n9243);
   U1901 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_5_port, B1 => 
                           n9370, B2 => REGISTERS_23_5_port, ZN => n9242);
   U1902 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_5_port, B1 => 
                           n9372, B2 => REGISTERS_24_5_port, ZN => n9241);
   U1903 : NAND4_X1 port map( A1 => n9244, A2 => n9243, A3 => n9242, A4 => 
                           n9241, ZN => n9245);
   U1904 : NOR2_X1 port map( A1 => n9246, A2 => n9245, ZN => n9260);
   U1905 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_5_port, B1 => 
                           n9322, B2 => REGISTERS_2_5_port, ZN => n9250);
   U1906 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_5_port, B1 => 
                           n9407, B2 => REGISTERS_0_5_port, ZN => n9249);
   U1907 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_5_port, B1 => 
                           n9351, B2 => REGISTERS_7_5_port, ZN => n9248);
   U1908 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_5_port, B1 => 
                           n9294, B2 => REGISTERS_3_5_port, ZN => n9247);
   U1909 : NAND4_X1 port map( A1 => n9250, A2 => n9249, A3 => n9248, A4 => 
                           n9247, ZN => n9257);
   U1910 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_5_port, B1 => 
                           n9405, B2 => REGISTERS_10_5_port, ZN => n9254);
   U1911 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_5_port, B1 => 
                           n9394, B2 => REGISTERS_9_5_port, ZN => n9253);
   U1912 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_5_port, B1 => 
                           n9351, B2 => REGISTERS_15_5_port, ZN => n9252);
   U1913 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_5_port, B1 => 
                           n9407, B2 => REGISTERS_8_5_port, ZN => n9251);
   U1914 : NAND4_X1 port map( A1 => n9254, A2 => n9253, A3 => n9252, A4 => 
                           n9251, ZN => n9255);
   U1915 : AOI22_X1 port map( A1 => n9258, A2 => n9257, B1 => n9256, B2 => 
                           n9255, ZN => n9259);
   U1916 : OAI21_X1 port map( B1 => n9365, B2 => n9260, A => n9259, ZN => N422)
                           ;
   U1917 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_4_port, B1 => 
                           n9336, B2 => REGISTERS_18_4_port, ZN => n9265);
   U1918 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_4_port, B1 => 
                           n9366, B2 => REGISTERS_16_4_port, ZN => n9264);
   U1919 : AOI22_X1 port map( A1 => n9261, A2 => REGISTERS_23_4_port, B1 => 
                           n9378, B2 => REGISTERS_17_4_port, ZN => n9263);
   U1920 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_4_port, B1 => 
                           n9380, B2 => REGISTERS_27_4_port, ZN => n9262);
   U1921 : NAND4_X1 port map( A1 => n9265, A2 => n9264, A3 => n9263, A4 => 
                           n9262, ZN => n9271);
   U1922 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_4_port, B1 => 
                           n9307, B2 => REGISTERS_31_4_port, ZN => n9269);
   U1923 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_4_port, B1 => 
                           n9384, B2 => REGISTERS_26_4_port, ZN => n9268);
   U1924 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_4_port, B1 => 
                           n9342, B2 => REGISTERS_29_4_port, ZN => n9267);
   U1925 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_4_port, B1 => 
                           n9373, B2 => REGISTERS_25_4_port, ZN => n9266);
   U1926 : NAND4_X1 port map( A1 => n9269, A2 => n9268, A3 => n9267, A4 => 
                           n9266, ZN => n9270);
   U1927 : NOR2_X1 port map( A1 => n9271, A2 => n9270, ZN => n9283);
   U1928 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_4_port, B1 => 
                           n9392, B2 => REGISTERS_0_4_port, ZN => n9275);
   U1929 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_4_port, B1 => 
                           n9408, B2 => REGISTERS_7_4_port, ZN => n9274);
   U1930 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_4_port, B1 => 
                           n9322, B2 => REGISTERS_2_4_port, ZN => n9273);
   U1931 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_4_port, B1 => 
                           n9403, B2 => REGISTERS_3_4_port, ZN => n9272);
   U1932 : NAND4_X1 port map( A1 => n9275, A2 => n9274, A3 => n9273, A4 => 
                           n9272, ZN => n9281);
   U1933 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_4_port, B1 => 
                           n9351, B2 => REGISTERS_15_4_port, ZN => n9279);
   U1934 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_9_4_port, B1 => 
                           n9405, B2 => REGISTERS_10_4_port, ZN => n9278);
   U1935 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_4_port, B1 => 
                           n9392, B2 => REGISTERS_8_4_port, ZN => n9277);
   U1936 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_4_port, B1 => 
                           n9403, B2 => REGISTERS_11_4_port, ZN => n9276);
   U1937 : NAND4_X1 port map( A1 => n9279, A2 => n9278, A3 => n9277, A4 => 
                           n9276, ZN => n9280);
   U1938 : AOI22_X1 port map( A1 => n9416, A2 => n9281, B1 => n9414, B2 => 
                           n9280, ZN => n9282);
   U1939 : OAI21_X1 port map( B1 => n9419, B2 => n9283, A => n9282, ZN => N421)
                           ;
   U1940 : AOI22_X1 port map( A1 => n9384, A2 => REGISTERS_26_3_port, B1 => 
                           n9336, B2 => REGISTERS_18_3_port, ZN => n9287);
   U1941 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_3_port, B1 => 
                           n9370, B2 => REGISTERS_23_3_port, ZN => n9286);
   U1942 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_3_port, B1 => 
                           n9366, B2 => REGISTERS_16_3_port, ZN => n9285);
   U1943 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_3_port, B1 => 
                           n9373, B2 => REGISTERS_25_3_port, ZN => n9284);
   U1944 : NAND4_X1 port map( A1 => n9287, A2 => n9286, A3 => n9285, A4 => 
                           n9284, ZN => n9293);
   U1945 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_3_port, B1 => 
                           n9343, B2 => REGISTERS_19_3_port, ZN => n9291);
   U1946 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_3_port, B1 => 
                           n9378, B2 => REGISTERS_17_3_port, ZN => n9290);
   U1947 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_3_port, B1 => 
                           n9380, B2 => REGISTERS_27_3_port, ZN => n9289);
   U1948 : AOI22_X1 port map( A1 => n9372, A2 => REGISTERS_24_3_port, B1 => 
                           n9307, B2 => REGISTERS_31_3_port, ZN => n9288);
   U1949 : NAND4_X1 port map( A1 => n9291, A2 => n9290, A3 => n9289, A4 => 
                           n9288, ZN => n9292);
   U1950 : NOR2_X1 port map( A1 => n9293, A2 => n9292, ZN => n9306);
   U1951 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_3_port, B1 => 
                           n9406, B2 => REGISTERS_1_3_port, ZN => n9298);
   U1952 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_7_3_port, B1 => 
                           n9322, B2 => REGISTERS_2_3_port, ZN => n9297);
   U1953 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_3_port, B1 => 
                           n9327, B2 => REGISTERS_0_3_port, ZN => n9296);
   U1954 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_3_port, B1 => 
                           n9294, B2 => REGISTERS_3_3_port, ZN => n9295);
   U1955 : NAND4_X1 port map( A1 => n9298, A2 => n9297, A3 => n9296, A4 => 
                           n9295, ZN => n9304);
   U1956 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_3_port, B1 => 
                           n9356, B2 => REGISTERS_13_3_port, ZN => n9302);
   U1957 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_3_port, B1 => 
                           n9392, B2 => REGISTERS_8_3_port, ZN => n9301);
   U1958 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_3_port, B1 => 
                           n9320, B2 => REGISTERS_9_3_port, ZN => n9300);
   U1959 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_3_port, B1 => 
                           n9405, B2 => REGISTERS_10_3_port, ZN => n9299);
   U1960 : NAND4_X1 port map( A1 => n9302, A2 => n9301, A3 => n9300, A4 => 
                           n9299, ZN => n9303);
   U1961 : AOI22_X1 port map( A1 => n9416, A2 => n9304, B1 => n9414, B2 => 
                           n9303, ZN => n9305);
   U1962 : OAI21_X1 port map( B1 => n9365, B2 => n9306, A => n9305, ZN => N420)
                           ;
   U1963 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_2_port, B1 => 
                           n9382, B2 => REGISTERS_20_2_port, ZN => n9311);
   U1964 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_2_port, B1 => 
                           n9307, B2 => REGISTERS_31_2_port, ZN => n9310);
   U1965 : AOI22_X1 port map( A1 => n9366, A2 => REGISTERS_16_2_port, B1 => 
                           n9336, B2 => REGISTERS_18_2_port, ZN => n9309);
   U1966 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_2_port, B1 => 
                           n9384, B2 => REGISTERS_26_2_port, ZN => n9308);
   U1967 : NAND4_X1 port map( A1 => n9311, A2 => n9310, A3 => n9309, A4 => 
                           n9308, ZN => n9318);
   U1968 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_2_port, B1 => 
                           n9312, B2 => REGISTERS_22_2_port, ZN => n9316);
   U1969 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_2_port, B1 => 
                           n9378, B2 => REGISTERS_17_2_port, ZN => n9315);
   U1970 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_2_port, B1 => 
                           n9372, B2 => REGISTERS_24_2_port, ZN => n9314);
   U1971 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_2_port, B1 => 
                           n9380, B2 => REGISTERS_27_2_port, ZN => n9313);
   U1972 : NAND4_X1 port map( A1 => n9316, A2 => n9315, A3 => n9314, A4 => 
                           n9313, ZN => n9317);
   U1973 : NOR2_X1 port map( A1 => n9318, A2 => n9317, ZN => n9335);
   U1974 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_2_port, B1 => 
                           n9319, B2 => REGISTERS_5_2_port, ZN => n9326);
   U1975 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_2_port, B1 => 
                           n9320, B2 => REGISTERS_1_2_port, ZN => n9325);
   U1976 : AOI22_X1 port map( A1 => n9321, A2 => REGISTERS_6_2_port, B1 => 
                           n9408, B2 => REGISTERS_7_2_port, ZN => n9324);
   U1977 : AOI22_X1 port map( A1 => n9327, A2 => REGISTERS_0_2_port, B1 => 
                           n9322, B2 => REGISTERS_2_2_port, ZN => n9323);
   U1978 : NAND4_X1 port map( A1 => n9326, A2 => n9325, A3 => n9324, A4 => 
                           n9323, ZN => n9333);
   U1979 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_11_2_port, B1 => 
                           n9395, B2 => REGISTERS_15_2_port, ZN => n9331);
   U1980 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_2_port, B1 => 
                           n9327, B2 => REGISTERS_8_2_port, ZN => n9330);
   U1981 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_9_2_port, B1 => 
                           n9405, B2 => REGISTERS_10_2_port, ZN => n9329);
   U1982 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_2_port, B1 => 
                           n9356, B2 => REGISTERS_13_2_port, ZN => n9328);
   U1983 : NAND4_X1 port map( A1 => n9331, A2 => n9330, A3 => n9329, A4 => 
                           n9328, ZN => n9332);
   U1984 : AOI22_X1 port map( A1 => n9416, A2 => n9333, B1 => n9414, B2 => 
                           n9332, ZN => n9334);
   U1985 : OAI21_X1 port map( B1 => n9419, B2 => n9335, A => n9334, ZN => N419)
                           ;
   U1986 : AOI22_X1 port map( A1 => n9370, A2 => REGISTERS_23_1_port, B1 => 
                           n9372, B2 => REGISTERS_24_1_port, ZN => n9341);
   U1987 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_1_port, B1 => 
                           n9336, B2 => REGISTERS_18_1_port, ZN => n9340);
   U1988 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_1_port, B1 => 
                           n9378, B2 => REGISTERS_17_1_port, ZN => n9339);
   U1989 : AOI22_X1 port map( A1 => n9337, A2 => REGISTERS_20_1_port, B1 => 
                           n9384, B2 => REGISTERS_26_1_port, ZN => n9338);
   U1990 : NAND4_X1 port map( A1 => n9341, A2 => n9340, A3 => n9339, A4 => 
                           n9338, ZN => n9350);
   U1991 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_1_port, B1 => 
                           n9366, B2 => REGISTERS_16_1_port, ZN => n9348);
   U1992 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_1_port, B1 => 
                           n9342, B2 => REGISTERS_29_1_port, ZN => n9347);
   U1993 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_1_port, B1 => 
                           n9380, B2 => REGISTERS_27_1_port, ZN => n9346);
   U1994 : AOI22_X1 port map( A1 => n9344, A2 => REGISTERS_21_1_port, B1 => 
                           n9343, B2 => REGISTERS_19_1_port, ZN => n9345);
   U1995 : NAND4_X1 port map( A1 => n9348, A2 => n9347, A3 => n9346, A4 => 
                           n9345, ZN => n9349);
   U1996 : NOR2_X1 port map( A1 => n9350, A2 => n9349, ZN => n9364);
   U1997 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_1_1_port, B1 => 
                           n9407, B2 => REGISTERS_0_1_port, ZN => n9355);
   U1998 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_1_port, B1 => 
                           n9351, B2 => REGISTERS_7_1_port, ZN => n9354);
   U1999 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_6_1_port, B1 => 
                           n9403, B2 => REGISTERS_3_1_port, ZN => n9353);
   U2000 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_1_port, B1 => 
                           n9405, B2 => REGISTERS_2_1_port, ZN => n9352);
   U2001 : NAND4_X1 port map( A1 => n9355, A2 => n9354, A3 => n9353, A4 => 
                           n9352, ZN => n9362);
   U2002 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_1_port, B1 => 
                           n9403, B2 => REGISTERS_11_1_port, ZN => n9360);
   U2003 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_12_1_port, B1 => 
                           n9356, B2 => REGISTERS_13_1_port, ZN => n9359);
   U2004 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_9_1_port, B1 => 
                           n9407, B2 => REGISTERS_8_1_port, ZN => n9358);
   U2005 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_1_port, B1 => 
                           n9405, B2 => REGISTERS_10_1_port, ZN => n9357);
   U2006 : NAND4_X1 port map( A1 => n9360, A2 => n9359, A3 => n9358, A4 => 
                           n9357, ZN => n9361);
   U2007 : AOI22_X1 port map( A1 => n9416, A2 => n9362, B1 => n9414, B2 => 
                           n9361, ZN => n9363);
   U2008 : OAI21_X1 port map( B1 => n9365, B2 => n9364, A => n9363, ZN => N418)
                           ;
   U2009 : AOI22_X1 port map( A1 => n9367, A2 => REGISTERS_22_0_port, B1 => 
                           n9366, B2 => REGISTERS_16_0_port, ZN => n9377);
   U2010 : AOI22_X1 port map( A1 => n9369, A2 => REGISTERS_30_0_port, B1 => 
                           n9368, B2 => REGISTERS_21_0_port, ZN => n9376);
   U2011 : AOI22_X1 port map( A1 => n9371, A2 => REGISTERS_29_0_port, B1 => 
                           n9370, B2 => REGISTERS_23_0_port, ZN => n9375);
   U2012 : AOI22_X1 port map( A1 => n9373, A2 => REGISTERS_25_0_port, B1 => 
                           n9372, B2 => REGISTERS_24_0_port, ZN => n9374);
   U2013 : NAND4_X1 port map( A1 => n9377, A2 => n9376, A3 => n9375, A4 => 
                           n9374, ZN => n9391);
   U2014 : AOI22_X1 port map( A1 => n9379, A2 => REGISTERS_18_0_port, B1 => 
                           n9378, B2 => REGISTERS_17_0_port, ZN => n9389);
   U2015 : AOI22_X1 port map( A1 => n9381, A2 => REGISTERS_31_0_port, B1 => 
                           n9380, B2 => REGISTERS_27_0_port, ZN => n9388);
   U2016 : AOI22_X1 port map( A1 => n9383, A2 => REGISTERS_19_0_port, B1 => 
                           n9382, B2 => REGISTERS_20_0_port, ZN => n9387);
   U2017 : AOI22_X1 port map( A1 => n9385, A2 => REGISTERS_28_0_port, B1 => 
                           n9384, B2 => REGISTERS_26_0_port, ZN => n9386);
   U2018 : NAND4_X1 port map( A1 => n9389, A2 => n9388, A3 => n9387, A4 => 
                           n9386, ZN => n9390);
   U2019 : NOR2_X1 port map( A1 => n9391, A2 => n9390, ZN => n9418);
   U2020 : AOI22_X1 port map( A1 => n9393, A2 => REGISTERS_4_0_port, B1 => 
                           n9392, B2 => REGISTERS_0_0_port, ZN => n9400);
   U2021 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_5_0_port, B1 => 
                           n9394, B2 => REGISTERS_1_0_port, ZN => n9399);
   U2022 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_6_0_port, B1 => 
                           n9405, B2 => REGISTERS_2_0_port, ZN => n9398);
   U2023 : AOI22_X1 port map( A1 => n9396, A2 => REGISTERS_3_0_port, B1 => 
                           n9395, B2 => REGISTERS_7_0_port, ZN => n9397);
   U2024 : NAND4_X1 port map( A1 => n9400, A2 => n9399, A3 => n9398, A4 => 
                           n9397, ZN => n9415);
   U2025 : AOI22_X1 port map( A1 => n9402, A2 => REGISTERS_14_0_port, B1 => 
                           n9401, B2 => REGISTERS_12_0_port, ZN => n9412);
   U2026 : AOI22_X1 port map( A1 => n9404, A2 => REGISTERS_13_0_port, B1 => 
                           n9403, B2 => REGISTERS_11_0_port, ZN => n9411);
   U2027 : AOI22_X1 port map( A1 => n9406, A2 => REGISTERS_9_0_port, B1 => 
                           n9405, B2 => REGISTERS_10_0_port, ZN => n9410);
   U2028 : AOI22_X1 port map( A1 => n9408, A2 => REGISTERS_15_0_port, B1 => 
                           n9407, B2 => REGISTERS_8_0_port, ZN => n9409);
   U2029 : NAND4_X1 port map( A1 => n9412, A2 => n9411, A3 => n9410, A4 => 
                           n9409, ZN => n9413);
   U2030 : AOI22_X1 port map( A1 => n9416, A2 => n9415, B1 => n9414, B2 => 
                           n9413, ZN => n9417);
   U2031 : OAI21_X1 port map( B1 => n9419, B2 => n9418, A => n9417, ZN => N417)
                           ;
   U2032 : NAND3_X1 port map( A1 => n8451, A2 => ENABLE, A3 => RD1, ZN => 
                           n10201);
   U2033 : INV_X1 port map( A => ADD_RD1(3), ZN => n9448);
   U2034 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => n9448, ZN => n9428);
   U2035 : INV_X1 port map( A => ADD_RD1(1), ZN => n9420);
   U2036 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n9420, 
                           ZN => n9442);
   U2037 : NOR2_X1 port map( A1 => n9428, A2 => n9442, ZN => n9898);
   U2038 : CLKBUF_X1 port map( A => n9898, Z => n10161);
   U2039 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n9429);
   U2040 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), A3 => 
                           ADD_RD1(2), ZN => n9443);
   U2041 : NOR2_X1 port map( A1 => n9429, A2 => n9443, ZN => n10061);
   U2042 : AOI22_X1 port map( A1 => REGISTERS_21_31_port, A2 => n10161, B1 => 
                           REGISTERS_31_31_port, B2 => n10061, ZN => n9426);
   U2043 : INV_X1 port map( A => ADD_RD1(0), ZN => n9422);
   U2044 : NAND3_X1 port map( A1 => ADD_RD1(2), A2 => n9422, A3 => n9420, ZN =>
                           n9436);
   U2045 : NOR2_X1 port map( A1 => n9436, A2 => n9429, ZN => n10166);
   U2046 : CLKBUF_X1 port map( A => n10166, Z => n10121);
   U2047 : INV_X1 port map( A => ADD_RD1(2), ZN => n9421);
   U2048 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => n9422, A3 => n9421, ZN =>
                           n9440);
   U2049 : NOR2_X1 port map( A1 => n9428, A2 => n9440, ZN => n9835);
   U2050 : CLKBUF_X1 port map( A => n9835, Z => n10154);
   U2051 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n10121, B1 => 
                           REGISTERS_18_31_port, B2 => n10154, ZN => n9425);
   U2052 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n9427);
   U2053 : NAND2_X1 port map( A1 => n9427, A2 => n9422, ZN => n9441);
   U2054 : NOR2_X1 port map( A1 => n9429, A2 => n9441, ZN => n10066);
   U2055 : CLKBUF_X1 port map( A => n10066, Z => n10165);
   U2056 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => n9421, 
                           ZN => n9437);
   U2057 : NOR2_X1 port map( A1 => n9429, A2 => n9437, ZN => n10168);
   U2058 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n10165, B1 => 
                           REGISTERS_27_31_port, B2 => n10168, ZN => n9424);
   U2059 : NAND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n9422, 
                           ZN => n9439);
   U2060 : NOR2_X1 port map( A1 => n9428, A2 => n9439, ZN => n10163);
   U2061 : CLKBUF_X1 port map( A => n10163, Z => n10087);
   U2062 : NOR2_X1 port map( A1 => n9428, A2 => n9443, ZN => n9992);
   U2063 : CLKBUF_X1 port map( A => n9992, Z => n10167);
   U2064 : AOI22_X1 port map( A1 => REGISTERS_22_31_port, A2 => n10087, B1 => 
                           REGISTERS_23_31_port, B2 => n10167, ZN => n9423);
   U2065 : NAND4_X1 port map( A1 => n9426, A2 => n9425, A3 => n9424, A4 => 
                           n9423, ZN => n9435);
   U2066 : NOR2_X1 port map( A1 => n9429, A2 => n9439, ZN => n10116);
   U2067 : CLKBUF_X1 port map( A => n10116, Z => n10150);
   U2068 : NOR2_X1 port map( A1 => n9428, A2 => n9441, ZN => n10153);
   U2069 : AOI22_X1 port map( A1 => REGISTERS_30_31_port, A2 => n10150, B1 => 
                           REGISTERS_16_31_port, B2 => n10153, ZN => n9433);
   U2070 : NOR2_X1 port map( A1 => n9428, A2 => n9436, ZN => n10162);
   U2071 : CLKBUF_X1 port map( A => n10162, Z => n10067);
   U2072 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n9427, ZN => n9438);
   U2073 : NOR2_X1 port map( A1 => n9429, A2 => n9438, ZN => n10093);
   U2074 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n10067, B1 => 
                           REGISTERS_25_31_port, B2 => n10093, ZN => n9432);
   U2075 : NOR2_X1 port map( A1 => n9429, A2 => n9440, ZN => n10122);
   U2076 : CLKBUF_X1 port map( A => n10122, Z => n10152);
   U2077 : NOR2_X1 port map( A1 => n9428, A2 => n9438, ZN => n10156);
   U2078 : AOI22_X1 port map( A1 => REGISTERS_26_31_port, A2 => n10152, B1 => 
                           REGISTERS_17_31_port, B2 => n10156, ZN => n9431);
   U2079 : NOR2_X1 port map( A1 => n9428, A2 => n9437, ZN => n10012);
   U2080 : CLKBUF_X1 port map( A => n10012, Z => n10155);
   U2081 : NOR2_X1 port map( A1 => n9429, A2 => n9442, ZN => n9921);
   U2082 : CLKBUF_X1 port map( A => n9921, Z => n10149);
   U2083 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n10155, B1 => 
                           REGISTERS_29_31_port, B2 => n10149, ZN => n9430);
   U2084 : NAND4_X1 port map( A1 => n9433, A2 => n9432, A3 => n9431, A4 => 
                           n9430, ZN => n9434);
   U2085 : NOR2_X1 port map( A1 => n9435, A2 => n9434, ZN => n9456);
   U2086 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n10148, 
                           ZN => n10198);
   U2087 : CLKBUF_X1 port map( A => n10198, Z => n10009);
   U2088 : INV_X1 port map( A => n9436, ZN => n10188);
   U2089 : CLKBUF_X1 port map( A => n10188, Z => n10101);
   U2090 : INV_X1 port map( A => n9437, ZN => n10187);
   U2091 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n10101, B1 => 
                           REGISTERS_3_31_port, B2 => n10187, ZN => n9447);
   U2092 : INV_X1 port map( A => n9438, ZN => n10189);
   U2093 : CLKBUF_X1 port map( A => n10189, Z => n10130);
   U2094 : INV_X1 port map( A => n9439, ZN => n10078);
   U2095 : CLKBUF_X1 port map( A => n10078, Z => n10175);
   U2096 : AOI22_X1 port map( A1 => REGISTERS_1_31_port, A2 => n10130, B1 => 
                           REGISTERS_6_31_port, B2 => n10175, ZN => n9446);
   U2097 : INV_X1 port map( A => n9440, ZN => n10102);
   U2098 : CLKBUF_X1 port map( A => n10102, Z => n10184);
   U2099 : INV_X1 port map( A => n9441, ZN => n10052);
   U2100 : CLKBUF_X1 port map( A => n10052, Z => n10185);
   U2101 : AOI22_X1 port map( A1 => REGISTERS_2_31_port, A2 => n10184, B1 => 
                           REGISTERS_0_31_port, B2 => n10185, ZN => n9445);
   U2102 : INV_X1 port map( A => n9442, ZN => n10047);
   U2103 : INV_X1 port map( A => n9443, ZN => n10176);
   U2104 : AOI22_X1 port map( A1 => REGISTERS_5_31_port, A2 => n10047, B1 => 
                           REGISTERS_7_31_port, B2 => n10176, ZN => n9444);
   U2105 : NAND4_X1 port map( A1 => n9447, A2 => n9446, A3 => n9445, A4 => 
                           n9444, ZN => n9454);
   U2106 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => n9448, A3 => n10148, ZN =>
                           n10196);
   U2107 : CLKBUF_X1 port map( A => n10196, Z => n10032);
   U2108 : CLKBUF_X1 port map( A => n10047, Z => n10129);
   U2109 : AOI22_X1 port map( A1 => REGISTERS_14_31_port, A2 => n10078, B1 => 
                           REGISTERS_13_31_port, B2 => n10129, ZN => n9452);
   U2110 : CLKBUF_X1 port map( A => n10102, Z => n10136);
   U2111 : AOI22_X1 port map( A1 => REGISTERS_9_31_port, A2 => n10130, B1 => 
                           REGISTERS_10_31_port, B2 => n10136, ZN => n9451);
   U2112 : CLKBUF_X1 port map( A => n10187, Z => n10178);
   U2113 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n10101, B1 => 
                           REGISTERS_11_31_port, B2 => n10178, ZN => n9450);
   U2114 : CLKBUF_X1 port map( A => n10176, Z => n10131);
   U2115 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n10131, B1 => 
                           REGISTERS_8_31_port, B2 => n10185, ZN => n9449);
   U2116 : NAND4_X1 port map( A1 => n9452, A2 => n9451, A3 => n9450, A4 => 
                           n9449, ZN => n9453);
   U2117 : AOI22_X1 port map( A1 => n10009, A2 => n9454, B1 => n10032, B2 => 
                           n9453, ZN => n9455);
   U2118 : OAI21_X1 port map( B1 => n10148, B2 => n9456, A => n9455, ZN => N416
                           );
   U2119 : AOI22_X1 port map( A1 => REGISTERS_26_30_port, A2 => n10152, B1 => 
                           REGISTERS_25_30_port, B2 => n10093, ZN => n9460);
   U2120 : AOI22_X1 port map( A1 => REGISTERS_22_30_port, A2 => n10087, B1 => 
                           REGISTERS_17_30_port, B2 => n10156, ZN => n9459);
   U2121 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n10067, B1 => 
                           REGISTERS_16_30_port, B2 => n10153, ZN => n9458);
   U2122 : AOI22_X1 port map( A1 => REGISTERS_30_30_port, A2 => n10150, B1 => 
                           REGISTERS_18_30_port, B2 => n9835, ZN => n9457);
   U2123 : NAND4_X1 port map( A1 => n9460, A2 => n9459, A3 => n9458, A4 => 
                           n9457, ZN => n9466);
   U2124 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n10121, B1 => 
                           REGISTERS_24_30_port, B2 => n10165, ZN => n9464);
   U2125 : CLKBUF_X1 port map( A => n10168, Z => n10094);
   U2126 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n10094, B1 => 
                           REGISTERS_31_30_port, B2 => n10061, ZN => n9463);
   U2127 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n10149, B1 => 
                           REGISTERS_23_30_port, B2 => n9992, ZN => n9462);
   U2128 : AOI22_X1 port map( A1 => REGISTERS_19_30_port, A2 => n10155, B1 => 
                           REGISTERS_21_30_port, B2 => n10161, ZN => n9461);
   U2129 : NAND4_X1 port map( A1 => n9464, A2 => n9463, A3 => n9462, A4 => 
                           n9461, ZN => n9465);
   U2130 : NOR2_X1 port map( A1 => n9466, A2 => n9465, ZN => n9478);
   U2131 : AOI22_X1 port map( A1 => REGISTERS_1_30_port, A2 => n10130, B1 => 
                           REGISTERS_0_30_port, B2 => n10185, ZN => n9470);
   U2132 : AOI22_X1 port map( A1 => REGISTERS_5_30_port, A2 => n10047, B1 => 
                           REGISTERS_2_30_port, B2 => n10136, ZN => n9469);
   U2133 : CLKBUF_X1 port map( A => n10176, Z => n10183);
   U2134 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n10101, B1 => 
                           REGISTERS_7_30_port, B2 => n10183, ZN => n9468);
   U2135 : CLKBUF_X1 port map( A => n10187, Z => n10137);
   U2136 : AOI22_X1 port map( A1 => REGISTERS_3_30_port, A2 => n10137, B1 => 
                           REGISTERS_6_30_port, B2 => n10175, ZN => n9467);
   U2137 : NAND4_X1 port map( A1 => n9470, A2 => n9469, A3 => n9468, A4 => 
                           n9467, ZN => n9476);
   U2138 : AOI22_X1 port map( A1 => REGISTERS_9_30_port, A2 => n10130, B1 => 
                           REGISTERS_13_30_port, B2 => n10129, ZN => n9474);
   U2139 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n10101, B1 => 
                           REGISTERS_10_30_port, B2 => n10136, ZN => n9473);
   U2140 : AOI22_X1 port map( A1 => REGISTERS_14_30_port, A2 => n10078, B1 => 
                           REGISTERS_11_30_port, B2 => n10178, ZN => n9472);
   U2141 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n10052, B1 => 
                           REGISTERS_15_30_port, B2 => n10183, ZN => n9471);
   U2142 : NAND4_X1 port map( A1 => n9474, A2 => n9473, A3 => n9472, A4 => 
                           n9471, ZN => n9475);
   U2143 : AOI22_X1 port map( A1 => n10009, A2 => n9476, B1 => n10032, B2 => 
                           n9475, ZN => n9477);
   U2144 : OAI21_X1 port map( B1 => n10148, B2 => n9478, A => n9477, ZN => N415
                           );
   U2145 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n10094, B1 => 
                           REGISTERS_19_29_port, B2 => n10155, ZN => n9482);
   U2146 : CLKBUF_X1 port map( A => n10156, Z => n10088);
   U2147 : AOI22_X1 port map( A1 => REGISTERS_17_29_port, A2 => n10088, B1 => 
                           REGISTERS_31_29_port, B2 => n10061, ZN => n9481);
   U2148 : AOI22_X1 port map( A1 => REGISTERS_26_29_port, A2 => n10152, B1 => 
                           REGISTERS_28_29_port, B2 => n10121, ZN => n9480);
   U2149 : AOI22_X1 port map( A1 => REGISTERS_18_29_port, A2 => n10154, B1 => 
                           REGISTERS_30_29_port, B2 => n10116, ZN => n9479);
   U2150 : NAND4_X1 port map( A1 => n9482, A2 => n9481, A3 => n9480, A4 => 
                           n9479, ZN => n9488);
   U2151 : CLKBUF_X1 port map( A => n10153, Z => n10115);
   U2152 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n10115, B1 => 
                           REGISTERS_21_29_port, B2 => n9898, ZN => n9486);
   U2153 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n10167, B1 => 
                           REGISTERS_24_29_port, B2 => n10066, ZN => n9485);
   U2154 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n10067, B1 => 
                           REGISTERS_25_29_port, B2 => n10093, ZN => n9484);
   U2155 : AOI22_X1 port map( A1 => REGISTERS_22_29_port, A2 => n10087, B1 => 
                           REGISTERS_29_29_port, B2 => n9921, ZN => n9483);
   U2156 : NAND4_X1 port map( A1 => n9486, A2 => n9485, A3 => n9484, A4 => 
                           n9483, ZN => n9487);
   U2157 : NOR2_X1 port map( A1 => n9488, A2 => n9487, ZN => n9500);
   U2158 : CLKBUF_X1 port map( A => n10189, Z => n10138);
   U2159 : AOI22_X1 port map( A1 => REGISTERS_7_29_port, A2 => n10131, B1 => 
                           REGISTERS_1_29_port, B2 => n10138, ZN => n9492);
   U2160 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n10137, B1 => 
                           REGISTERS_5_29_port, B2 => n10129, ZN => n9491);
   U2161 : AOI22_X1 port map( A1 => REGISTERS_2_29_port, A2 => n10102, B1 => 
                           REGISTERS_6_29_port, B2 => n10175, ZN => n9490);
   U2162 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n10101, B1 => 
                           REGISTERS_0_29_port, B2 => n10052, ZN => n9489);
   U2163 : NAND4_X1 port map( A1 => n9492, A2 => n9491, A3 => n9490, A4 => 
                           n9489, ZN => n9498);
   U2164 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n10101, B1 => 
                           REGISTERS_8_29_port, B2 => n10185, ZN => n9496);
   U2165 : AOI22_X1 port map( A1 => REGISTERS_13_29_port, A2 => n10047, B1 => 
                           REGISTERS_11_29_port, B2 => n10178, ZN => n9495);
   U2166 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n10131, B1 => 
                           REGISTERS_10_29_port, B2 => n10102, ZN => n9494);
   U2167 : AOI22_X1 port map( A1 => REGISTERS_14_29_port, A2 => n10078, B1 => 
                           REGISTERS_9_29_port, B2 => n10138, ZN => n9493);
   U2168 : NAND4_X1 port map( A1 => n9496, A2 => n9495, A3 => n9494, A4 => 
                           n9493, ZN => n9497);
   U2169 : AOI22_X1 port map( A1 => n10009, A2 => n9498, B1 => n10032, B2 => 
                           n9497, ZN => n9499);
   U2170 : OAI21_X1 port map( B1 => n10148, B2 => n9500, A => n9499, ZN => N414
                           );
   U2171 : AOI22_X1 port map( A1 => REGISTERS_19_28_port, A2 => n10155, B1 => 
                           REGISTERS_30_28_port, B2 => n10116, ZN => n9504);
   U2172 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n10094, B1 => 
                           REGISTERS_22_28_port, B2 => n10087, ZN => n9503);
   U2173 : CLKBUF_X1 port map( A => n10061, Z => n10164);
   U2174 : AOI22_X1 port map( A1 => REGISTERS_31_28_port, A2 => n10164, B1 => 
                           REGISTERS_25_28_port, B2 => n10093, ZN => n9502);
   U2175 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n10149, B1 => 
                           REGISTERS_18_28_port, B2 => n9835, ZN => n9501);
   U2176 : NAND4_X1 port map( A1 => n9504, A2 => n9503, A3 => n9502, A4 => 
                           n9501, ZN => n9510);
   U2177 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n10115, B1 => 
                           REGISTERS_20_28_port, B2 => n10162, ZN => n9508);
   U2178 : AOI22_X1 port map( A1 => REGISTERS_26_28_port, A2 => n10152, B1 => 
                           REGISTERS_23_28_port, B2 => n9992, ZN => n9507);
   U2179 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n10165, B1 => 
                           REGISTERS_17_28_port, B2 => n10156, ZN => n9506);
   U2180 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n10121, B1 => 
                           REGISTERS_21_28_port, B2 => n9898, ZN => n9505);
   U2181 : NAND4_X1 port map( A1 => n9508, A2 => n9507, A3 => n9506, A4 => 
                           n9505, ZN => n9509);
   U2182 : NOR2_X1 port map( A1 => n9510, A2 => n9509, ZN => n9522);
   U2183 : AOI22_X1 port map( A1 => REGISTERS_1_28_port, A2 => n10130, B1 => 
                           REGISTERS_2_28_port, B2 => n10102, ZN => n9514);
   U2184 : AOI22_X1 port map( A1 => REGISTERS_5_28_port, A2 => n10047, B1 => 
                           REGISTERS_0_28_port, B2 => n10185, ZN => n9513);
   U2185 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n10101, B1 => 
                           REGISTERS_3_28_port, B2 => n10178, ZN => n9512);
   U2186 : CLKBUF_X1 port map( A => n10078, Z => n10186);
   U2187 : AOI22_X1 port map( A1 => REGISTERS_6_28_port, A2 => n10186, B1 => 
                           REGISTERS_7_28_port, B2 => n10183, ZN => n9511);
   U2188 : NAND4_X1 port map( A1 => n9514, A2 => n9513, A3 => n9512, A4 => 
                           n9511, ZN => n9520);
   U2189 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n10052, B1 => 
                           REGISTERS_14_28_port, B2 => n10078, ZN => n9518);
   U2190 : CLKBUF_X1 port map( A => n10047, Z => n10190);
   U2191 : AOI22_X1 port map( A1 => REGISTERS_13_28_port, A2 => n10190, B1 => 
                           REGISTERS_12_28_port, B2 => n10101, ZN => n9517);
   U2192 : AOI22_X1 port map( A1 => REGISTERS_9_28_port, A2 => n10130, B1 => 
                           REGISTERS_15_28_port, B2 => n10183, ZN => n9516);
   U2193 : AOI22_X1 port map( A1 => REGISTERS_10_28_port, A2 => n10102, B1 => 
                           REGISTERS_11_28_port, B2 => n10178, ZN => n9515);
   U2194 : NAND4_X1 port map( A1 => n9518, A2 => n9517, A3 => n9516, A4 => 
                           n9515, ZN => n9519);
   U2195 : AOI22_X1 port map( A1 => n10009, A2 => n9520, B1 => n10032, B2 => 
                           n9519, ZN => n9521);
   U2196 : OAI21_X1 port map( B1 => n10148, B2 => n9522, A => n9521, ZN => N413
                           );
   U2197 : AOI22_X1 port map( A1 => REGISTERS_17_27_port, A2 => n10088, B1 => 
                           REGISTERS_21_27_port, B2 => n9898, ZN => n9526);
   U2198 : AOI22_X1 port map( A1 => REGISTERS_22_27_port, A2 => n10087, B1 => 
                           REGISTERS_18_27_port, B2 => n9835, ZN => n9525);
   U2199 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n10165, B1 => 
                           REGISTERS_19_27_port, B2 => n10012, ZN => n9524);
   U2200 : AOI22_X1 port map( A1 => REGISTERS_31_27_port, A2 => n10164, B1 => 
                           REGISTERS_26_27_port, B2 => n10122, ZN => n9523);
   U2201 : NAND4_X1 port map( A1 => n9526, A2 => n9525, A3 => n9524, A4 => 
                           n9523, ZN => n9532);
   U2202 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n10121, B1 => 
                           REGISTERS_27_27_port, B2 => n10168, ZN => n9530);
   U2203 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n10067, B1 => 
                           REGISTERS_29_27_port, B2 => n9921, ZN => n9529);
   U2204 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n10115, B1 => 
                           REGISTERS_30_27_port, B2 => n10116, ZN => n9528);
   U2205 : AOI22_X1 port map( A1 => REGISTERS_23_27_port, A2 => n10167, B1 => 
                           REGISTERS_25_27_port, B2 => n10093, ZN => n9527);
   U2206 : NAND4_X1 port map( A1 => n9530, A2 => n9529, A3 => n9528, A4 => 
                           n9527, ZN => n9531);
   U2207 : NOR2_X1 port map( A1 => n9532, A2 => n9531, ZN => n9544);
   U2208 : AOI22_X1 port map( A1 => REGISTERS_5_27_port, A2 => n10047, B1 => 
                           REGISTERS_1_27_port, B2 => n10138, ZN => n9536);
   U2209 : CLKBUF_X1 port map( A => n10052, Z => n10177);
   U2210 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n10177, B1 => 
                           REGISTERS_3_27_port, B2 => n10187, ZN => n9535);
   U2211 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n10101, B1 => 
                           REGISTERS_6_27_port, B2 => n10078, ZN => n9534);
   U2212 : AOI22_X1 port map( A1 => REGISTERS_2_27_port, A2 => n10102, B1 => 
                           REGISTERS_7_27_port, B2 => n10183, ZN => n9533);
   U2213 : NAND4_X1 port map( A1 => n9536, A2 => n9535, A3 => n9534, A4 => 
                           n9533, ZN => n9542);
   U2214 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n10101, B1 => 
                           REGISTERS_10_27_port, B2 => n10136, ZN => n9540);
   U2215 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n10137, B1 => 
                           REGISTERS_13_27_port, B2 => n10129, ZN => n9539);
   U2216 : AOI22_X1 port map( A1 => REGISTERS_15_27_port, A2 => n10131, B1 => 
                           REGISTERS_8_27_port, B2 => n10185, ZN => n9538);
   U2217 : AOI22_X1 port map( A1 => REGISTERS_9_27_port, A2 => n10130, B1 => 
                           REGISTERS_14_27_port, B2 => n10175, ZN => n9537);
   U2218 : NAND4_X1 port map( A1 => n9540, A2 => n9539, A3 => n9538, A4 => 
                           n9537, ZN => n9541);
   U2219 : AOI22_X1 port map( A1 => n10009, A2 => n9542, B1 => n10032, B2 => 
                           n9541, ZN => n9543);
   U2220 : OAI21_X1 port map( B1 => n10148, B2 => n9544, A => n9543, ZN => N412
                           );
   U2221 : AOI22_X1 port map( A1 => REGISTERS_23_26_port, A2 => n10167, B1 => 
                           REGISTERS_28_26_port, B2 => n10166, ZN => n9548);
   U2222 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n10115, B1 => 
                           REGISTERS_18_26_port, B2 => n9835, ZN => n9547);
   U2223 : AOI22_X1 port map( A1 => REGISTERS_26_26_port, A2 => n10152, B1 => 
                           REGISTERS_31_26_port, B2 => n10061, ZN => n9546);
   U2224 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n10067, B1 => 
                           REGISTERS_29_26_port, B2 => n9921, ZN => n9545);
   U2225 : NAND4_X1 port map( A1 => n9548, A2 => n9547, A3 => n9546, A4 => 
                           n9545, ZN => n9554);
   U2226 : CLKBUF_X1 port map( A => n10093, Z => n10151);
   U2227 : AOI22_X1 port map( A1 => REGISTERS_17_26_port, A2 => n10088, B1 => 
                           REGISTERS_25_26_port, B2 => n10151, ZN => n9552);
   U2228 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n10155, B1 => 
                           REGISTERS_27_26_port, B2 => n10168, ZN => n9551);
   U2229 : AOI22_X1 port map( A1 => REGISTERS_30_26_port, A2 => n10150, B1 => 
                           REGISTERS_24_26_port, B2 => n10066, ZN => n9550);
   U2230 : AOI22_X1 port map( A1 => REGISTERS_22_26_port, A2 => n10087, B1 => 
                           REGISTERS_21_26_port, B2 => n9898, ZN => n9549);
   U2231 : NAND4_X1 port map( A1 => n9552, A2 => n9551, A3 => n9550, A4 => 
                           n9549, ZN => n9553);
   U2232 : NOR2_X1 port map( A1 => n9554, A2 => n9553, ZN => n9566);
   U2233 : AOI22_X1 port map( A1 => REGISTERS_6_26_port, A2 => n10186, B1 => 
                           REGISTERS_1_26_port, B2 => n10138, ZN => n9558);
   U2234 : AOI22_X1 port map( A1 => REGISTERS_5_26_port, A2 => n10190, B1 => 
                           REGISTERS_0_26_port, B2 => n10052, ZN => n9557);
   U2235 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n10137, B1 => 
                           REGISTERS_2_26_port, B2 => n10102, ZN => n9556);
   U2236 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n10101, B1 => 
                           REGISTERS_7_26_port, B2 => n10176, ZN => n9555);
   U2237 : NAND4_X1 port map( A1 => n9558, A2 => n9557, A3 => n9556, A4 => 
                           n9555, ZN => n9564);
   U2238 : AOI22_X1 port map( A1 => REGISTERS_10_26_port, A2 => n10184, B1 => 
                           REGISTERS_11_26_port, B2 => n10178, ZN => n9562);
   U2239 : AOI22_X1 port map( A1 => REGISTERS_9_26_port, A2 => n10130, B1 => 
                           REGISTERS_8_26_port, B2 => n10052, ZN => n9561);
   U2240 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n10101, B1 => 
                           REGISTERS_13_26_port, B2 => n10047, ZN => n9560);
   U2241 : AOI22_X1 port map( A1 => REGISTERS_14_26_port, A2 => n10186, B1 => 
                           REGISTERS_15_26_port, B2 => n10183, ZN => n9559);
   U2242 : NAND4_X1 port map( A1 => n9562, A2 => n9561, A3 => n9560, A4 => 
                           n9559, ZN => n9563);
   U2243 : AOI22_X1 port map( A1 => n10009, A2 => n9564, B1 => n10032, B2 => 
                           n9563, ZN => n9565);
   U2244 : OAI21_X1 port map( B1 => n10148, B2 => n9566, A => n9565, ZN => N411
                           );
   U2245 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n10165, B1 => 
                           REGISTERS_31_25_port, B2 => n10061, ZN => n9570);
   U2246 : AOI22_X1 port map( A1 => REGISTERS_21_25_port, A2 => n10161, B1 => 
                           REGISTERS_18_25_port, B2 => n9835, ZN => n9569);
   U2247 : AOI22_X1 port map( A1 => REGISTERS_25_25_port, A2 => n10093, B1 => 
                           REGISTERS_19_25_port, B2 => n10012, ZN => n9568);
   U2248 : AOI22_X1 port map( A1 => REGISTERS_17_25_port, A2 => n10088, B1 => 
                           REGISTERS_30_25_port, B2 => n10150, ZN => n9567);
   U2249 : NAND4_X1 port map( A1 => n9570, A2 => n9569, A3 => n9568, A4 => 
                           n9567, ZN => n9576);
   U2250 : AOI22_X1 port map( A1 => REGISTERS_22_25_port, A2 => n10087, B1 => 
                           REGISTERS_16_25_port, B2 => n10153, ZN => n9574);
   U2251 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n10067, B1 => 
                           REGISTERS_26_25_port, B2 => n10152, ZN => n9573);
   U2252 : AOI22_X1 port map( A1 => REGISTERS_27_25_port, A2 => n10094, B1 => 
                           REGISTERS_28_25_port, B2 => n10166, ZN => n9572);
   U2253 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n10149, B1 => 
                           REGISTERS_23_25_port, B2 => n9992, ZN => n9571);
   U2254 : NAND4_X1 port map( A1 => n9574, A2 => n9573, A3 => n9572, A4 => 
                           n9571, ZN => n9575);
   U2255 : NOR2_X1 port map( A1 => n9576, A2 => n9575, ZN => n9588);
   U2256 : AOI22_X1 port map( A1 => REGISTERS_1_25_port, A2 => n10130, B1 => 
                           REGISTERS_3_25_port, B2 => n10187, ZN => n9580);
   U2257 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n10101, B1 => 
                           REGISTERS_7_25_port, B2 => n10176, ZN => n9579);
   U2258 : AOI22_X1 port map( A1 => REGISTERS_2_25_port, A2 => n10184, B1 => 
                           REGISTERS_5_25_port, B2 => n10190, ZN => n9578);
   U2259 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n10177, B1 => 
                           REGISTERS_6_25_port, B2 => n10175, ZN => n9577);
   U2260 : NAND4_X1 port map( A1 => n9580, A2 => n9579, A3 => n9578, A4 => 
                           n9577, ZN => n9586);
   U2261 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n10052, B1 => 
                           REGISTERS_11_25_port, B2 => n10178, ZN => n9584);
   U2262 : AOI22_X1 port map( A1 => REGISTERS_9_25_port, A2 => n10130, B1 => 
                           REGISTERS_15_25_port, B2 => n10183, ZN => n9583);
   U2263 : CLKBUF_X1 port map( A => n10188, Z => n10139);
   U2264 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n10139, B1 => 
                           REGISTERS_10_25_port, B2 => n10102, ZN => n9582);
   U2265 : AOI22_X1 port map( A1 => REGISTERS_13_25_port, A2 => n10129, B1 => 
                           REGISTERS_14_25_port, B2 => n10078, ZN => n9581);
   U2266 : NAND4_X1 port map( A1 => n9584, A2 => n9583, A3 => n9582, A4 => 
                           n9581, ZN => n9585);
   U2267 : AOI22_X1 port map( A1 => n10009, A2 => n9586, B1 => n10032, B2 => 
                           n9585, ZN => n9587);
   U2268 : OAI21_X1 port map( B1 => n10148, B2 => n9588, A => n9587, ZN => N410
                           );
   U2269 : AOI22_X1 port map( A1 => REGISTERS_21_24_port, A2 => n10161, B1 => 
                           REGISTERS_19_24_port, B2 => n10012, ZN => n9592);
   U2270 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n10165, B1 => 
                           REGISTERS_18_24_port, B2 => n9835, ZN => n9591);
   U2271 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n10094, B1 => 
                           REGISTERS_28_24_port, B2 => n10166, ZN => n9590);
   U2272 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n10162, B1 => 
                           REGISTERS_17_24_port, B2 => n10088, ZN => n9589);
   U2273 : NAND4_X1 port map( A1 => n9592, A2 => n9591, A3 => n9590, A4 => 
                           n9589, ZN => n9598);
   U2274 : AOI22_X1 port map( A1 => REGISTERS_26_24_port, A2 => n10152, B1 => 
                           REGISTERS_25_24_port, B2 => n10151, ZN => n9596);
   U2275 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n10167, B1 => 
                           REGISTERS_30_24_port, B2 => n10150, ZN => n9595);
   U2276 : AOI22_X1 port map( A1 => REGISTERS_22_24_port, A2 => n10087, B1 => 
                           REGISTERS_29_24_port, B2 => n9921, ZN => n9594);
   U2277 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n10115, B1 => 
                           REGISTERS_31_24_port, B2 => n10164, ZN => n9593);
   U2278 : NAND4_X1 port map( A1 => n9596, A2 => n9595, A3 => n9594, A4 => 
                           n9593, ZN => n9597);
   U2279 : NOR2_X1 port map( A1 => n9598, A2 => n9597, ZN => n9610);
   U2280 : AOI22_X1 port map( A1 => REGISTERS_2_24_port, A2 => n10102, B1 => 
                           REGISTERS_6_24_port, B2 => n10078, ZN => n9602);
   U2281 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n10177, B1 => 
                           REGISTERS_1_24_port, B2 => n10138, ZN => n9601);
   U2282 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n10131, B1 => 
                           REGISTERS_5_24_port, B2 => n10129, ZN => n9600);
   U2283 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n10137, B1 => 
                           REGISTERS_4_24_port, B2 => n10139, ZN => n9599);
   U2284 : NAND4_X1 port map( A1 => n9602, A2 => n9601, A3 => n9600, A4 => 
                           n9599, ZN => n9608);
   U2285 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n10101, B1 => 
                           REGISTERS_11_24_port, B2 => n10187, ZN => n9606);
   U2286 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n10185, B1 => 
                           REGISTERS_9_24_port, B2 => n10138, ZN => n9605);
   U2287 : AOI22_X1 port map( A1 => REGISTERS_15_24_port, A2 => n10131, B1 => 
                           REGISTERS_10_24_port, B2 => n10136, ZN => n9604);
   U2288 : AOI22_X1 port map( A1 => REGISTERS_13_24_port, A2 => n10047, B1 => 
                           REGISTERS_14_24_port, B2 => n10186, ZN => n9603);
   U2289 : NAND4_X1 port map( A1 => n9606, A2 => n9605, A3 => n9604, A4 => 
                           n9603, ZN => n9607);
   U2290 : AOI22_X1 port map( A1 => n10009, A2 => n9608, B1 => n10032, B2 => 
                           n9607, ZN => n9609);
   U2291 : OAI21_X1 port map( B1 => n10148, B2 => n9610, A => n9609, ZN => N409
                           );
   U2292 : AOI22_X1 port map( A1 => REGISTERS_17_23_port, A2 => n10088, B1 => 
                           REGISTERS_28_23_port, B2 => n10166, ZN => n9614);
   U2293 : AOI22_X1 port map( A1 => REGISTERS_21_23_port, A2 => n10161, B1 => 
                           REGISTERS_23_23_port, B2 => n9992, ZN => n9613);
   U2294 : AOI22_X1 port map( A1 => REGISTERS_19_23_port, A2 => n10155, B1 => 
                           REGISTERS_20_23_port, B2 => n10067, ZN => n9612);
   U2295 : AOI22_X1 port map( A1 => REGISTERS_26_23_port, A2 => n10122, B1 => 
                           REGISTERS_29_23_port, B2 => n9921, ZN => n9611);
   U2296 : NAND4_X1 port map( A1 => n9614, A2 => n9613, A3 => n9612, A4 => 
                           n9611, ZN => n9620);
   U2297 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n10165, B1 => 
                           REGISTERS_18_23_port, B2 => n9835, ZN => n9618);
   U2298 : AOI22_X1 port map( A1 => REGISTERS_31_23_port, A2 => n10164, B1 => 
                           REGISTERS_27_23_port, B2 => n10094, ZN => n9617);
   U2299 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n10115, B1 => 
                           REGISTERS_25_23_port, B2 => n10151, ZN => n9616);
   U2300 : AOI22_X1 port map( A1 => REGISTERS_22_23_port, A2 => n10087, B1 => 
                           REGISTERS_30_23_port, B2 => n10150, ZN => n9615);
   U2301 : NAND4_X1 port map( A1 => n9618, A2 => n9617, A3 => n9616, A4 => 
                           n9615, ZN => n9619);
   U2302 : NOR2_X1 port map( A1 => n9620, A2 => n9619, ZN => n9632);
   U2303 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n10131, B1 => 
                           REGISTERS_2_23_port, B2 => n10102, ZN => n9624);
   U2304 : AOI22_X1 port map( A1 => REGISTERS_6_23_port, A2 => n10175, B1 => 
                           REGISTERS_1_23_port, B2 => n10189, ZN => n9623);
   U2305 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n10177, B1 => 
                           REGISTERS_3_23_port, B2 => n10178, ZN => n9622);
   U2306 : AOI22_X1 port map( A1 => REGISTERS_5_23_port, A2 => n10190, B1 => 
                           REGISTERS_4_23_port, B2 => n10139, ZN => n9621);
   U2307 : NAND4_X1 port map( A1 => n9624, A2 => n9623, A3 => n9622, A4 => 
                           n9621, ZN => n9630);
   U2308 : AOI22_X1 port map( A1 => REGISTERS_10_23_port, A2 => n10184, B1 => 
                           REGISTERS_9_23_port, B2 => n10138, ZN => n9628);
   U2309 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n10137, B1 => 
                           REGISTERS_14_23_port, B2 => n10078, ZN => n9627);
   U2310 : AOI22_X1 port map( A1 => REGISTERS_13_23_port, A2 => n10129, B1 => 
                           REGISTERS_12_23_port, B2 => n10139, ZN => n9626);
   U2311 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n10052, B1 => 
                           REGISTERS_15_23_port, B2 => n10176, ZN => n9625);
   U2312 : NAND4_X1 port map( A1 => n9628, A2 => n9627, A3 => n9626, A4 => 
                           n9625, ZN => n9629);
   U2313 : AOI22_X1 port map( A1 => n10009, A2 => n9630, B1 => n10032, B2 => 
                           n9629, ZN => n9631);
   U2314 : OAI21_X1 port map( B1 => n10201, B2 => n9632, A => n9631, ZN => N408
                           );
   U2315 : AOI22_X1 port map( A1 => REGISTERS_17_22_port, A2 => n10088, B1 => 
                           REGISTERS_21_22_port, B2 => n9898, ZN => n9636);
   U2316 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n10115, B1 => 
                           REGISTERS_25_22_port, B2 => n10151, ZN => n9635);
   U2317 : AOI22_X1 port map( A1 => REGISTERS_30_22_port, A2 => n10150, B1 => 
                           REGISTERS_29_22_port, B2 => n9921, ZN => n9634);
   U2318 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n10155, B1 => 
                           REGISTERS_26_22_port, B2 => n10152, ZN => n9633);
   U2319 : NAND4_X1 port map( A1 => n9636, A2 => n9635, A3 => n9634, A4 => 
                           n9633, ZN => n9642);
   U2320 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n10121, B1 => 
                           REGISTERS_20_22_port, B2 => n10162, ZN => n9640);
   U2321 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n10165, B1 => 
                           REGISTERS_22_22_port, B2 => n10163, ZN => n9639);
   U2322 : AOI22_X1 port map( A1 => REGISTERS_31_22_port, A2 => n10164, B1 => 
                           REGISTERS_18_22_port, B2 => n9835, ZN => n9638);
   U2323 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n10167, B1 => 
                           REGISTERS_27_22_port, B2 => n10168, ZN => n9637);
   U2324 : NAND4_X1 port map( A1 => n9640, A2 => n9639, A3 => n9638, A4 => 
                           n9637, ZN => n9641);
   U2325 : NOR2_X1 port map( A1 => n9642, A2 => n9641, ZN => n9654);
   U2326 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n10137, B1 => 
                           REGISTERS_1_22_port, B2 => n10189, ZN => n9646);
   U2327 : AOI22_X1 port map( A1 => REGISTERS_6_22_port, A2 => n10078, B1 => 
                           REGISTERS_2_22_port, B2 => n10136, ZN => n9645);
   U2328 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n10176, B1 => 
                           REGISTERS_5_22_port, B2 => n10047, ZN => n9644);
   U2329 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n10185, B1 => 
                           REGISTERS_4_22_port, B2 => n10139, ZN => n9643);
   U2330 : NAND4_X1 port map( A1 => n9646, A2 => n9645, A3 => n9644, A4 => 
                           n9643, ZN => n9652);
   U2331 : AOI22_X1 port map( A1 => REGISTERS_14_22_port, A2 => n10186, B1 => 
                           REGISTERS_13_22_port, B2 => n10047, ZN => n9650);
   U2332 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n10131, B1 => 
                           REGISTERS_9_22_port, B2 => n10138, ZN => n9649);
   U2333 : AOI22_X1 port map( A1 => REGISTERS_10_22_port, A2 => n10136, B1 => 
                           REGISTERS_8_22_port, B2 => n10177, ZN => n9648);
   U2334 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n10101, B1 => 
                           REGISTERS_11_22_port, B2 => n10187, ZN => n9647);
   U2335 : NAND4_X1 port map( A1 => n9650, A2 => n9649, A3 => n9648, A4 => 
                           n9647, ZN => n9651);
   U2336 : AOI22_X1 port map( A1 => n10009, A2 => n9652, B1 => n10032, B2 => 
                           n9651, ZN => n9653);
   U2337 : OAI21_X1 port map( B1 => n10201, B2 => n9654, A => n9653, ZN => N407
                           );
   U2338 : AOI22_X1 port map( A1 => REGISTERS_30_21_port, A2 => n10150, B1 => 
                           REGISTERS_18_21_port, B2 => n10154, ZN => n9658);
   U2339 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n10162, B1 => 
                           REGISTERS_25_21_port, B2 => n10151, ZN => n9657);
   U2340 : AOI22_X1 port map( A1 => REGISTERS_22_21_port, A2 => n10163, B1 => 
                           REGISTERS_23_21_port, B2 => n9992, ZN => n9656);
   U2341 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n10115, B1 => 
                           REGISTERS_29_21_port, B2 => n9921, ZN => n9655);
   U2342 : NAND4_X1 port map( A1 => n9658, A2 => n9657, A3 => n9656, A4 => 
                           n9655, ZN => n9664);
   U2343 : AOI22_X1 port map( A1 => REGISTERS_26_21_port, A2 => n10152, B1 => 
                           REGISTERS_21_21_port, B2 => n9898, ZN => n9662);
   U2344 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n10012, B1 => 
                           REGISTERS_17_21_port, B2 => n10088, ZN => n9661);
   U2345 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n10165, B1 => 
                           REGISTERS_27_21_port, B2 => n10094, ZN => n9660);
   U2346 : AOI22_X1 port map( A1 => REGISTERS_31_21_port, A2 => n10164, B1 => 
                           REGISTERS_28_21_port, B2 => n10166, ZN => n9659);
   U2347 : NAND4_X1 port map( A1 => n9662, A2 => n9661, A3 => n9660, A4 => 
                           n9659, ZN => n9663);
   U2348 : NOR2_X1 port map( A1 => n9664, A2 => n9663, ZN => n9676);
   U2349 : AOI22_X1 port map( A1 => REGISTERS_5_21_port, A2 => n10129, B1 => 
                           REGISTERS_7_21_port, B2 => n10183, ZN => n9668);
   U2350 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n10185, B1 => 
                           REGISTERS_2_21_port, B2 => n10136, ZN => n9667);
   U2351 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n10139, B1 => 
                           REGISTERS_3_21_port, B2 => n10178, ZN => n9666);
   U2352 : AOI22_X1 port map( A1 => REGISTERS_6_21_port, A2 => n10078, B1 => 
                           REGISTERS_1_21_port, B2 => n10189, ZN => n9665);
   U2353 : NAND4_X1 port map( A1 => n9668, A2 => n9667, A3 => n9666, A4 => 
                           n9665, ZN => n9674);
   U2354 : AOI22_X1 port map( A1 => REGISTERS_14_21_port, A2 => n10175, B1 => 
                           REGISTERS_10_21_port, B2 => n10184, ZN => n9672);
   U2355 : AOI22_X1 port map( A1 => REGISTERS_15_21_port, A2 => n10183, B1 => 
                           REGISTERS_9_21_port, B2 => n10138, ZN => n9671);
   U2356 : AOI22_X1 port map( A1 => REGISTERS_13_21_port, A2 => n10190, B1 => 
                           REGISTERS_8_21_port, B2 => n10052, ZN => n9670);
   U2357 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n10188, B1 => 
                           REGISTERS_11_21_port, B2 => n10187, ZN => n9669);
   U2358 : NAND4_X1 port map( A1 => n9672, A2 => n9671, A3 => n9670, A4 => 
                           n9669, ZN => n9673);
   U2359 : AOI22_X1 port map( A1 => n10009, A2 => n9674, B1 => n10032, B2 => 
                           n9673, ZN => n9675);
   U2360 : OAI21_X1 port map( B1 => n10201, B2 => n9676, A => n9675, ZN => N406
                           );
   U2361 : AOI22_X1 port map( A1 => REGISTERS_30_20_port, A2 => n10116, B1 => 
                           REGISTERS_31_20_port, B2 => n10164, ZN => n9680);
   U2362 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n10115, B1 => 
                           REGISTERS_21_20_port, B2 => n9898, ZN => n9679);
   U2363 : AOI22_X1 port map( A1 => REGISTERS_18_20_port, A2 => n9835, B1 => 
                           REGISTERS_28_20_port, B2 => n10166, ZN => n9678);
   U2364 : AOI22_X1 port map( A1 => REGISTERS_25_20_port, A2 => n10093, B1 => 
                           REGISTERS_19_20_port, B2 => n10012, ZN => n9677);
   U2365 : NAND4_X1 port map( A1 => n9680, A2 => n9679, A3 => n9678, A4 => 
                           n9677, ZN => n9686);
   U2366 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n10094, B1 => 
                           REGISTERS_20_20_port, B2 => n10067, ZN => n9684);
   U2367 : AOI22_X1 port map( A1 => REGISTERS_23_20_port, A2 => n10167, B1 => 
                           REGISTERS_26_20_port, B2 => n10122, ZN => n9683);
   U2368 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n10149, B1 => 
                           REGISTERS_24_20_port, B2 => n10066, ZN => n9682);
   U2369 : AOI22_X1 port map( A1 => REGISTERS_17_20_port, A2 => n10088, B1 => 
                           REGISTERS_22_20_port, B2 => n10163, ZN => n9681);
   U2370 : NAND4_X1 port map( A1 => n9684, A2 => n9683, A3 => n9682, A4 => 
                           n9681, ZN => n9685);
   U2371 : NOR2_X1 port map( A1 => n9686, A2 => n9685, ZN => n9698);
   U2372 : AOI22_X1 port map( A1 => REGISTERS_5_20_port, A2 => n10129, B1 => 
                           REGISTERS_6_20_port, B2 => n10175, ZN => n9690);
   U2373 : AOI22_X1 port map( A1 => REGISTERS_2_20_port, A2 => n10136, B1 => 
                           REGISTERS_4_20_port, B2 => n10139, ZN => n9689);
   U2374 : AOI22_X1 port map( A1 => REGISTERS_1_20_port, A2 => n10189, B1 => 
                           REGISTERS_3_20_port, B2 => n10178, ZN => n9688);
   U2375 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n10183, B1 => 
                           REGISTERS_0_20_port, B2 => n10185, ZN => n9687);
   U2376 : NAND4_X1 port map( A1 => n9690, A2 => n9689, A3 => n9688, A4 => 
                           n9687, ZN => n9696);
   U2377 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n10052, B1 => 
                           REGISTERS_12_20_port, B2 => n10188, ZN => n9694);
   U2378 : AOI22_X1 port map( A1 => REGISTERS_9_20_port, A2 => n10130, B1 => 
                           REGISTERS_14_20_port, B2 => n10186, ZN => n9693);
   U2379 : AOI22_X1 port map( A1 => REGISTERS_13_20_port, A2 => n10190, B1 => 
                           REGISTERS_11_20_port, B2 => n10187, ZN => n9692);
   U2380 : AOI22_X1 port map( A1 => REGISTERS_10_20_port, A2 => n10102, B1 => 
                           REGISTERS_15_20_port, B2 => n10176, ZN => n9691);
   U2381 : NAND4_X1 port map( A1 => n9694, A2 => n9693, A3 => n9692, A4 => 
                           n9691, ZN => n9695);
   U2382 : AOI22_X1 port map( A1 => n10009, A2 => n9696, B1 => n10196, B2 => 
                           n9695, ZN => n9697);
   U2383 : OAI21_X1 port map( B1 => n10201, B2 => n9698, A => n9697, ZN => N405
                           );
   U2384 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n10121, B1 => 
                           REGISTERS_27_19_port, B2 => n10094, ZN => n9702);
   U2385 : AOI22_X1 port map( A1 => REGISTERS_19_19_port, A2 => n10155, B1 => 
                           REGISTERS_23_19_port, B2 => n9992, ZN => n9701);
   U2386 : AOI22_X1 port map( A1 => REGISTERS_17_19_port, A2 => n10156, B1 => 
                           REGISTERS_29_19_port, B2 => n9921, ZN => n9700);
   U2387 : AOI22_X1 port map( A1 => REGISTERS_26_19_port, A2 => n10122, B1 => 
                           REGISTERS_20_19_port, B2 => n10067, ZN => n9699);
   U2388 : NAND4_X1 port map( A1 => n9702, A2 => n9701, A3 => n9700, A4 => 
                           n9699, ZN => n9708);
   U2389 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n10153, B1 => 
                           REGISTERS_22_19_port, B2 => n10163, ZN => n9706);
   U2390 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n10066, B1 => 
                           REGISTERS_31_19_port, B2 => n10164, ZN => n9705);
   U2391 : AOI22_X1 port map( A1 => REGISTERS_30_19_port, A2 => n10116, B1 => 
                           REGISTERS_18_19_port, B2 => n10154, ZN => n9704);
   U2392 : AOI22_X1 port map( A1 => REGISTERS_25_19_port, A2 => n10151, B1 => 
                           REGISTERS_21_19_port, B2 => n9898, ZN => n9703);
   U2393 : NAND4_X1 port map( A1 => n9706, A2 => n9705, A3 => n9704, A4 => 
                           n9703, ZN => n9707);
   U2394 : NOR2_X1 port map( A1 => n9708, A2 => n9707, ZN => n9720);
   U2395 : CLKBUF_X1 port map( A => n10198, Z => n10034);
   U2396 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n10131, B1 => 
                           REGISTERS_3_19_port, B2 => n10187, ZN => n9712);
   U2397 : AOI22_X1 port map( A1 => REGISTERS_6_19_port, A2 => n10186, B1 => 
                           REGISTERS_4_19_port, B2 => n10139, ZN => n9711);
   U2398 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n10185, B1 => 
                           REGISTERS_2_19_port, B2 => n10136, ZN => n9710);
   U2399 : AOI22_X1 port map( A1 => REGISTERS_5_19_port, A2 => n10047, B1 => 
                           REGISTERS_1_19_port, B2 => n10189, ZN => n9709);
   U2400 : NAND4_X1 port map( A1 => n9712, A2 => n9711, A3 => n9710, A4 => 
                           n9709, ZN => n9718);
   U2401 : AOI22_X1 port map( A1 => REGISTERS_9_19_port, A2 => n10189, B1 => 
                           REGISTERS_10_19_port, B2 => n10102, ZN => n9716);
   U2402 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n10101, B1 => 
                           REGISTERS_8_19_port, B2 => n10052, ZN => n9715);
   U2403 : AOI22_X1 port map( A1 => REGISTERS_13_19_port, A2 => n10129, B1 => 
                           REGISTERS_14_19_port, B2 => n10186, ZN => n9714);
   U2404 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n10131, B1 => 
                           REGISTERS_11_19_port, B2 => n10178, ZN => n9713);
   U2405 : NAND4_X1 port map( A1 => n9716, A2 => n9715, A3 => n9714, A4 => 
                           n9713, ZN => n9717);
   U2406 : AOI22_X1 port map( A1 => n10034, A2 => n9718, B1 => n10032, B2 => 
                           n9717, ZN => n9719);
   U2407 : OAI21_X1 port map( B1 => n10201, B2 => n9720, A => n9719, ZN => N404
                           );
   U2408 : AOI22_X1 port map( A1 => REGISTERS_25_18_port, A2 => n10151, B1 => 
                           REGISTERS_28_18_port, B2 => n10166, ZN => n9724);
   U2409 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n10167, B1 => 
                           REGISTERS_30_18_port, B2 => n10150, ZN => n9723);
   U2410 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n10153, B1 => 
                           REGISTERS_31_18_port, B2 => n10164, ZN => n9722);
   U2411 : AOI22_X1 port map( A1 => REGISTERS_22_18_port, A2 => n10087, B1 => 
                           REGISTERS_29_18_port, B2 => n10149, ZN => n9721);
   U2412 : NAND4_X1 port map( A1 => n9724, A2 => n9723, A3 => n9722, A4 => 
                           n9721, ZN => n9730);
   U2413 : AOI22_X1 port map( A1 => REGISTERS_26_18_port, A2 => n10152, B1 => 
                           REGISTERS_27_18_port, B2 => n10168, ZN => n9728);
   U2414 : AOI22_X1 port map( A1 => REGISTERS_21_18_port, A2 => n9898, B1 => 
                           REGISTERS_18_18_port, B2 => n10154, ZN => n9727);
   U2415 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n10067, B1 => 
                           REGISTERS_19_18_port, B2 => n10012, ZN => n9726);
   U2416 : AOI22_X1 port map( A1 => REGISTERS_17_18_port, A2 => n10156, B1 => 
                           REGISTERS_24_18_port, B2 => n10066, ZN => n9725);
   U2417 : NAND4_X1 port map( A1 => n9728, A2 => n9727, A3 => n9726, A4 => 
                           n9725, ZN => n9729);
   U2418 : NOR2_X1 port map( A1 => n9730, A2 => n9729, ZN => n9742);
   U2419 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n10176, B1 => 
                           REGISTERS_2_18_port, B2 => n10136, ZN => n9734);
   U2420 : AOI22_X1 port map( A1 => REGISTERS_3_18_port, A2 => n10187, B1 => 
                           REGISTERS_0_18_port, B2 => n10185, ZN => n9733);
   U2421 : AOI22_X1 port map( A1 => REGISTERS_5_18_port, A2 => n10190, B1 => 
                           REGISTERS_4_18_port, B2 => n10188, ZN => n9732);
   U2422 : AOI22_X1 port map( A1 => REGISTERS_1_18_port, A2 => n10130, B1 => 
                           REGISTERS_6_18_port, B2 => n10186, ZN => n9731);
   U2423 : NAND4_X1 port map( A1 => n9734, A2 => n9733, A3 => n9732, A4 => 
                           n9731, ZN => n9740);
   U2424 : AOI22_X1 port map( A1 => REGISTERS_14_18_port, A2 => n10078, B1 => 
                           REGISTERS_10_18_port, B2 => n10136, ZN => n9738);
   U2425 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n10139, B1 => 
                           REGISTERS_11_18_port, B2 => n10187, ZN => n9737);
   U2426 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n10177, B1 => 
                           REGISTERS_13_18_port, B2 => n10190, ZN => n9736);
   U2427 : AOI22_X1 port map( A1 => REGISTERS_9_18_port, A2 => n10138, B1 => 
                           REGISTERS_15_18_port, B2 => n10183, ZN => n9735);
   U2428 : NAND4_X1 port map( A1 => n9738, A2 => n9737, A3 => n9736, A4 => 
                           n9735, ZN => n9739);
   U2429 : AOI22_X1 port map( A1 => n10034, A2 => n9740, B1 => n10032, B2 => 
                           n9739, ZN => n9741);
   U2430 : OAI21_X1 port map( B1 => n10201, B2 => n9742, A => n9741, ZN => N403
                           );
   U2431 : AOI22_X1 port map( A1 => REGISTERS_21_17_port, A2 => n9898, B1 => 
                           REGISTERS_22_17_port, B2 => n10163, ZN => n9746);
   U2432 : AOI22_X1 port map( A1 => REGISTERS_30_17_port, A2 => n10150, B1 => 
                           REGISTERS_19_17_port, B2 => n10012, ZN => n9745);
   U2433 : AOI22_X1 port map( A1 => REGISTERS_31_17_port, A2 => n10061, B1 => 
                           REGISTERS_27_17_port, B2 => n10094, ZN => n9744);
   U2434 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n10067, B1 => 
                           REGISTERS_29_17_port, B2 => n10149, ZN => n9743);
   U2435 : NAND4_X1 port map( A1 => n9746, A2 => n9745, A3 => n9744, A4 => 
                           n9743, ZN => n9752);
   U2436 : AOI22_X1 port map( A1 => REGISTERS_18_17_port, A2 => n9835, B1 => 
                           REGISTERS_16_17_port, B2 => n10115, ZN => n9750);
   U2437 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n10166, B1 => 
                           REGISTERS_23_17_port, B2 => n9992, ZN => n9749);
   U2438 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n10165, B1 => 
                           REGISTERS_26_17_port, B2 => n10152, ZN => n9748);
   U2439 : AOI22_X1 port map( A1 => REGISTERS_17_17_port, A2 => n10088, B1 => 
                           REGISTERS_25_17_port, B2 => n10151, ZN => n9747);
   U2440 : NAND4_X1 port map( A1 => n9750, A2 => n9749, A3 => n9748, A4 => 
                           n9747, ZN => n9751);
   U2441 : NOR2_X1 port map( A1 => n9752, A2 => n9751, ZN => n9764);
   U2442 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n10052, B1 => 
                           REGISTERS_3_17_port, B2 => n10178, ZN => n9756);
   U2443 : AOI22_X1 port map( A1 => REGISTERS_1_17_port, A2 => n10189, B1 => 
                           REGISTERS_5_17_port, B2 => n10129, ZN => n9755);
   U2444 : AOI22_X1 port map( A1 => REGISTERS_6_17_port, A2 => n10175, B1 => 
                           REGISTERS_7_17_port, B2 => n10176, ZN => n9754);
   U2445 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n10101, B1 => 
                           REGISTERS_2_17_port, B2 => n10184, ZN => n9753);
   U2446 : NAND4_X1 port map( A1 => n9756, A2 => n9755, A3 => n9754, A4 => 
                           n9753, ZN => n9762);
   U2447 : AOI22_X1 port map( A1 => REGISTERS_10_17_port, A2 => n10136, B1 => 
                           REGISTERS_14_17_port, B2 => n10175, ZN => n9760);
   U2448 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n10187, B1 => 
                           REGISTERS_9_17_port, B2 => n10138, ZN => n9759);
   U2449 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n10188, B1 => 
                           REGISTERS_15_17_port, B2 => n10183, ZN => n9758);
   U2450 : AOI22_X1 port map( A1 => REGISTERS_13_17_port, A2 => n10047, B1 => 
                           REGISTERS_8_17_port, B2 => n10177, ZN => n9757);
   U2451 : NAND4_X1 port map( A1 => n9760, A2 => n9759, A3 => n9758, A4 => 
                           n9757, ZN => n9761);
   U2452 : AOI22_X1 port map( A1 => n10034, A2 => n9762, B1 => n10032, B2 => 
                           n9761, ZN => n9763);
   U2453 : OAI21_X1 port map( B1 => n10201, B2 => n9764, A => n9763, ZN => N402
                           );
   U2454 : AOI22_X1 port map( A1 => REGISTERS_23_16_port, A2 => n9992, B1 => 
                           REGISTERS_21_16_port, B2 => n10161, ZN => n9768);
   U2455 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n10067, B1 => 
                           REGISTERS_30_16_port, B2 => n10150, ZN => n9767);
   U2456 : AOI22_X1 port map( A1 => REGISTERS_31_16_port, A2 => n10061, B1 => 
                           REGISTERS_25_16_port, B2 => n10151, ZN => n9766);
   U2457 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n10155, B1 => 
                           REGISTERS_17_16_port, B2 => n10088, ZN => n9765);
   U2458 : NAND4_X1 port map( A1 => n9768, A2 => n9767, A3 => n9766, A4 => 
                           n9765, ZN => n9774);
   U2459 : AOI22_X1 port map( A1 => REGISTERS_22_16_port, A2 => n10163, B1 => 
                           REGISTERS_28_16_port, B2 => n10166, ZN => n9772);
   U2460 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n10165, B1 => 
                           REGISTERS_18_16_port, B2 => n10154, ZN => n9771);
   U2461 : AOI22_X1 port map( A1 => REGISTERS_27_16_port, A2 => n10168, B1 => 
                           REGISTERS_16_16_port, B2 => n10115, ZN => n9770);
   U2462 : AOI22_X1 port map( A1 => REGISTERS_26_16_port, A2 => n10152, B1 => 
                           REGISTERS_29_16_port, B2 => n10149, ZN => n9769);
   U2463 : NAND4_X1 port map( A1 => n9772, A2 => n9771, A3 => n9770, A4 => 
                           n9769, ZN => n9773);
   U2464 : NOR2_X1 port map( A1 => n9774, A2 => n9773, ZN => n9786);
   U2465 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n10139, B1 => 
                           REGISTERS_6_16_port, B2 => n10175, ZN => n9778);
   U2466 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n10137, B1 => 
                           REGISTERS_7_16_port, B2 => n10176, ZN => n9777);
   U2467 : AOI22_X1 port map( A1 => REGISTERS_5_16_port, A2 => n10129, B1 => 
                           REGISTERS_0_16_port, B2 => n10052, ZN => n9776);
   U2468 : AOI22_X1 port map( A1 => REGISTERS_2_16_port, A2 => n10184, B1 => 
                           REGISTERS_1_16_port, B2 => n10189, ZN => n9775);
   U2469 : NAND4_X1 port map( A1 => n9778, A2 => n9777, A3 => n9776, A4 => 
                           n9775, ZN => n9784);
   U2470 : AOI22_X1 port map( A1 => REGISTERS_14_16_port, A2 => n10175, B1 => 
                           REGISTERS_11_16_port, B2 => n10187, ZN => n9782);
   U2471 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n10176, B1 => 
                           REGISTERS_9_16_port, B2 => n10138, ZN => n9781);
   U2472 : AOI22_X1 port map( A1 => REGISTERS_10_16_port, A2 => n10102, B1 => 
                           REGISTERS_13_16_port, B2 => n10190, ZN => n9780);
   U2473 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n10185, B1 => 
                           REGISTERS_12_16_port, B2 => n10139, ZN => n9779);
   U2474 : NAND4_X1 port map( A1 => n9782, A2 => n9781, A3 => n9780, A4 => 
                           n9779, ZN => n9783);
   U2475 : AOI22_X1 port map( A1 => n10034, A2 => n9784, B1 => n10032, B2 => 
                           n9783, ZN => n9785);
   U2476 : OAI21_X1 port map( B1 => n10201, B2 => n9786, A => n9785, ZN => N401
                           );
   U2477 : AOI22_X1 port map( A1 => REGISTERS_31_15_port, A2 => n10061, B1 => 
                           REGISTERS_16_15_port, B2 => n10153, ZN => n9790);
   U2478 : AOI22_X1 port map( A1 => REGISTERS_22_15_port, A2 => n10087, B1 => 
                           REGISTERS_18_15_port, B2 => n10154, ZN => n9789);
   U2479 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n9921, B1 => 
                           REGISTERS_27_15_port, B2 => n10094, ZN => n9788);
   U2480 : AOI22_X1 port map( A1 => REGISTERS_17_15_port, A2 => n10088, B1 => 
                           REGISTERS_26_15_port, B2 => n10152, ZN => n9787);
   U2481 : NAND4_X1 port map( A1 => n9790, A2 => n9789, A3 => n9788, A4 => 
                           n9787, ZN => n9796);
   U2482 : AOI22_X1 port map( A1 => REGISTERS_21_15_port, A2 => n10161, B1 => 
                           REGISTERS_28_15_port, B2 => n10121, ZN => n9794);
   U2483 : AOI22_X1 port map( A1 => REGISTERS_30_15_port, A2 => n10150, B1 => 
                           REGISTERS_23_15_port, B2 => n9992, ZN => n9793);
   U2484 : AOI22_X1 port map( A1 => REGISTERS_25_15_port, A2 => n10151, B1 => 
                           REGISTERS_19_15_port, B2 => n10012, ZN => n9792);
   U2485 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n10067, B1 => 
                           REGISTERS_24_15_port, B2 => n10066, ZN => n9791);
   U2486 : NAND4_X1 port map( A1 => n9794, A2 => n9793, A3 => n9792, A4 => 
                           n9791, ZN => n9795);
   U2487 : NOR2_X1 port map( A1 => n9796, A2 => n9795, ZN => n9808);
   U2488 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n10131, B1 => 
                           REGISTERS_1_15_port, B2 => n10189, ZN => n9800);
   U2489 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n10188, B1 => 
                           REGISTERS_5_15_port, B2 => n10129, ZN => n9799);
   U2490 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n10177, B1 => 
                           REGISTERS_6_15_port, B2 => n10078, ZN => n9798);
   U2491 : AOI22_X1 port map( A1 => REGISTERS_3_15_port, A2 => n10178, B1 => 
                           REGISTERS_2_15_port, B2 => n10102, ZN => n9797);
   U2492 : NAND4_X1 port map( A1 => n9800, A2 => n9799, A3 => n9798, A4 => 
                           n9797, ZN => n9806);
   U2493 : AOI22_X1 port map( A1 => REGISTERS_10_15_port, A2 => n10136, B1 => 
                           REGISTERS_13_15_port, B2 => n10047, ZN => n9804);
   U2494 : AOI22_X1 port map( A1 => REGISTERS_11_15_port, A2 => n10137, B1 => 
                           REGISTERS_8_15_port, B2 => n10052, ZN => n9803);
   U2495 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n10101, B1 => 
                           REGISTERS_14_15_port, B2 => n10175, ZN => n9802);
   U2496 : AOI22_X1 port map( A1 => REGISTERS_9_15_port, A2 => n10138, B1 => 
                           REGISTERS_15_15_port, B2 => n10176, ZN => n9801);
   U2497 : NAND4_X1 port map( A1 => n9804, A2 => n9803, A3 => n9802, A4 => 
                           n9801, ZN => n9805);
   U2498 : AOI22_X1 port map( A1 => n10034, A2 => n9806, B1 => n10032, B2 => 
                           n9805, ZN => n9807);
   U2499 : OAI21_X1 port map( B1 => n10148, B2 => n9808, A => n9807, ZN => N400
                           );
   U2500 : AOI22_X1 port map( A1 => REGISTERS_27_14_port, A2 => n10168, B1 => 
                           REGISTERS_20_14_port, B2 => n10067, ZN => n9812);
   U2501 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n9921, B1 => 
                           REGISTERS_31_14_port, B2 => n10164, ZN => n9811);
   U2502 : AOI22_X1 port map( A1 => REGISTERS_21_14_port, A2 => n10161, B1 => 
                           REGISTERS_18_14_port, B2 => n10154, ZN => n9810);
   U2503 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n10166, B1 => 
                           REGISTERS_24_14_port, B2 => n10066, ZN => n9809);
   U2504 : NAND4_X1 port map( A1 => n9812, A2 => n9811, A3 => n9810, A4 => 
                           n9809, ZN => n9818);
   U2505 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n10153, B1 => 
                           REGISTERS_17_14_port, B2 => n10088, ZN => n9816);
   U2506 : AOI22_X1 port map( A1 => REGISTERS_22_14_port, A2 => n10087, B1 => 
                           REGISTERS_19_14_port, B2 => n10012, ZN => n9815);
   U2507 : AOI22_X1 port map( A1 => REGISTERS_23_14_port, A2 => n9992, B1 => 
                           REGISTERS_25_14_port, B2 => n10151, ZN => n9814);
   U2508 : AOI22_X1 port map( A1 => REGISTERS_26_14_port, A2 => n10152, B1 => 
                           REGISTERS_30_14_port, B2 => n10150, ZN => n9813);
   U2509 : NAND4_X1 port map( A1 => n9816, A2 => n9815, A3 => n9814, A4 => 
                           n9813, ZN => n9817);
   U2510 : NOR2_X1 port map( A1 => n9818, A2 => n9817, ZN => n9830);
   U2511 : AOI22_X1 port map( A1 => REGISTERS_5_14_port, A2 => n10190, B1 => 
                           REGISTERS_3_14_port, B2 => n10178, ZN => n9822);
   U2512 : AOI22_X1 port map( A1 => REGISTERS_1_14_port, A2 => n10130, B1 => 
                           REGISTERS_4_14_port, B2 => n10188, ZN => n9821);
   U2513 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n10052, B1 => 
                           REGISTERS_2_14_port, B2 => n10102, ZN => n9820);
   U2514 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n10183, B1 => 
                           REGISTERS_6_14_port, B2 => n10078, ZN => n9819);
   U2515 : NAND4_X1 port map( A1 => n9822, A2 => n9821, A3 => n9820, A4 => 
                           n9819, ZN => n9828);
   U2516 : AOI22_X1 port map( A1 => REGISTERS_15_14_port, A2 => n10131, B1 => 
                           REGISTERS_12_14_port, B2 => n10139, ZN => n9826);
   U2517 : AOI22_X1 port map( A1 => REGISTERS_13_14_port, A2 => n10047, B1 => 
                           REGISTERS_14_14_port, B2 => n10078, ZN => n9825);
   U2518 : AOI22_X1 port map( A1 => REGISTERS_10_14_port, A2 => n10184, B1 => 
                           REGISTERS_8_14_port, B2 => n10177, ZN => n9824);
   U2519 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n10178, B1 => 
                           REGISTERS_9_14_port, B2 => n10189, ZN => n9823);
   U2520 : NAND4_X1 port map( A1 => n9826, A2 => n9825, A3 => n9824, A4 => 
                           n9823, ZN => n9827);
   U2521 : AOI22_X1 port map( A1 => n10034, A2 => n9828, B1 => n10032, B2 => 
                           n9827, ZN => n9829);
   U2522 : OAI21_X1 port map( B1 => n10201, B2 => n9830, A => n9829, ZN => N399
                           );
   U2523 : AOI22_X1 port map( A1 => REGISTERS_31_13_port, A2 => n10164, B1 => 
                           REGISTERS_20_13_port, B2 => n10067, ZN => n9834);
   U2524 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n10165, B1 => 
                           REGISTERS_17_13_port, B2 => n10088, ZN => n9833);
   U2525 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n10115, B1 => 
                           REGISTERS_19_13_port, B2 => n10155, ZN => n9832);
   U2526 : AOI22_X1 port map( A1 => REGISTERS_25_13_port, A2 => n10151, B1 => 
                           REGISTERS_27_13_port, B2 => n10094, ZN => n9831);
   U2527 : NAND4_X1 port map( A1 => n9834, A2 => n9833, A3 => n9832, A4 => 
                           n9831, ZN => n9841);
   U2528 : AOI22_X1 port map( A1 => REGISTERS_18_13_port, A2 => n9835, B1 => 
                           REGISTERS_28_13_port, B2 => n10121, ZN => n9839);
   U2529 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n10149, B1 => 
                           REGISTERS_23_13_port, B2 => n10167, ZN => n9838);
   U2530 : AOI22_X1 port map( A1 => REGISTERS_26_13_port, A2 => n10152, B1 => 
                           REGISTERS_22_13_port, B2 => n10163, ZN => n9837);
   U2531 : AOI22_X1 port map( A1 => REGISTERS_21_13_port, A2 => n10161, B1 => 
                           REGISTERS_30_13_port, B2 => n10150, ZN => n9836);
   U2532 : NAND4_X1 port map( A1 => n9839, A2 => n9838, A3 => n9837, A4 => 
                           n9836, ZN => n9840);
   U2533 : NOR2_X1 port map( A1 => n9841, A2 => n9840, ZN => n9853);
   U2534 : AOI22_X1 port map( A1 => REGISTERS_1_13_port, A2 => n10189, B1 => 
                           REGISTERS_7_13_port, B2 => n10183, ZN => n9845);
   U2535 : AOI22_X1 port map( A1 => REGISTERS_2_13_port, A2 => n10102, B1 => 
                           REGISTERS_0_13_port, B2 => n10052, ZN => n9844);
   U2536 : AOI22_X1 port map( A1 => REGISTERS_3_13_port, A2 => n10187, B1 => 
                           REGISTERS_5_13_port, B2 => n10047, ZN => n9843);
   U2537 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n10101, B1 => 
                           REGISTERS_6_13_port, B2 => n10078, ZN => n9842);
   U2538 : NAND4_X1 port map( A1 => n9845, A2 => n9844, A3 => n9843, A4 => 
                           n9842, ZN => n9851);
   U2539 : AOI22_X1 port map( A1 => REGISTERS_13_13_port, A2 => n10190, B1 => 
                           REGISTERS_15_13_port, B2 => n10176, ZN => n9849);
   U2540 : AOI22_X1 port map( A1 => REGISTERS_11_13_port, A2 => n10187, B1 => 
                           REGISTERS_14_13_port, B2 => n10175, ZN => n9848);
   U2541 : AOI22_X1 port map( A1 => REGISTERS_9_13_port, A2 => n10130, B1 => 
                           REGISTERS_8_13_port, B2 => n10185, ZN => n9847);
   U2542 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n10188, B1 => 
                           REGISTERS_10_13_port, B2 => n10184, ZN => n9846);
   U2543 : NAND4_X1 port map( A1 => n9849, A2 => n9848, A3 => n9847, A4 => 
                           n9846, ZN => n9850);
   U2544 : AOI22_X1 port map( A1 => n10034, A2 => n9851, B1 => n10032, B2 => 
                           n9850, ZN => n9852);
   U2545 : OAI21_X1 port map( B1 => n10148, B2 => n9853, A => n9852, ZN => N398
                           );
   U2546 : AOI22_X1 port map( A1 => REGISTERS_21_12_port, A2 => n10161, B1 => 
                           REGISTERS_24_12_port, B2 => n10066, ZN => n9857);
   U2547 : AOI22_X1 port map( A1 => REGISTERS_27_12_port, A2 => n10094, B1 => 
                           REGISTERS_19_12_port, B2 => n10155, ZN => n9856);
   U2548 : AOI22_X1 port map( A1 => REGISTERS_23_12_port, A2 => n10167, B1 => 
                           REGISTERS_28_12_port, B2 => n10121, ZN => n9855);
   U2549 : AOI22_X1 port map( A1 => REGISTERS_26_12_port, A2 => n10152, B1 => 
                           REGISTERS_18_12_port, B2 => n10154, ZN => n9854);
   U2550 : NAND4_X1 port map( A1 => n9857, A2 => n9856, A3 => n9855, A4 => 
                           n9854, ZN => n9863);
   U2551 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n10067, B1 => 
                           REGISTERS_29_12_port, B2 => n10149, ZN => n9861);
   U2552 : AOI22_X1 port map( A1 => REGISTERS_25_12_port, A2 => n10093, B1 => 
                           REGISTERS_31_12_port, B2 => n10164, ZN => n9860);
   U2553 : AOI22_X1 port map( A1 => REGISTERS_30_12_port, A2 => n10116, B1 => 
                           REGISTERS_22_12_port, B2 => n10163, ZN => n9859);
   U2554 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n10115, B1 => 
                           REGISTERS_17_12_port, B2 => n10156, ZN => n9858);
   U2555 : NAND4_X1 port map( A1 => n9861, A2 => n9860, A3 => n9859, A4 => 
                           n9858, ZN => n9862);
   U2556 : NOR2_X1 port map( A1 => n9863, A2 => n9862, ZN => n9875);
   U2557 : AOI22_X1 port map( A1 => REGISTERS_2_12_port, A2 => n10136, B1 => 
                           REGISTERS_1_12_port, B2 => n10138, ZN => n9867);
   U2558 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n10176, B1 => 
                           REGISTERS_6_12_port, B2 => n10175, ZN => n9866);
   U2559 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n10188, B1 => 
                           REGISTERS_5_12_port, B2 => n10129, ZN => n9865);
   U2560 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n10185, B1 => 
                           REGISTERS_3_12_port, B2 => n10187, ZN => n9864);
   U2561 : NAND4_X1 port map( A1 => n9867, A2 => n9866, A3 => n9865, A4 => 
                           n9864, ZN => n9873);
   U2562 : AOI22_X1 port map( A1 => REGISTERS_14_12_port, A2 => n10186, B1 => 
                           REGISTERS_15_12_port, B2 => n10183, ZN => n9871);
   U2563 : AOI22_X1 port map( A1 => REGISTERS_13_12_port, A2 => n10190, B1 => 
                           REGISTERS_8_12_port, B2 => n10052, ZN => n9870);
   U2564 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n10188, B1 => 
                           REGISTERS_11_12_port, B2 => n10137, ZN => n9869);
   U2565 : AOI22_X1 port map( A1 => REGISTERS_10_12_port, A2 => n10184, B1 => 
                           REGISTERS_9_12_port, B2 => n10189, ZN => n9868);
   U2566 : NAND4_X1 port map( A1 => n9871, A2 => n9870, A3 => n9869, A4 => 
                           n9868, ZN => n9872);
   U2567 : AOI22_X1 port map( A1 => n10034, A2 => n9873, B1 => n10032, B2 => 
                           n9872, ZN => n9874);
   U2568 : OAI21_X1 port map( B1 => n10201, B2 => n9875, A => n9874, ZN => N397
                           );
   U2569 : AOI22_X1 port map( A1 => REGISTERS_27_11_port, A2 => n10094, B1 => 
                           REGISTERS_18_11_port, B2 => n10154, ZN => n9879);
   U2570 : AOI22_X1 port map( A1 => REGISTERS_22_11_port, A2 => n10087, B1 => 
                           REGISTERS_28_11_port, B2 => n10121, ZN => n9878);
   U2571 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n10167, B1 => 
                           REGISTERS_20_11_port, B2 => n10067, ZN => n9877);
   U2572 : AOI22_X1 port map( A1 => REGISTERS_17_11_port, A2 => n10088, B1 => 
                           REGISTERS_29_11_port, B2 => n10149, ZN => n9876);
   U2573 : NAND4_X1 port map( A1 => n9879, A2 => n9878, A3 => n9877, A4 => 
                           n9876, ZN => n9885);
   U2574 : AOI22_X1 port map( A1 => REGISTERS_31_11_port, A2 => n10164, B1 => 
                           REGISTERS_25_11_port, B2 => n10151, ZN => n9883);
   U2575 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n10165, B1 => 
                           REGISTERS_21_11_port, B2 => n10161, ZN => n9882);
   U2576 : AOI22_X1 port map( A1 => REGISTERS_30_11_port, A2 => n10150, B1 => 
                           REGISTERS_26_11_port, B2 => n10152, ZN => n9881);
   U2577 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n10155, B1 => 
                           REGISTERS_16_11_port, B2 => n10115, ZN => n9880);
   U2578 : NAND4_X1 port map( A1 => n9883, A2 => n9882, A3 => n9881, A4 => 
                           n9880, ZN => n9884);
   U2579 : NOR2_X1 port map( A1 => n9885, A2 => n9884, ZN => n9897);
   U2580 : AOI22_X1 port map( A1 => REGISTERS_6_11_port, A2 => n10186, B1 => 
                           REGISTERS_3_11_port, B2 => n10187, ZN => n9889);
   U2581 : AOI22_X1 port map( A1 => REGISTERS_5_11_port, A2 => n10190, B1 => 
                           REGISTERS_7_11_port, B2 => n10176, ZN => n9888);
   U2582 : AOI22_X1 port map( A1 => REGISTERS_2_11_port, A2 => n10102, B1 => 
                           REGISTERS_0_11_port, B2 => n10185, ZN => n9887);
   U2583 : AOI22_X1 port map( A1 => REGISTERS_1_11_port, A2 => n10189, B1 => 
                           REGISTERS_4_11_port, B2 => n10188, ZN => n9886);
   U2584 : NAND4_X1 port map( A1 => n9889, A2 => n9888, A3 => n9887, A4 => 
                           n9886, ZN => n9895);
   U2585 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n10177, B1 => 
                           REGISTERS_15_11_port, B2 => n10183, ZN => n9893);
   U2586 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n10188, B1 => 
                           REGISTERS_11_11_port, B2 => n10137, ZN => n9892);
   U2587 : AOI22_X1 port map( A1 => REGISTERS_10_11_port, A2 => n10184, B1 => 
                           REGISTERS_9_11_port, B2 => n10138, ZN => n9891);
   U2588 : AOI22_X1 port map( A1 => REGISTERS_13_11_port, A2 => n10190, B1 => 
                           REGISTERS_14_11_port, B2 => n10175, ZN => n9890);
   U2589 : NAND4_X1 port map( A1 => n9893, A2 => n9892, A3 => n9891, A4 => 
                           n9890, ZN => n9894);
   U2590 : AOI22_X1 port map( A1 => n10034, A2 => n9895, B1 => n10032, B2 => 
                           n9894, ZN => n9896);
   U2591 : OAI21_X1 port map( B1 => n10201, B2 => n9897, A => n9896, ZN => N396
                           );
   U2592 : AOI22_X1 port map( A1 => REGISTERS_21_10_port, A2 => n9898, B1 => 
                           REGISTERS_20_10_port, B2 => n10067, ZN => n9902);
   U2593 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n10165, B1 => 
                           REGISTERS_28_10_port, B2 => n10121, ZN => n9901);
   U2594 : AOI22_X1 port map( A1 => REGISTERS_31_10_port, A2 => n10164, B1 => 
                           REGISTERS_16_10_port, B2 => n10153, ZN => n9900);
   U2595 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n10094, B1 => 
                           REGISTERS_25_10_port, B2 => n10151, ZN => n9899);
   U2596 : NAND4_X1 port map( A1 => n9902, A2 => n9901, A3 => n9900, A4 => 
                           n9899, ZN => n9908);
   U2597 : AOI22_X1 port map( A1 => REGISTERS_22_10_port, A2 => n10087, B1 => 
                           REGISTERS_26_10_port, B2 => n10152, ZN => n9906);
   U2598 : AOI22_X1 port map( A1 => REGISTERS_23_10_port, A2 => n10167, B1 => 
                           REGISTERS_18_10_port, B2 => n10154, ZN => n9905);
   U2599 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n10155, B1 => 
                           REGISTERS_29_10_port, B2 => n10149, ZN => n9904);
   U2600 : AOI22_X1 port map( A1 => REGISTERS_17_10_port, A2 => n10088, B1 => 
                           REGISTERS_30_10_port, B2 => n10150, ZN => n9903);
   U2601 : NAND4_X1 port map( A1 => n9906, A2 => n9905, A3 => n9904, A4 => 
                           n9903, ZN => n9907);
   U2602 : NOR2_X1 port map( A1 => n9908, A2 => n9907, ZN => n9920);
   U2603 : AOI22_X1 port map( A1 => REGISTERS_1_10_port, A2 => n10130, B1 => 
                           REGISTERS_4_10_port, B2 => n10139, ZN => n9912);
   U2604 : AOI22_X1 port map( A1 => REGISTERS_2_10_port, A2 => n10184, B1 => 
                           REGISTERS_6_10_port, B2 => n10078, ZN => n9911);
   U2605 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n10052, B1 => 
                           REGISTERS_3_10_port, B2 => n10178, ZN => n9910);
   U2606 : AOI22_X1 port map( A1 => REGISTERS_5_10_port, A2 => n10190, B1 => 
                           REGISTERS_7_10_port, B2 => n10131, ZN => n9909);
   U2607 : NAND4_X1 port map( A1 => n9912, A2 => n9911, A3 => n9910, A4 => 
                           n9909, ZN => n9918);
   U2608 : AOI22_X1 port map( A1 => REGISTERS_9_10_port, A2 => n10189, B1 => 
                           REGISTERS_14_10_port, B2 => n10078, ZN => n9916);
   U2609 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n10178, B1 => 
                           REGISTERS_8_10_port, B2 => n10185, ZN => n9915);
   U2610 : AOI22_X1 port map( A1 => REGISTERS_15_10_port, A2 => n10176, B1 => 
                           REGISTERS_12_10_port, B2 => n10188, ZN => n9914);
   U2611 : AOI22_X1 port map( A1 => REGISTERS_10_10_port, A2 => n10184, B1 => 
                           REGISTERS_13_10_port, B2 => n10129, ZN => n9913);
   U2612 : NAND4_X1 port map( A1 => n9916, A2 => n9915, A3 => n9914, A4 => 
                           n9913, ZN => n9917);
   U2613 : AOI22_X1 port map( A1 => n10034, A2 => n9918, B1 => n10032, B2 => 
                           n9917, ZN => n9919);
   U2614 : OAI21_X1 port map( B1 => n10201, B2 => n9920, A => n9919, ZN => N395
                           );
   U2615 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n9921, B1 => 
                           REGISTERS_30_9_port, B2 => n10116, ZN => n9925);
   U2616 : AOI22_X1 port map( A1 => REGISTERS_17_9_port, A2 => n10088, B1 => 
                           REGISTERS_24_9_port, B2 => n10066, ZN => n9924);
   U2617 : AOI22_X1 port map( A1 => REGISTERS_31_9_port, A2 => n10164, B1 => 
                           REGISTERS_26_9_port, B2 => n10122, ZN => n9923);
   U2618 : AOI22_X1 port map( A1 => REGISTERS_19_9_port, A2 => n10155, B1 => 
                           REGISTERS_23_9_port, B2 => n10167, ZN => n9922);
   U2619 : NAND4_X1 port map( A1 => n9925, A2 => n9924, A3 => n9923, A4 => 
                           n9922, ZN => n9931);
   U2620 : AOI22_X1 port map( A1 => REGISTERS_21_9_port, A2 => n10161, B1 => 
                           REGISTERS_18_9_port, B2 => n10154, ZN => n9929);
   U2621 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n10115, B1 => 
                           REGISTERS_22_9_port, B2 => n10163, ZN => n9928);
   U2622 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n10067, B1 => 
                           REGISTERS_25_9_port, B2 => n10151, ZN => n9927);
   U2623 : AOI22_X1 port map( A1 => REGISTERS_27_9_port, A2 => n10094, B1 => 
                           REGISTERS_28_9_port, B2 => n10121, ZN => n9926);
   U2624 : NAND4_X1 port map( A1 => n9929, A2 => n9928, A3 => n9927, A4 => 
                           n9926, ZN => n9930);
   U2625 : NOR2_X1 port map( A1 => n9931, A2 => n9930, ZN => n9943);
   U2626 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n10177, B1 => 
                           REGISTERS_5_9_port, B2 => n10047, ZN => n9935);
   U2627 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n10187, B1 => 
                           REGISTERS_4_9_port, B2 => n10139, ZN => n9934);
   U2628 : AOI22_X1 port map( A1 => REGISTERS_1_9_port, A2 => n10138, B1 => 
                           REGISTERS_2_9_port, B2 => n10136, ZN => n9933);
   U2629 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n10183, B1 => 
                           REGISTERS_6_9_port, B2 => n10078, ZN => n9932);
   U2630 : NAND4_X1 port map( A1 => n9935, A2 => n9934, A3 => n9933, A4 => 
                           n9932, ZN => n9941);
   U2631 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n10177, B1 => 
                           REGISTERS_13_9_port, B2 => n10129, ZN => n9939);
   U2632 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n10131, B1 => 
                           REGISTERS_12_9_port, B2 => n10188, ZN => n9938);
   U2633 : AOI22_X1 port map( A1 => REGISTERS_14_9_port, A2 => n10186, B1 => 
                           REGISTERS_10_9_port, B2 => n10102, ZN => n9937);
   U2634 : AOI22_X1 port map( A1 => REGISTERS_11_9_port, A2 => n10137, B1 => 
                           REGISTERS_9_9_port, B2 => n10130, ZN => n9936);
   U2635 : NAND4_X1 port map( A1 => n9939, A2 => n9938, A3 => n9937, A4 => 
                           n9936, ZN => n9940);
   U2636 : AOI22_X1 port map( A1 => n10034, A2 => n9941, B1 => n10032, B2 => 
                           n9940, ZN => n9942);
   U2637 : OAI21_X1 port map( B1 => n10148, B2 => n9943, A => n9942, ZN => N394
                           );
   U2638 : AOI22_X1 port map( A1 => REGISTERS_22_8_port, A2 => n10087, B1 => 
                           REGISTERS_26_8_port, B2 => n10122, ZN => n9947);
   U2639 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n10155, B1 => 
                           REGISTERS_31_8_port, B2 => n10061, ZN => n9946);
   U2640 : AOI22_X1 port map( A1 => REGISTERS_25_8_port, A2 => n10151, B1 => 
                           REGISTERS_27_8_port, B2 => n10168, ZN => n9945);
   U2641 : AOI22_X1 port map( A1 => REGISTERS_30_8_port, A2 => n10150, B1 => 
                           REGISTERS_24_8_port, B2 => n10165, ZN => n9944);
   U2642 : NAND4_X1 port map( A1 => n9947, A2 => n9946, A3 => n9945, A4 => 
                           n9944, ZN => n9953);
   U2643 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n10149, B1 => 
                           REGISTERS_18_8_port, B2 => n10154, ZN => n9951);
   U2644 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n10067, B1 => 
                           REGISTERS_21_8_port, B2 => n10161, ZN => n9950);
   U2645 : AOI22_X1 port map( A1 => REGISTERS_17_8_port, A2 => n10088, B1 => 
                           REGISTERS_16_8_port, B2 => n10153, ZN => n9949);
   U2646 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n10167, B1 => 
                           REGISTERS_28_8_port, B2 => n10121, ZN => n9948);
   U2647 : NAND4_X1 port map( A1 => n9951, A2 => n9950, A3 => n9949, A4 => 
                           n9948, ZN => n9952);
   U2648 : NOR2_X1 port map( A1 => n9953, A2 => n9952, ZN => n9965);
   U2649 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n10183, B1 => 
                           REGISTERS_5_8_port, B2 => n10129, ZN => n9957);
   U2650 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n10177, B1 => 
                           REGISTERS_6_8_port, B2 => n10175, ZN => n9956);
   U2651 : AOI22_X1 port map( A1 => REGISTERS_3_8_port, A2 => n10187, B1 => 
                           REGISTERS_1_8_port, B2 => n10189, ZN => n9955);
   U2652 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n10139, B1 => 
                           REGISTERS_2_8_port, B2 => n10102, ZN => n9954);
   U2653 : NAND4_X1 port map( A1 => n9957, A2 => n9956, A3 => n9955, A4 => 
                           n9954, ZN => n9963);
   U2654 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n10176, B1 => 
                           REGISTERS_13_8_port, B2 => n10047, ZN => n9961);
   U2655 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n10137, B1 => 
                           REGISTERS_14_8_port, B2 => n10078, ZN => n9960);
   U2656 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n10177, B1 => 
                           REGISTERS_9_8_port, B2 => n10138, ZN => n9959);
   U2657 : AOI22_X1 port map( A1 => REGISTERS_10_8_port, A2 => n10184, B1 => 
                           REGISTERS_12_8_port, B2 => n10139, ZN => n9958);
   U2658 : NAND4_X1 port map( A1 => n9961, A2 => n9960, A3 => n9959, A4 => 
                           n9958, ZN => n9962);
   U2659 : AOI22_X1 port map( A1 => n10034, A2 => n9963, B1 => n10032, B2 => 
                           n9962, ZN => n9964);
   U2660 : OAI21_X1 port map( B1 => n10201, B2 => n9965, A => n9964, ZN => N393
                           );
   U2661 : AOI22_X1 port map( A1 => REGISTERS_25_7_port, A2 => n10151, B1 => 
                           REGISTERS_22_7_port, B2 => n10087, ZN => n9969);
   U2662 : AOI22_X1 port map( A1 => REGISTERS_31_7_port, A2 => n10164, B1 => 
                           REGISTERS_27_7_port, B2 => n10168, ZN => n9968);
   U2663 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n10165, B1 => 
                           REGISTERS_20_7_port, B2 => n10162, ZN => n9967);
   U2664 : AOI22_X1 port map( A1 => REGISTERS_18_7_port, A2 => n10154, B1 => 
                           REGISTERS_28_7_port, B2 => n10121, ZN => n9966);
   U2665 : NAND4_X1 port map( A1 => n9969, A2 => n9968, A3 => n9967, A4 => 
                           n9966, ZN => n9975);
   U2666 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n10115, B1 => 
                           REGISTERS_19_7_port, B2 => n10155, ZN => n9973);
   U2667 : AOI22_X1 port map( A1 => REGISTERS_26_7_port, A2 => n10152, B1 => 
                           REGISTERS_17_7_port, B2 => n10156, ZN => n9972);
   U2668 : AOI22_X1 port map( A1 => REGISTERS_21_7_port, A2 => n10161, B1 => 
                           REGISTERS_29_7_port, B2 => n10149, ZN => n9971);
   U2669 : AOI22_X1 port map( A1 => REGISTERS_30_7_port, A2 => n10150, B1 => 
                           REGISTERS_23_7_port, B2 => n10167, ZN => n9970);
   U2670 : NAND4_X1 port map( A1 => n9973, A2 => n9972, A3 => n9971, A4 => 
                           n9970, ZN => n9974);
   U2671 : NOR2_X1 port map( A1 => n9975, A2 => n9974, ZN => n9987);
   U2672 : AOI22_X1 port map( A1 => REGISTERS_2_7_port, A2 => n10184, B1 => 
                           REGISTERS_7_7_port, B2 => n10183, ZN => n9979);
   U2673 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n10177, B1 => 
                           REGISTERS_3_7_port, B2 => n10137, ZN => n9978);
   U2674 : AOI22_X1 port map( A1 => REGISTERS_6_7_port, A2 => n10186, B1 => 
                           REGISTERS_5_7_port, B2 => n10129, ZN => n9977);
   U2675 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n10139, B1 => 
                           REGISTERS_1_7_port, B2 => n10189, ZN => n9976);
   U2676 : NAND4_X1 port map( A1 => n9979, A2 => n9978, A3 => n9977, A4 => 
                           n9976, ZN => n9985);
   U2677 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n10177, B1 => 
                           REGISTERS_15_7_port, B2 => n10176, ZN => n9983);
   U2678 : AOI22_X1 port map( A1 => REGISTERS_14_7_port, A2 => n10186, B1 => 
                           REGISTERS_9_7_port, B2 => n10138, ZN => n9982);
   U2679 : AOI22_X1 port map( A1 => REGISTERS_10_7_port, A2 => n10184, B1 => 
                           REGISTERS_13_7_port, B2 => n10047, ZN => n9981);
   U2680 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n10137, B1 => 
                           REGISTERS_12_7_port, B2 => n10139, ZN => n9980);
   U2681 : NAND4_X1 port map( A1 => n9983, A2 => n9982, A3 => n9981, A4 => 
                           n9980, ZN => n9984);
   U2682 : AOI22_X1 port map( A1 => n10034, A2 => n9985, B1 => n10032, B2 => 
                           n9984, ZN => n9986);
   U2683 : OAI21_X1 port map( B1 => n10148, B2 => n9987, A => n9986, ZN => N392
                           );
   U2684 : AOI22_X1 port map( A1 => REGISTERS_25_6_port, A2 => n10151, B1 => 
                           REGISTERS_26_6_port, B2 => n10122, ZN => n9991);
   U2685 : AOI22_X1 port map( A1 => REGISTERS_31_6_port, A2 => n10164, B1 => 
                           REGISTERS_17_6_port, B2 => n10156, ZN => n9990);
   U2686 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n10115, B1 => 
                           REGISTERS_24_6_port, B2 => n10165, ZN => n9989);
   U2687 : AOI22_X1 port map( A1 => REGISTERS_18_6_port, A2 => n10154, B1 => 
                           REGISTERS_20_6_port, B2 => n10162, ZN => n9988);
   U2688 : NAND4_X1 port map( A1 => n9991, A2 => n9990, A3 => n9989, A4 => 
                           n9988, ZN => n9998);
   U2689 : AOI22_X1 port map( A1 => REGISTERS_27_6_port, A2 => n10094, B1 => 
                           REGISTERS_28_6_port, B2 => n10121, ZN => n9996);
   U2690 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n10149, B1 => 
                           REGISTERS_21_6_port, B2 => n10161, ZN => n9995);
   U2691 : AOI22_X1 port map( A1 => REGISTERS_23_6_port, A2 => n9992, B1 => 
                           REGISTERS_30_6_port, B2 => n10116, ZN => n9994);
   U2692 : AOI22_X1 port map( A1 => REGISTERS_19_6_port, A2 => n10012, B1 => 
                           REGISTERS_22_6_port, B2 => n10087, ZN => n9993);
   U2693 : NAND4_X1 port map( A1 => n9996, A2 => n9995, A3 => n9994, A4 => 
                           n9993, ZN => n9997);
   U2694 : NOR2_X1 port map( A1 => n9998, A2 => n9997, ZN => n10011);
   U2695 : AOI22_X1 port map( A1 => REGISTERS_1_6_port, A2 => n10130, B1 => 
                           REGISTERS_2_6_port, B2 => n10136, ZN => n10002);
   U2696 : AOI22_X1 port map( A1 => REGISTERS_7_6_port, A2 => n10131, B1 => 
                           REGISTERS_0_6_port, B2 => n10185, ZN => n10001);
   U2697 : AOI22_X1 port map( A1 => REGISTERS_5_6_port, A2 => n10190, B1 => 
                           REGISTERS_4_6_port, B2 => n10101, ZN => n10000);
   U2698 : AOI22_X1 port map( A1 => REGISTERS_3_6_port, A2 => n10137, B1 => 
                           REGISTERS_6_6_port, B2 => n10175, ZN => n9999);
   U2699 : NAND4_X1 port map( A1 => n10002, A2 => n10001, A3 => n10000, A4 => 
                           n9999, ZN => n10008);
   U2700 : AOI22_X1 port map( A1 => REGISTERS_14_6_port, A2 => n10186, B1 => 
                           REGISTERS_9_6_port, B2 => n10138, ZN => n10006);
   U2701 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n10178, B1 => 
                           REGISTERS_12_6_port, B2 => n10101, ZN => n10005);
   U2702 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n10131, B1 => 
                           REGISTERS_8_6_port, B2 => n10052, ZN => n10004);
   U2703 : AOI22_X1 port map( A1 => REGISTERS_10_6_port, A2 => n10184, B1 => 
                           REGISTERS_13_6_port, B2 => n10047, ZN => n10003);
   U2704 : NAND4_X1 port map( A1 => n10006, A2 => n10005, A3 => n10004, A4 => 
                           n10003, ZN => n10007);
   U2705 : AOI22_X1 port map( A1 => n10009, A2 => n10008, B1 => n10032, B2 => 
                           n10007, ZN => n10010);
   U2706 : OAI21_X1 port map( B1 => n10201, B2 => n10011, A => n10010, ZN => 
                           N391);
   U2707 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n10121, B1 => 
                           REGISTERS_29_5_port, B2 => n10149, ZN => n10016);
   U2708 : AOI22_X1 port map( A1 => REGISTERS_22_5_port, A2 => n10087, B1 => 
                           REGISTERS_30_5_port, B2 => n10116, ZN => n10015);
   U2709 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n10115, B1 => 
                           REGISTERS_24_5_port, B2 => n10165, ZN => n10014);
   U2710 : AOI22_X1 port map( A1 => REGISTERS_19_5_port, A2 => n10012, B1 => 
                           REGISTERS_25_5_port, B2 => n10093, ZN => n10013);
   U2711 : NAND4_X1 port map( A1 => n10016, A2 => n10015, A3 => n10014, A4 => 
                           n10013, ZN => n10022);
   U2712 : AOI22_X1 port map( A1 => REGISTERS_18_5_port, A2 => n10154, B1 => 
                           REGISTERS_21_5_port, B2 => n10161, ZN => n10020);
   U2713 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n10167, B1 => 
                           REGISTERS_31_5_port, B2 => n10061, ZN => n10019);
   U2714 : AOI22_X1 port map( A1 => REGISTERS_26_5_port, A2 => n10152, B1 => 
                           REGISTERS_17_5_port, B2 => n10156, ZN => n10018);
   U2715 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n10094, B1 => 
                           REGISTERS_20_5_port, B2 => n10162, ZN => n10017);
   U2716 : NAND4_X1 port map( A1 => n10020, A2 => n10019, A3 => n10018, A4 => 
                           n10017, ZN => n10021);
   U2717 : NOR2_X1 port map( A1 => n10022, A2 => n10021, ZN => n10036);
   U2718 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n10177, B1 => 
                           REGISTERS_5_5_port, B2 => n10047, ZN => n10026);
   U2719 : AOI22_X1 port map( A1 => REGISTERS_6_5_port, A2 => n10186, B1 => 
                           REGISTERS_7_5_port, B2 => n10176, ZN => n10025);
   U2720 : AOI22_X1 port map( A1 => REGISTERS_1_5_port, A2 => n10138, B1 => 
                           REGISTERS_2_5_port, B2 => n10136, ZN => n10024);
   U2721 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n10139, B1 => 
                           REGISTERS_3_5_port, B2 => n10137, ZN => n10023);
   U2722 : NAND4_X1 port map( A1 => n10026, A2 => n10025, A3 => n10024, A4 => 
                           n10023, ZN => n10033);
   U2723 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n10178, B1 => 
                           REGISTERS_13_5_port, B2 => n10129, ZN => n10030);
   U2724 : AOI22_X1 port map( A1 => REGISTERS_10_5_port, A2 => n10184, B1 => 
                           REGISTERS_12_5_port, B2 => n10188, ZN => n10029);
   U2725 : AOI22_X1 port map( A1 => REGISTERS_9_5_port, A2 => n10130, B1 => 
                           REGISTERS_15_5_port, B2 => n10131, ZN => n10028);
   U2726 : AOI22_X1 port map( A1 => REGISTERS_14_5_port, A2 => n10186, B1 => 
                           REGISTERS_8_5_port, B2 => n10052, ZN => n10027);
   U2727 : NAND4_X1 port map( A1 => n10030, A2 => n10029, A3 => n10028, A4 => 
                           n10027, ZN => n10031);
   U2728 : AOI22_X1 port map( A1 => n10034, A2 => n10033, B1 => n10032, B2 => 
                           n10031, ZN => n10035);
   U2729 : OAI21_X1 port map( B1 => n10148, B2 => n10036, A => n10035, ZN => 
                           N390);
   U2730 : AOI22_X1 port map( A1 => REGISTERS_26_4_port, A2 => n10122, B1 => 
                           REGISTERS_18_4_port, B2 => n10154, ZN => n10040);
   U2731 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n10094, B1 => 
                           REGISTERS_19_4_port, B2 => n10155, ZN => n10039);
   U2732 : AOI22_X1 port map( A1 => REGISTERS_21_4_port, A2 => n10161, B1 => 
                           REGISTERS_20_4_port, B2 => n10162, ZN => n10038);
   U2733 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n10066, B1 => 
                           REGISTERS_30_4_port, B2 => n10116, ZN => n10037);
   U2734 : NAND4_X1 port map( A1 => n10040, A2 => n10039, A3 => n10038, A4 => 
                           n10037, ZN => n10046);
   U2735 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n10115, B1 => 
                           REGISTERS_28_4_port, B2 => n10121, ZN => n10044);
   U2736 : AOI22_X1 port map( A1 => REGISTERS_25_4_port, A2 => n10151, B1 => 
                           REGISTERS_29_4_port, B2 => n10149, ZN => n10043);
   U2737 : AOI22_X1 port map( A1 => REGISTERS_31_4_port, A2 => n10164, B1 => 
                           REGISTERS_22_4_port, B2 => n10087, ZN => n10042);
   U2738 : AOI22_X1 port map( A1 => REGISTERS_17_4_port, A2 => n10088, B1 => 
                           REGISTERS_23_4_port, B2 => n10167, ZN => n10041);
   U2739 : NAND4_X1 port map( A1 => n10044, A2 => n10043, A3 => n10042, A4 => 
                           n10041, ZN => n10045);
   U2740 : NOR2_X1 port map( A1 => n10046, A2 => n10045, ZN => n10060);
   U2741 : AOI22_X1 port map( A1 => REGISTERS_3_4_port, A2 => n10137, B1 => 
                           REGISTERS_5_4_port, B2 => n10047, ZN => n10051);
   U2742 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n10131, B1 => 
                           REGISTERS_1_4_port, B2 => n10130, ZN => n10050);
   U2743 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n10177, B1 => 
                           REGISTERS_4_4_port, B2 => n10188, ZN => n10049);
   U2744 : AOI22_X1 port map( A1 => REGISTERS_6_4_port, A2 => n10186, B1 => 
                           REGISTERS_2_4_port, B2 => n10136, ZN => n10048);
   U2745 : NAND4_X1 port map( A1 => n10051, A2 => n10050, A3 => n10049, A4 => 
                           n10048, ZN => n10058);
   U2746 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n10137, B1 => 
                           REGISTERS_12_4_port, B2 => n10188, ZN => n10056);
   U2747 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n10131, B1 => 
                           REGISTERS_13_4_port, B2 => n10129, ZN => n10055);
   U2748 : AOI22_X1 port map( A1 => REGISTERS_9_4_port, A2 => n10189, B1 => 
                           REGISTERS_8_4_port, B2 => n10052, ZN => n10054);
   U2749 : AOI22_X1 port map( A1 => REGISTERS_14_4_port, A2 => n10186, B1 => 
                           REGISTERS_10_4_port, B2 => n10102, ZN => n10053);
   U2750 : NAND4_X1 port map( A1 => n10056, A2 => n10055, A3 => n10054, A4 => 
                           n10053, ZN => n10057);
   U2751 : AOI22_X1 port map( A1 => n10198, A2 => n10058, B1 => n10196, B2 => 
                           n10057, ZN => n10059);
   U2752 : OAI21_X1 port map( B1 => n10201, B2 => n10060, A => n10059, ZN => 
                           N389);
   U2753 : AOI22_X1 port map( A1 => REGISTERS_22_3_port, A2 => n10087, B1 => 
                           REGISTERS_25_3_port, B2 => n10093, ZN => n10065);
   U2754 : AOI22_X1 port map( A1 => REGISTERS_30_3_port, A2 => n10150, B1 => 
                           REGISTERS_31_3_port, B2 => n10061, ZN => n10064);
   U2755 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n10155, B1 => 
                           REGISTERS_29_3_port, B2 => n10149, ZN => n10063);
   U2756 : AOI22_X1 port map( A1 => REGISTERS_18_3_port, A2 => n10154, B1 => 
                           REGISTERS_16_3_port, B2 => n10153, ZN => n10062);
   U2757 : NAND4_X1 port map( A1 => n10065, A2 => n10064, A3 => n10063, A4 => 
                           n10062, ZN => n10073);
   U2758 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n10066, B1 => 
                           REGISTERS_28_3_port, B2 => n10121, ZN => n10071);
   U2759 : AOI22_X1 port map( A1 => REGISTERS_27_3_port, A2 => n10094, B1 => 
                           REGISTERS_21_3_port, B2 => n10161, ZN => n10070);
   U2760 : AOI22_X1 port map( A1 => REGISTERS_17_3_port, A2 => n10088, B1 => 
                           REGISTERS_26_3_port, B2 => n10122, ZN => n10069);
   U2761 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n10067, B1 => 
                           REGISTERS_23_3_port, B2 => n10167, ZN => n10068);
   U2762 : NAND4_X1 port map( A1 => n10071, A2 => n10070, A3 => n10069, A4 => 
                           n10068, ZN => n10072);
   U2763 : NOR2_X1 port map( A1 => n10073, A2 => n10072, ZN => n10086);
   U2764 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n10188, B1 => 
                           REGISTERS_3_3_port, B2 => n10178, ZN => n10077);
   U2765 : AOI22_X1 port map( A1 => REGISTERS_1_3_port, A2 => n10138, B1 => 
                           REGISTERS_7_3_port, B2 => n10131, ZN => n10076);
   U2766 : AOI22_X1 port map( A1 => REGISTERS_2_3_port, A2 => n10184, B1 => 
                           REGISTERS_6_3_port, B2 => n10175, ZN => n10075);
   U2767 : AOI22_X1 port map( A1 => REGISTERS_5_3_port, A2 => n10190, B1 => 
                           REGISTERS_0_3_port, B2 => n10185, ZN => n10074);
   U2768 : NAND4_X1 port map( A1 => n10077, A2 => n10076, A3 => n10075, A4 => 
                           n10074, ZN => n10084);
   U2769 : AOI22_X1 port map( A1 => REGISTERS_9_3_port, A2 => n10130, B1 => 
                           REGISTERS_10_3_port, B2 => n10136, ZN => n10082);
   U2770 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n10177, B1 => 
                           REGISTERS_11_3_port, B2 => n10178, ZN => n10081);
   U2771 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n10139, B1 => 
                           REGISTERS_15_3_port, B2 => n10176, ZN => n10080);
   U2772 : AOI22_X1 port map( A1 => REGISTERS_13_3_port, A2 => n10190, B1 => 
                           REGISTERS_14_3_port, B2 => n10078, ZN => n10079);
   U2773 : NAND4_X1 port map( A1 => n10082, A2 => n10081, A3 => n10080, A4 => 
                           n10079, ZN => n10083);
   U2774 : AOI22_X1 port map( A1 => n10198, A2 => n10084, B1 => n10196, B2 => 
                           n10083, ZN => n10085);
   U2775 : OAI21_X1 port map( B1 => n10148, B2 => n10086, A => n10085, ZN => 
                           N388);
   U2776 : AOI22_X1 port map( A1 => REGISTERS_30_2_port, A2 => n10150, B1 => 
                           REGISTERS_26_2_port, B2 => n10122, ZN => n10092);
   U2777 : AOI22_X1 port map( A1 => REGISTERS_17_2_port, A2 => n10088, B1 => 
                           REGISTERS_22_2_port, B2 => n10087, ZN => n10091);
   U2778 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n10115, B1 => 
                           REGISTERS_18_2_port, B2 => n10154, ZN => n10090);
   U2779 : AOI22_X1 port map( A1 => REGISTERS_21_2_port, A2 => n10161, B1 => 
                           REGISTERS_19_2_port, B2 => n10155, ZN => n10089);
   U2780 : NAND4_X1 port map( A1 => n10092, A2 => n10091, A3 => n10090, A4 => 
                           n10089, ZN => n10100);
   U2781 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n10167, B1 => 
                           REGISTERS_28_2_port, B2 => n10121, ZN => n10098);
   U2782 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n10149, B1 => 
                           REGISTERS_25_2_port, B2 => n10093, ZN => n10097);
   U2783 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n10094, B1 => 
                           REGISTERS_24_2_port, B2 => n10165, ZN => n10096);
   U2784 : AOI22_X1 port map( A1 => REGISTERS_31_2_port, A2 => n10164, B1 => 
                           REGISTERS_20_2_port, B2 => n10162, ZN => n10095);
   U2785 : NAND4_X1 port map( A1 => n10098, A2 => n10097, A3 => n10096, A4 => 
                           n10095, ZN => n10099);
   U2786 : NOR2_X1 port map( A1 => n10100, A2 => n10099, ZN => n10114);
   U2787 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n10137, B1 => 
                           REGISTERS_6_2_port, B2 => n10175, ZN => n10106);
   U2788 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n10101, B1 => 
                           REGISTERS_7_2_port, B2 => n10183, ZN => n10105);
   U2789 : AOI22_X1 port map( A1 => REGISTERS_1_2_port, A2 => n10189, B1 => 
                           REGISTERS_0_2_port, B2 => n10185, ZN => n10104);
   U2790 : AOI22_X1 port map( A1 => REGISTERS_5_2_port, A2 => n10190, B1 => 
                           REGISTERS_2_2_port, B2 => n10102, ZN => n10103);
   U2791 : NAND4_X1 port map( A1 => n10106, A2 => n10105, A3 => n10104, A4 => 
                           n10103, ZN => n10112);
   U2792 : AOI22_X1 port map( A1 => REGISTERS_11_2_port, A2 => n10137, B1 => 
                           REGISTERS_15_2_port, B2 => n10131, ZN => n10110);
   U2793 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n10188, B1 => 
                           REGISTERS_13_2_port, B2 => n10129, ZN => n10109);
   U2794 : AOI22_X1 port map( A1 => REGISTERS_10_2_port, A2 => n10184, B1 => 
                           REGISTERS_14_2_port, B2 => n10175, ZN => n10108);
   U2795 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n10177, B1 => 
                           REGISTERS_9_2_port, B2 => n10130, ZN => n10107);
   U2796 : NAND4_X1 port map( A1 => n10110, A2 => n10109, A3 => n10108, A4 => 
                           n10107, ZN => n10111);
   U2797 : AOI22_X1 port map( A1 => n10198, A2 => n10112, B1 => n10196, B2 => 
                           n10111, ZN => n10113);
   U2798 : OAI21_X1 port map( B1 => n10201, B2 => n10114, A => n10113, ZN => 
                           N387);
   U2799 : AOI22_X1 port map( A1 => REGISTERS_22_1_port, A2 => n10163, B1 => 
                           REGISTERS_20_1_port, B2 => n10162, ZN => n10120);
   U2800 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n10149, B1 => 
                           REGISTERS_19_1_port, B2 => n10155, ZN => n10119);
   U2801 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n10115, B1 => 
                           REGISTERS_27_1_port, B2 => n10168, ZN => n10118);
   U2802 : AOI22_X1 port map( A1 => REGISTERS_21_1_port, A2 => n10161, B1 => 
                           REGISTERS_30_1_port, B2 => n10116, ZN => n10117);
   U2803 : NAND4_X1 port map( A1 => n10120, A2 => n10119, A3 => n10118, A4 => 
                           n10117, ZN => n10128);
   U2804 : AOI22_X1 port map( A1 => REGISTERS_31_1_port, A2 => n10164, B1 => 
                           REGISTERS_23_1_port, B2 => n10167, ZN => n10126);
   U2805 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n10165, B1 => 
                           REGISTERS_17_1_port, B2 => n10156, ZN => n10125);
   U2806 : AOI22_X1 port map( A1 => REGISTERS_25_1_port, A2 => n10151, B1 => 
                           REGISTERS_28_1_port, B2 => n10121, ZN => n10124);
   U2807 : AOI22_X1 port map( A1 => REGISTERS_18_1_port, A2 => n10154, B1 => 
                           REGISTERS_26_1_port, B2 => n10122, ZN => n10123);
   U2808 : NAND4_X1 port map( A1 => n10126, A2 => n10125, A3 => n10124, A4 => 
                           n10123, ZN => n10127);
   U2809 : NOR2_X1 port map( A1 => n10128, A2 => n10127, ZN => n10147);
   U2810 : AOI22_X1 port map( A1 => REGISTERS_1_1_port, A2 => n10130, B1 => 
                           REGISTERS_5_1_port, B2 => n10129, ZN => n10135);
   U2811 : AOI22_X1 port map( A1 => REGISTERS_6_1_port, A2 => n10186, B1 => 
                           REGISTERS_2_1_port, B2 => n10136, ZN => n10134);
   U2812 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n10131, B1 => 
                           REGISTERS_4_1_port, B2 => n10139, ZN => n10133);
   U2813 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n10177, B1 => 
                           REGISTERS_3_1_port, B2 => n10187, ZN => n10132);
   U2814 : NAND4_X1 port map( A1 => n10135, A2 => n10134, A3 => n10133, A4 => 
                           n10132, ZN => n10145);
   U2815 : AOI22_X1 port map( A1 => REGISTERS_14_1_port, A2 => n10186, B1 => 
                           REGISTERS_10_1_port, B2 => n10136, ZN => n10143);
   U2816 : AOI22_X1 port map( A1 => REGISTERS_13_1_port, A2 => n10190, B1 => 
                           REGISTERS_8_1_port, B2 => n10185, ZN => n10142);
   U2817 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n10137, B1 => 
                           REGISTERS_15_1_port, B2 => n10183, ZN => n10141);
   U2818 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n10139, B1 => 
                           REGISTERS_9_1_port, B2 => n10138, ZN => n10140);
   U2819 : NAND4_X1 port map( A1 => n10143, A2 => n10142, A3 => n10141, A4 => 
                           n10140, ZN => n10144);
   U2820 : AOI22_X1 port map( A1 => n10198, A2 => n10145, B1 => n10196, B2 => 
                           n10144, ZN => n10146);
   U2821 : OAI21_X1 port map( B1 => n10148, B2 => n10147, A => n10146, ZN => 
                           N386);
   U2822 : AOI22_X1 port map( A1 => REGISTERS_30_0_port, A2 => n10150, B1 => 
                           REGISTERS_29_0_port, B2 => n10149, ZN => n10160);
   U2823 : AOI22_X1 port map( A1 => REGISTERS_26_0_port, A2 => n10152, B1 => 
                           REGISTERS_25_0_port, B2 => n10151, ZN => n10159);
   U2824 : AOI22_X1 port map( A1 => REGISTERS_18_0_port, A2 => n10154, B1 => 
                           REGISTERS_16_0_port, B2 => n10153, ZN => n10158);
   U2825 : AOI22_X1 port map( A1 => REGISTERS_17_0_port, A2 => n10156, B1 => 
                           REGISTERS_19_0_port, B2 => n10155, ZN => n10157);
   U2826 : NAND4_X1 port map( A1 => n10160, A2 => n10159, A3 => n10158, A4 => 
                           n10157, ZN => n10174);
   U2827 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n10162, B1 => 
                           REGISTERS_21_0_port, B2 => n10161, ZN => n10172);
   U2828 : AOI22_X1 port map( A1 => REGISTERS_31_0_port, A2 => n10164, B1 => 
                           REGISTERS_22_0_port, B2 => n10163, ZN => n10171);
   U2829 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n10166, B1 => 
                           REGISTERS_24_0_port, B2 => n10165, ZN => n10170);
   U2830 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n10168, B1 => 
                           REGISTERS_23_0_port, B2 => n10167, ZN => n10169);
   U2831 : NAND4_X1 port map( A1 => n10172, A2 => n10171, A3 => n10170, A4 => 
                           n10169, ZN => n10173);
   U2832 : NOR2_X1 port map( A1 => n10174, A2 => n10173, ZN => n10200);
   U2833 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n10188, B1 => 
                           REGISTERS_6_0_port, B2 => n10175, ZN => n10182);
   U2834 : AOI22_X1 port map( A1 => REGISTERS_2_0_port, A2 => n10184, B1 => 
                           REGISTERS_7_0_port, B2 => n10176, ZN => n10181);
   U2835 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n10177, B1 => 
                           REGISTERS_1_0_port, B2 => n10189, ZN => n10180);
   U2836 : AOI22_X1 port map( A1 => REGISTERS_5_0_port, A2 => n10190, B1 => 
                           REGISTERS_3_0_port, B2 => n10178, ZN => n10179);
   U2837 : NAND4_X1 port map( A1 => n10182, A2 => n10181, A3 => n10180, A4 => 
                           n10179, ZN => n10197);
   U2838 : AOI22_X1 port map( A1 => REGISTERS_10_0_port, A2 => n10184, B1 => 
                           REGISTERS_15_0_port, B2 => n10183, ZN => n10194);
   U2839 : AOI22_X1 port map( A1 => REGISTERS_14_0_port, A2 => n10186, B1 => 
                           REGISTERS_8_0_port, B2 => n10185, ZN => n10193);
   U2840 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n10188, B1 => 
                           REGISTERS_11_0_port, B2 => n10187, ZN => n10192);
   U2841 : AOI22_X1 port map( A1 => REGISTERS_13_0_port, A2 => n10190, B1 => 
                           REGISTERS_9_0_port, B2 => n10189, ZN => n10191);
   U2842 : NAND4_X1 port map( A1 => n10194, A2 => n10193, A3 => n10192, A4 => 
                           n10191, ZN => n10195);
   U2843 : AOI22_X1 port map( A1 => n10198, A2 => n10197, B1 => n10196, B2 => 
                           n10195, ZN => n10199);
   U2844 : OAI21_X1 port map( B1 => n10201, B2 => n10200, A => n10199, ZN => 
                           N385);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ENABLE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ENABLE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component general_alu_N32
      port( clk : in std_logic;  zero_mul_detect, mul_exeception : out 
            std_logic;  FUNC : in std_logic_vector (0 to 3);  DATA1, DATA2 : in
            std_logic_vector (31 downto 0);  cin, signed_notsigned : in 
            std_logic;  overflow : out std_logic;  OUTALU : out 
            std_logic_vector (31 downto 0);  rst_BAR : in std_logic);
   end component;
   
   component register_file_NBITREG32_NBITADD5
      port( CLK, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2
            : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector 
            (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0);  
            RESET_BAR : in std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ENABLE_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, curr_instruction_to_cu_i_31_port, 
      curr_instruction_to_cu_i_30_port, curr_instruction_to_cu_i_28_port, 
      curr_instruction_to_cu_i_27_port, curr_instruction_to_cu_i_26_port, 
      curr_instruction_to_cu_i_20_port, curr_instruction_to_cu_i_19_port, 
      curr_instruction_to_cu_i_18_port, curr_instruction_to_cu_i_17_port, 
      curr_instruction_to_cu_i_16_port, curr_instruction_to_cu_i_15_port, 
      curr_instruction_to_cu_i_14_port, curr_instruction_to_cu_i_13_port, 
      curr_instruction_to_cu_i_12_port, curr_instruction_to_cu_i_11_port, 
      curr_instruction_to_cu_i_5_port, curr_instruction_to_cu_i_4_port, 
      curr_instruction_to_cu_i_3_port, curr_instruction_to_cu_i_2_port, 
      curr_instruction_to_cu_i_1_port, curr_instruction_to_cu_i_0_port, 
      enable_rf_i, read_rf_p2_i, alu_cin_i, write_rf_i, cu_i_n131, cu_i_n127, 
      cu_i_n126, cu_i_n125, cu_i_n124, cu_i_n123, cu_i_n210, cu_i_n209, 
      cu_i_n145, cu_i_n26, cu_i_n25, cu_i_n23, cu_i_cw1_i_4_port, 
      cu_i_cw1_i_7_port, cu_i_cw1_i_8_port, cu_i_cw3_6_port, cu_i_cw2_5_port, 
      cu_i_cw2_6_port, cu_i_cw2_7_port, cu_i_cw2_8_port, cu_i_cw1_0_port, 
      cu_i_cw1_1_port, cu_i_cw1_2_port, cu_i_cw1_3_port, cu_i_cw1_4_port, 
      cu_i_cw1_5_port, cu_i_cw1_6_port, cu_i_cw1_7_port, cu_i_cw1_8_port, 
      cu_i_cw1_10_port, cu_i_cw1_11_port, cu_i_cw1_12_port, cu_i_N279, 
      cu_i_N278, cu_i_N277, cu_i_N276, cu_i_N275, cu_i_N274, cu_i_N273, 
      cu_i_N267, cu_i_N266, cu_i_N265, cu_i_N264, cu_i_cmd_alu_op_type_0_port, 
      cu_i_cmd_alu_op_type_1_port, cu_i_cmd_alu_op_type_2_port, 
      cu_i_cmd_alu_op_type_3_port, cu_i_cmd_word_1_port, cu_i_cmd_word_3_port, 
      cu_i_cmd_word_4_port, cu_i_cmd_word_6_port, cu_i_cmd_word_7_port, 
      cu_i_cmd_word_8_port, cu_i_next_stall, cu_i_next_val_counter_mul_0_port, 
      cu_i_next_val_counter_mul_1_port, cu_i_next_val_counter_mul_2_port, 
      cu_i_next_val_counter_mul_3_port, datapath_i_data_from_alu_i_0_port, 
      datapath_i_data_from_alu_i_1_port, datapath_i_data_from_alu_i_2_port, 
      datapath_i_data_from_alu_i_3_port, datapath_i_data_from_alu_i_4_port, 
      datapath_i_data_from_alu_i_5_port, datapath_i_data_from_alu_i_6_port, 
      datapath_i_data_from_alu_i_7_port, datapath_i_data_from_alu_i_8_port, 
      datapath_i_data_from_alu_i_9_port, datapath_i_data_from_alu_i_10_port, 
      datapath_i_data_from_alu_i_11_port, datapath_i_data_from_alu_i_12_port, 
      datapath_i_data_from_alu_i_13_port, datapath_i_data_from_alu_i_14_port, 
      datapath_i_data_from_alu_i_15_port, datapath_i_data_from_alu_i_16_port, 
      datapath_i_data_from_alu_i_17_port, datapath_i_data_from_alu_i_18_port, 
      datapath_i_data_from_alu_i_19_port, datapath_i_data_from_alu_i_20_port, 
      datapath_i_data_from_alu_i_21_port, datapath_i_data_from_alu_i_22_port, 
      datapath_i_data_from_alu_i_23_port, datapath_i_data_from_alu_i_24_port, 
      datapath_i_data_from_alu_i_25_port, datapath_i_data_from_alu_i_26_port, 
      datapath_i_data_from_alu_i_27_port, datapath_i_data_from_alu_i_28_port, 
      datapath_i_data_from_alu_i_29_port, datapath_i_data_from_alu_i_30_port, 
      datapath_i_data_from_alu_i_31_port, datapath_i_data_from_memory_i_0_port,
      datapath_i_data_from_memory_i_1_port, 
      datapath_i_data_from_memory_i_2_port, 
      datapath_i_data_from_memory_i_3_port, 
      datapath_i_data_from_memory_i_4_port, 
      datapath_i_data_from_memory_i_5_port, 
      datapath_i_data_from_memory_i_6_port, 
      datapath_i_data_from_memory_i_7_port, 
      datapath_i_data_from_memory_i_8_port, 
      datapath_i_data_from_memory_i_9_port, 
      datapath_i_data_from_memory_i_10_port, 
      datapath_i_data_from_memory_i_11_port, 
      datapath_i_data_from_memory_i_12_port, 
      datapath_i_data_from_memory_i_13_port, 
      datapath_i_data_from_memory_i_14_port, 
      datapath_i_data_from_memory_i_15_port, 
      datapath_i_data_from_memory_i_16_port, 
      datapath_i_data_from_memory_i_17_port, 
      datapath_i_data_from_memory_i_18_port, 
      datapath_i_data_from_memory_i_19_port, 
      datapath_i_data_from_memory_i_20_port, 
      datapath_i_data_from_memory_i_21_port, 
      datapath_i_data_from_memory_i_22_port, 
      datapath_i_data_from_memory_i_23_port, 
      datapath_i_data_from_memory_i_24_port, 
      datapath_i_data_from_memory_i_25_port, 
      datapath_i_data_from_memory_i_26_port, 
      datapath_i_data_from_memory_i_27_port, 
      datapath_i_data_from_memory_i_28_port, 
      datapath_i_data_from_memory_i_29_port, 
      datapath_i_data_from_memory_i_30_port, 
      datapath_i_data_from_memory_i_31_port, datapath_i_value_to_mem_i_0_port, 
      datapath_i_value_to_mem_i_1_port, datapath_i_value_to_mem_i_2_port, 
      datapath_i_value_to_mem_i_3_port, datapath_i_value_to_mem_i_4_port, 
      datapath_i_value_to_mem_i_5_port, datapath_i_value_to_mem_i_6_port, 
      datapath_i_value_to_mem_i_7_port, datapath_i_value_to_mem_i_8_port, 
      datapath_i_value_to_mem_i_9_port, datapath_i_value_to_mem_i_10_port, 
      datapath_i_value_to_mem_i_11_port, datapath_i_value_to_mem_i_12_port, 
      datapath_i_value_to_mem_i_13_port, datapath_i_value_to_mem_i_14_port, 
      datapath_i_value_to_mem_i_15_port, datapath_i_value_to_mem_i_16_port, 
      datapath_i_value_to_mem_i_17_port, datapath_i_value_to_mem_i_18_port, 
      datapath_i_value_to_mem_i_19_port, datapath_i_value_to_mem_i_20_port, 
      datapath_i_value_to_mem_i_21_port, datapath_i_value_to_mem_i_22_port, 
      datapath_i_value_to_mem_i_23_port, datapath_i_value_to_mem_i_24_port, 
      datapath_i_value_to_mem_i_25_port, datapath_i_value_to_mem_i_26_port, 
      datapath_i_value_to_mem_i_27_port, datapath_i_value_to_mem_i_28_port, 
      datapath_i_value_to_mem_i_29_port, datapath_i_value_to_mem_i_30_port, 
      datapath_i_value_to_mem_i_31_port, datapath_i_alu_output_val_i_0_port, 
      datapath_i_alu_output_val_i_1_port, datapath_i_alu_output_val_i_2_port, 
      datapath_i_alu_output_val_i_3_port, datapath_i_alu_output_val_i_4_port, 
      datapath_i_alu_output_val_i_5_port, datapath_i_alu_output_val_i_6_port, 
      datapath_i_alu_output_val_i_7_port, datapath_i_alu_output_val_i_8_port, 
      datapath_i_alu_output_val_i_9_port, datapath_i_alu_output_val_i_10_port, 
      datapath_i_alu_output_val_i_11_port, datapath_i_alu_output_val_i_12_port,
      datapath_i_alu_output_val_i_13_port, datapath_i_alu_output_val_i_14_port,
      datapath_i_alu_output_val_i_15_port, datapath_i_alu_output_val_i_16_port,
      datapath_i_alu_output_val_i_17_port, datapath_i_alu_output_val_i_18_port,
      datapath_i_alu_output_val_i_19_port, datapath_i_alu_output_val_i_20_port,
      datapath_i_alu_output_val_i_21_port, datapath_i_alu_output_val_i_22_port,
      datapath_i_alu_output_val_i_23_port, datapath_i_alu_output_val_i_24_port,
      datapath_i_alu_output_val_i_25_port, datapath_i_alu_output_val_i_26_port,
      datapath_i_alu_output_val_i_27_port, datapath_i_alu_output_val_i_28_port,
      datapath_i_alu_output_val_i_29_port, datapath_i_alu_output_val_i_30_port,
      datapath_i_alu_output_val_i_31_port, datapath_i_val_immediate_i_0_port, 
      datapath_i_val_immediate_i_1_port, datapath_i_val_immediate_i_2_port, 
      datapath_i_val_immediate_i_3_port, datapath_i_val_immediate_i_4_port, 
      datapath_i_val_immediate_i_5_port, datapath_i_val_immediate_i_6_port, 
      datapath_i_val_immediate_i_7_port, datapath_i_val_immediate_i_8_port, 
      datapath_i_val_immediate_i_9_port, datapath_i_val_immediate_i_10_port, 
      datapath_i_val_immediate_i_11_port, datapath_i_val_immediate_i_12_port, 
      datapath_i_val_immediate_i_13_port, datapath_i_val_immediate_i_14_port, 
      datapath_i_val_immediate_i_15_port, datapath_i_val_immediate_i_16_port, 
      datapath_i_val_immediate_i_17_port, datapath_i_val_immediate_i_18_port, 
      datapath_i_val_immediate_i_19_port, datapath_i_val_immediate_i_20_port, 
      datapath_i_val_immediate_i_21_port, datapath_i_val_immediate_i_22_port, 
      datapath_i_val_immediate_i_23_port, datapath_i_val_immediate_i_24_port, 
      datapath_i_val_immediate_i_25_port, datapath_i_val_b_i_0_port, 
      datapath_i_val_b_i_1_port, datapath_i_val_b_i_2_port, 
      datapath_i_val_b_i_3_port, datapath_i_val_b_i_4_port, 
      datapath_i_val_b_i_5_port, datapath_i_val_b_i_6_port, 
      datapath_i_val_b_i_7_port, datapath_i_val_b_i_8_port, 
      datapath_i_val_b_i_9_port, datapath_i_val_b_i_10_port, 
      datapath_i_val_b_i_11_port, datapath_i_val_b_i_12_port, 
      datapath_i_val_b_i_13_port, datapath_i_val_b_i_14_port, 
      datapath_i_val_b_i_15_port, datapath_i_val_b_i_16_port, 
      datapath_i_val_b_i_17_port, datapath_i_val_b_i_18_port, 
      datapath_i_val_b_i_19_port, datapath_i_val_b_i_20_port, 
      datapath_i_val_b_i_21_port, datapath_i_val_b_i_22_port, 
      datapath_i_val_b_i_23_port, datapath_i_val_b_i_24_port, 
      datapath_i_val_b_i_25_port, datapath_i_val_b_i_26_port, 
      datapath_i_val_b_i_27_port, datapath_i_val_b_i_28_port, 
      datapath_i_val_b_i_29_port, datapath_i_val_b_i_30_port, 
      datapath_i_val_b_i_31_port, datapath_i_val_a_i_0_port, 
      datapath_i_val_a_i_1_port, datapath_i_val_a_i_2_port, 
      datapath_i_val_a_i_3_port, datapath_i_val_a_i_4_port, 
      datapath_i_val_a_i_5_port, datapath_i_val_a_i_6_port, 
      datapath_i_val_a_i_7_port, datapath_i_val_a_i_8_port, 
      datapath_i_val_a_i_9_port, datapath_i_val_a_i_10_port, 
      datapath_i_val_a_i_11_port, datapath_i_val_a_i_12_port, 
      datapath_i_val_a_i_13_port, datapath_i_val_a_i_14_port, 
      datapath_i_val_a_i_15_port, datapath_i_val_a_i_16_port, 
      datapath_i_val_a_i_17_port, datapath_i_val_a_i_18_port, 
      datapath_i_val_a_i_19_port, datapath_i_val_a_i_20_port, 
      datapath_i_val_a_i_21_port, datapath_i_val_a_i_22_port, 
      datapath_i_val_a_i_23_port, datapath_i_val_a_i_24_port, 
      datapath_i_val_a_i_25_port, datapath_i_val_a_i_26_port, 
      datapath_i_val_a_i_27_port, datapath_i_val_a_i_28_port, 
      datapath_i_val_a_i_29_port, datapath_i_val_a_i_30_port, 
      datapath_i_val_a_i_31_port, datapath_i_new_pc_value_decode_0_port, 
      datapath_i_new_pc_value_decode_1_port, 
      datapath_i_new_pc_value_decode_2_port, 
      datapath_i_new_pc_value_decode_3_port, 
      datapath_i_new_pc_value_decode_4_port, 
      datapath_i_new_pc_value_decode_5_port, 
      datapath_i_new_pc_value_decode_6_port, 
      datapath_i_new_pc_value_decode_7_port, 
      datapath_i_new_pc_value_decode_8_port, 
      datapath_i_new_pc_value_decode_9_port, 
      datapath_i_new_pc_value_decode_10_port, 
      datapath_i_new_pc_value_decode_11_port, 
      datapath_i_new_pc_value_decode_12_port, 
      datapath_i_new_pc_value_decode_13_port, 
      datapath_i_new_pc_value_decode_14_port, 
      datapath_i_new_pc_value_decode_15_port, 
      datapath_i_new_pc_value_decode_16_port, 
      datapath_i_new_pc_value_decode_17_port, 
      datapath_i_new_pc_value_decode_18_port, 
      datapath_i_new_pc_value_decode_19_port, 
      datapath_i_new_pc_value_decode_20_port, 
      datapath_i_new_pc_value_decode_21_port, 
      datapath_i_new_pc_value_decode_22_port, 
      datapath_i_new_pc_value_decode_23_port, 
      datapath_i_new_pc_value_decode_24_port, 
      datapath_i_new_pc_value_decode_25_port, 
      datapath_i_new_pc_value_decode_26_port, 
      datapath_i_new_pc_value_decode_27_port, 
      datapath_i_new_pc_value_decode_28_port, 
      datapath_i_new_pc_value_decode_29_port, 
      datapath_i_new_pc_value_decode_30_port, 
      datapath_i_new_pc_value_decode_31_port, 
      datapath_i_new_pc_value_mem_stage_i_2_port, 
      datapath_i_new_pc_value_mem_stage_i_3_port, 
      datapath_i_new_pc_value_mem_stage_i_4_port, 
      datapath_i_new_pc_value_mem_stage_i_5_port, 
      datapath_i_new_pc_value_mem_stage_i_6_port, 
      datapath_i_new_pc_value_mem_stage_i_7_port, 
      datapath_i_new_pc_value_mem_stage_i_8_port, 
      datapath_i_new_pc_value_mem_stage_i_9_port, 
      datapath_i_new_pc_value_mem_stage_i_10_port, 
      datapath_i_new_pc_value_mem_stage_i_11_port, 
      datapath_i_new_pc_value_mem_stage_i_12_port, 
      datapath_i_new_pc_value_mem_stage_i_13_port, 
      datapath_i_new_pc_value_mem_stage_i_14_port, 
      datapath_i_new_pc_value_mem_stage_i_15_port, 
      datapath_i_new_pc_value_mem_stage_i_16_port, 
      datapath_i_new_pc_value_mem_stage_i_17_port, 
      datapath_i_new_pc_value_mem_stage_i_18_port, 
      datapath_i_new_pc_value_mem_stage_i_19_port, 
      datapath_i_new_pc_value_mem_stage_i_20_port, 
      datapath_i_new_pc_value_mem_stage_i_21_port, 
      datapath_i_new_pc_value_mem_stage_i_22_port, 
      datapath_i_new_pc_value_mem_stage_i_23_port, 
      datapath_i_new_pc_value_mem_stage_i_24_port, 
      datapath_i_new_pc_value_mem_stage_i_25_port, 
      datapath_i_new_pc_value_mem_stage_i_26_port, 
      datapath_i_new_pc_value_mem_stage_i_27_port, 
      datapath_i_new_pc_value_mem_stage_i_28_port, 
      datapath_i_new_pc_value_mem_stage_i_29_port, 
      datapath_i_new_pc_value_mem_stage_i_30_port, 
      datapath_i_new_pc_value_mem_stage_i_31_port, datapath_i_n18, 
      datapath_i_n17, datapath_i_n16, datapath_i_n15, datapath_i_n14, 
      datapath_i_n13, datapath_i_n12, datapath_i_n11, datapath_i_n10, 
      datapath_i_n9, datapath_i_fetch_stage_dp_n69, 
      datapath_i_fetch_stage_dp_n68, datapath_i_fetch_stage_dp_n67, 
      datapath_i_fetch_stage_dp_n66, datapath_i_fetch_stage_dp_n65, 
      datapath_i_fetch_stage_dp_n64, datapath_i_fetch_stage_dp_n63, 
      datapath_i_fetch_stage_dp_n62, datapath_i_fetch_stage_dp_n61, 
      datapath_i_fetch_stage_dp_n60, datapath_i_fetch_stage_dp_n59, 
      datapath_i_fetch_stage_dp_n58, datapath_i_fetch_stage_dp_n57, 
      datapath_i_fetch_stage_dp_n56, datapath_i_fetch_stage_dp_n55, 
      datapath_i_fetch_stage_dp_n54, datapath_i_fetch_stage_dp_n53, 
      datapath_i_fetch_stage_dp_n52, datapath_i_fetch_stage_dp_n51, 
      datapath_i_fetch_stage_dp_n50, datapath_i_fetch_stage_dp_n49, 
      datapath_i_fetch_stage_dp_n48, datapath_i_fetch_stage_dp_n47, 
      datapath_i_fetch_stage_dp_n46, datapath_i_fetch_stage_dp_n45, 
      datapath_i_fetch_stage_dp_n44, datapath_i_fetch_stage_dp_n43, 
      datapath_i_fetch_stage_dp_n42, datapath_i_fetch_stage_dp_n41, 
      datapath_i_fetch_stage_dp_n40, datapath_i_fetch_stage_dp_n39, 
      datapath_i_fetch_stage_dp_n38, datapath_i_fetch_stage_dp_n37, 
      datapath_i_fetch_stage_dp_n36, datapath_i_fetch_stage_dp_n35, 
      datapath_i_fetch_stage_dp_n34, datapath_i_fetch_stage_dp_n33, 
      datapath_i_fetch_stage_dp_n32, datapath_i_fetch_stage_dp_n31, 
      datapath_i_fetch_stage_dp_n30, datapath_i_fetch_stage_dp_n29, 
      datapath_i_fetch_stage_dp_n28, datapath_i_fetch_stage_dp_n27, 
      datapath_i_fetch_stage_dp_n26, datapath_i_fetch_stage_dp_n25, 
      datapath_i_fetch_stage_dp_n24, datapath_i_fetch_stage_dp_n23, 
      datapath_i_fetch_stage_dp_n22, datapath_i_fetch_stage_dp_n21, 
      datapath_i_fetch_stage_dp_n20, datapath_i_fetch_stage_dp_n19, 
      datapath_i_fetch_stage_dp_n18, datapath_i_fetch_stage_dp_n17, 
      datapath_i_fetch_stage_dp_n16, datapath_i_fetch_stage_dp_n15, 
      datapath_i_fetch_stage_dp_n14, datapath_i_fetch_stage_dp_n13, 
      datapath_i_fetch_stage_dp_n12, datapath_i_fetch_stage_dp_n11, 
      datapath_i_fetch_stage_dp_n10, datapath_i_fetch_stage_dp_n9, 
      datapath_i_fetch_stage_dp_n4, datapath_i_fetch_stage_dp_n3, 
      datapath_i_fetch_stage_dp_n2, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port, datapath_i_fetch_stage_dp_N6, 
      datapath_i_fetch_stage_dp_N5, datapath_i_decode_stage_dp_n78, 
      datapath_i_decode_stage_dp_n43, datapath_i_decode_stage_dp_n42, 
      datapath_i_decode_stage_dp_n41, datapath_i_decode_stage_dp_n40, 
      datapath_i_decode_stage_dp_n39, datapath_i_decode_stage_dp_n38, 
      datapath_i_decode_stage_dp_n37, datapath_i_decode_stage_dp_n36, 
      datapath_i_decode_stage_dp_n35, datapath_i_decode_stage_dp_n34, 
      datapath_i_decode_stage_dp_n33, datapath_i_decode_stage_dp_n32, 
      datapath_i_decode_stage_dp_n31, datapath_i_decode_stage_dp_n30, 
      datapath_i_decode_stage_dp_n29, datapath_i_decode_stage_dp_n28, 
      datapath_i_decode_stage_dp_n27, datapath_i_decode_stage_dp_n26, 
      datapath_i_decode_stage_dp_n25, datapath_i_decode_stage_dp_n24, 
      datapath_i_decode_stage_dp_n23, datapath_i_decode_stage_dp_n22, 
      datapath_i_decode_stage_dp_n21, datapath_i_decode_stage_dp_n20, 
      datapath_i_decode_stage_dp_n19, datapath_i_decode_stage_dp_n18, 
      datapath_i_decode_stage_dp_n17, datapath_i_decode_stage_dp_n16, 
      datapath_i_decode_stage_dp_n15, datapath_i_decode_stage_dp_n14, 
      datapath_i_decode_stage_dp_n13, datapath_i_decode_stage_dp_n12, 
      datapath_i_decode_stage_dp_pc_delay3_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_0_port, 
      datapath_i_decode_stage_dp_pc_delay2_1_port, 
      datapath_i_decode_stage_dp_pc_delay2_2_port, 
      datapath_i_decode_stage_dp_pc_delay2_3_port, 
      datapath_i_decode_stage_dp_pc_delay2_4_port, 
      datapath_i_decode_stage_dp_pc_delay2_5_port, 
      datapath_i_decode_stage_dp_pc_delay2_6_port, 
      datapath_i_decode_stage_dp_pc_delay2_7_port, 
      datapath_i_decode_stage_dp_pc_delay2_8_port, 
      datapath_i_decode_stage_dp_pc_delay2_9_port, 
      datapath_i_decode_stage_dp_pc_delay2_10_port, 
      datapath_i_decode_stage_dp_pc_delay2_11_port, 
      datapath_i_decode_stage_dp_pc_delay2_12_port, 
      datapath_i_decode_stage_dp_pc_delay2_13_port, 
      datapath_i_decode_stage_dp_pc_delay2_14_port, 
      datapath_i_decode_stage_dp_pc_delay2_15_port, 
      datapath_i_decode_stage_dp_pc_delay2_16_port, 
      datapath_i_decode_stage_dp_pc_delay2_17_port, 
      datapath_i_decode_stage_dp_pc_delay2_18_port, 
      datapath_i_decode_stage_dp_pc_delay2_19_port, 
      datapath_i_decode_stage_dp_pc_delay2_20_port, 
      datapath_i_decode_stage_dp_pc_delay2_21_port, 
      datapath_i_decode_stage_dp_pc_delay2_22_port, 
      datapath_i_decode_stage_dp_pc_delay2_23_port, 
      datapath_i_decode_stage_dp_pc_delay2_24_port, 
      datapath_i_decode_stage_dp_pc_delay2_25_port, 
      datapath_i_decode_stage_dp_pc_delay2_26_port, 
      datapath_i_decode_stage_dp_pc_delay2_27_port, 
      datapath_i_decode_stage_dp_pc_delay2_28_port, 
      datapath_i_decode_stage_dp_pc_delay2_29_port, 
      datapath_i_decode_stage_dp_pc_delay2_30_port, 
      datapath_i_decode_stage_dp_pc_delay2_31_port, 
      datapath_i_decode_stage_dp_pc_delay2_32_port, 
      datapath_i_decode_stage_dp_clk_immediate, 
      datapath_i_decode_stage_dp_val_reg_immediate_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_31_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
      datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
      datapath_i_decode_stage_dp_enable_rf_i, 
      datapath_i_decode_stage_dp_address_rf_write_0_port, 
      datapath_i_decode_stage_dp_address_rf_write_1_port, 
      datapath_i_decode_stage_dp_address_rf_write_2_port, 
      datapath_i_decode_stage_dp_address_rf_write_3_port, 
      datapath_i_decode_stage_dp_address_rf_write_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
      datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
      datapath_i_execute_stage_dp_n9, datapath_i_execute_stage_dp_n7, 
      datapath_i_execute_stage_dp_alu_out_0_port, 
      datapath_i_execute_stage_dp_alu_out_1_port, 
      datapath_i_execute_stage_dp_alu_out_2_port, 
      datapath_i_execute_stage_dp_alu_out_3_port, 
      datapath_i_execute_stage_dp_alu_out_4_port, 
      datapath_i_execute_stage_dp_alu_out_5_port, 
      datapath_i_execute_stage_dp_alu_out_6_port, 
      datapath_i_execute_stage_dp_alu_out_7_port, 
      datapath_i_execute_stage_dp_alu_out_8_port, 
      datapath_i_execute_stage_dp_alu_out_9_port, 
      datapath_i_execute_stage_dp_alu_out_10_port, 
      datapath_i_execute_stage_dp_alu_out_11_port, 
      datapath_i_execute_stage_dp_alu_out_12_port, 
      datapath_i_execute_stage_dp_alu_out_13_port, 
      datapath_i_execute_stage_dp_alu_out_14_port, 
      datapath_i_execute_stage_dp_alu_out_15_port, 
      datapath_i_execute_stage_dp_alu_out_16_port, 
      datapath_i_execute_stage_dp_alu_out_17_port, 
      datapath_i_execute_stage_dp_alu_out_18_port, 
      datapath_i_execute_stage_dp_alu_out_19_port, 
      datapath_i_execute_stage_dp_alu_out_20_port, 
      datapath_i_execute_stage_dp_alu_out_21_port, 
      datapath_i_execute_stage_dp_alu_out_22_port, 
      datapath_i_execute_stage_dp_alu_out_23_port, 
      datapath_i_execute_stage_dp_alu_out_24_port, 
      datapath_i_execute_stage_dp_alu_out_25_port, 
      datapath_i_execute_stage_dp_alu_out_26_port, 
      datapath_i_execute_stage_dp_alu_out_27_port, 
      datapath_i_execute_stage_dp_alu_out_28_port, 
      datapath_i_execute_stage_dp_alu_out_29_port, 
      datapath_i_execute_stage_dp_alu_out_30_port, 
      datapath_i_execute_stage_dp_alu_out_31_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
      datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
      datapath_i_execute_stage_dp_opb_0_port, 
      datapath_i_execute_stage_dp_opb_1_port, 
      datapath_i_execute_stage_dp_opb_2_port, 
      datapath_i_execute_stage_dp_opb_3_port, 
      datapath_i_execute_stage_dp_opb_4_port, 
      datapath_i_execute_stage_dp_opb_5_port, 
      datapath_i_execute_stage_dp_opb_6_port, 
      datapath_i_execute_stage_dp_opb_7_port, 
      datapath_i_execute_stage_dp_opb_8_port, 
      datapath_i_execute_stage_dp_opb_9_port, 
      datapath_i_execute_stage_dp_opb_10_port, 
      datapath_i_execute_stage_dp_opb_11_port, 
      datapath_i_execute_stage_dp_opb_12_port, 
      datapath_i_execute_stage_dp_opb_13_port, 
      datapath_i_execute_stage_dp_opb_14_port, 
      datapath_i_execute_stage_dp_opb_15_port, 
      datapath_i_execute_stage_dp_opb_16_port, 
      datapath_i_execute_stage_dp_opb_17_port, 
      datapath_i_execute_stage_dp_opb_18_port, 
      datapath_i_execute_stage_dp_opb_19_port, 
      datapath_i_execute_stage_dp_opb_20_port, 
      datapath_i_execute_stage_dp_opb_21_port, 
      datapath_i_execute_stage_dp_opb_22_port, 
      datapath_i_execute_stage_dp_opb_23_port, 
      datapath_i_execute_stage_dp_opb_24_port, 
      datapath_i_execute_stage_dp_opb_25_port, 
      datapath_i_execute_stage_dp_opb_26_port, 
      datapath_i_execute_stage_dp_opb_27_port, 
      datapath_i_execute_stage_dp_opb_28_port, 
      datapath_i_execute_stage_dp_opb_29_port, 
      datapath_i_execute_stage_dp_opb_30_port, 
      datapath_i_execute_stage_dp_opb_31_port, 
      datapath_i_execute_stage_dp_opa_0_port, 
      datapath_i_execute_stage_dp_opa_1_port, 
      datapath_i_execute_stage_dp_opa_2_port, 
      datapath_i_execute_stage_dp_opa_3_port, 
      datapath_i_execute_stage_dp_opa_4_port, 
      datapath_i_execute_stage_dp_opa_5_port, 
      datapath_i_execute_stage_dp_opa_6_port, 
      datapath_i_execute_stage_dp_opa_7_port, 
      datapath_i_execute_stage_dp_opa_8_port, 
      datapath_i_execute_stage_dp_opa_9_port, 
      datapath_i_execute_stage_dp_opa_10_port, 
      datapath_i_execute_stage_dp_opa_11_port, 
      datapath_i_execute_stage_dp_opa_12_port, 
      datapath_i_execute_stage_dp_opa_13_port, 
      datapath_i_execute_stage_dp_opa_14_port, 
      datapath_i_execute_stage_dp_opa_15_port, 
      datapath_i_execute_stage_dp_opa_16_port, 
      datapath_i_execute_stage_dp_opa_17_port, 
      datapath_i_execute_stage_dp_opa_18_port, 
      datapath_i_execute_stage_dp_opa_19_port, 
      datapath_i_execute_stage_dp_opa_20_port, 
      datapath_i_execute_stage_dp_opa_21_port, 
      datapath_i_execute_stage_dp_opa_22_port, 
      datapath_i_execute_stage_dp_opa_23_port, 
      datapath_i_execute_stage_dp_opa_24_port, 
      datapath_i_execute_stage_dp_opa_25_port, 
      datapath_i_execute_stage_dp_opa_26_port, 
      datapath_i_execute_stage_dp_opa_27_port, 
      datapath_i_execute_stage_dp_opa_28_port, 
      datapath_i_execute_stage_dp_opa_29_port, 
      datapath_i_execute_stage_dp_opa_30_port, 
      datapath_i_execute_stage_dp_opa_31_port, 
      datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
      datapath_i_memory_stage_dp_n2, datapath_i_memory_stage_dp_data_ir_0_port,
      datapath_i_memory_stage_dp_data_ir_1_port, 
      datapath_i_memory_stage_dp_data_ir_2_port, 
      datapath_i_memory_stage_dp_data_ir_3_port, 
      datapath_i_memory_stage_dp_data_ir_4_port, 
      datapath_i_memory_stage_dp_data_ir_5_port, 
      datapath_i_memory_stage_dp_data_ir_6_port, 
      datapath_i_memory_stage_dp_data_ir_7_port, 
      datapath_i_memory_stage_dp_data_ir_8_port, 
      datapath_i_memory_stage_dp_data_ir_9_port, 
      datapath_i_memory_stage_dp_data_ir_10_port, 
      datapath_i_memory_stage_dp_data_ir_11_port, 
      datapath_i_memory_stage_dp_data_ir_12_port, 
      datapath_i_memory_stage_dp_data_ir_13_port, 
      datapath_i_memory_stage_dp_data_ir_14_port, 
      datapath_i_memory_stage_dp_data_ir_15_port, 
      datapath_i_memory_stage_dp_data_ir_16_port, 
      datapath_i_memory_stage_dp_data_ir_17_port, 
      datapath_i_memory_stage_dp_data_ir_18_port, 
      datapath_i_memory_stage_dp_data_ir_19_port, 
      datapath_i_memory_stage_dp_data_ir_20_port, 
      datapath_i_memory_stage_dp_data_ir_21_port, 
      datapath_i_memory_stage_dp_data_ir_22_port, 
      datapath_i_memory_stage_dp_data_ir_23_port, 
      datapath_i_memory_stage_dp_data_ir_24_port, 
      datapath_i_memory_stage_dp_data_ir_25_port, 
      datapath_i_memory_stage_dp_data_ir_26_port, 
      datapath_i_memory_stage_dp_data_ir_27_port, 
      datapath_i_memory_stage_dp_data_ir_28_port, 
      datapath_i_memory_stage_dp_data_ir_29_port, 
      datapath_i_memory_stage_dp_data_ir_30_port, 
      datapath_i_memory_stage_dp_data_ir_31_port, n309, n310, n311, n691, n697,
      n699, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n737, n740, n741, 
      n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, 
      n756, n758, n759, n760, n761, n762, n763, n764, n1152, n1534, n1925, 
      n1926, n1927, n1928, n1929, n1932, n1933, n1934, n1935, n1936, n1937, 
      n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, 
      n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, 
      n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, 
      n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, 
      n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, 
      n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, 
      n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, 
      n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, 
      n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
      n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, 
      n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, 
      n2318, n2319, n2320, n2321, DRAM_ENABLE_port, n2323, n2324, n_1413, 
      n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, 
      n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, 
      n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, 
      n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, 
      n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, 
      n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, 
      n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, 
      n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, 
      n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, 
      n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, 
      n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, 
      n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, 
      n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, 
      n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, 
      n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, 
      n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, 
      n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, 
      n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, 
      n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, 
      n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, 
      n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, 
      n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, 
      n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, 
      n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, 
      n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, 
      n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, 
      n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, 
      n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, 
      n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, 
      n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, 
      n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, 
      n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, 
      n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, 
      n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, 
      n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, 
      n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, 
      n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, 
      n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, 
      n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, 
      n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, 
      n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, 
      n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, 
      n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, datapath_i_fetch_stage_dp_N40_port, 
      datapath_i_fetch_stage_dp_N39_port );
   IRAM_ENABLE <= IRAM_ENABLE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, datapath_i_execute_stage_dp_n9, 
      datapath_i_execute_stage_dp_n9 );
   DRAM_ENABLE <= DRAM_ENABLE_port;
   
   cu_i_cmd_alu_op_type_reg_3_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N267, Q => cu_i_cmd_alu_op_type_3_port);
   cu_i_next_val_counter_mul_reg_1_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N275, Q => cu_i_next_val_counter_mul_1_port);
   cu_i_next_val_counter_mul_reg_2_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N276, Q => cu_i_next_val_counter_mul_2_port);
   cu_i_counter_mul_reg_3_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_3_port, CK => CLK, RN => 
                           RST, Q => n2313, QN => cu_i_n124);
   cu_i_next_val_counter_mul_reg_3_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N277, Q => cu_i_next_val_counter_mul_3_port);
   cu_i_counter_mul_reg_0_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_0_port, CK => CLK, RN => 
                           RST, Q => n2303, QN => cu_i_n125);
   cu_i_next_val_counter_mul_reg_0_inst : DLH_X1 port map( G => cu_i_N274, D =>
                           cu_i_N273, Q => cu_i_next_val_counter_mul_0_port);
   cu_i_next_stall_reg : DLH_X1 port map( G => cu_i_N279, D => cu_i_n145, Q => 
                           cu_i_next_stall);
   cu_i_curr_state_reg_1_inst : DFFR_X1 port map( D => cu_i_n209, CK => CLK, RN
                           => RST, Q => n_1413, QN => cu_i_n123);
   datapath_i_decode_stage_dp_reg_file : register_file_NBITREG32_NBITADD5 port 
                           map( CLK => CLK, ENABLE => 
                           datapath_i_decode_stage_dp_enable_rf_i, RD1 => 
                           enable_rf_i, RD2 => read_rf_p2_i, WR => write_rf_i, 
                           ADD_WR(4) => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           ADD_WR(3) => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           ADD_WR(2) => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ADD_WR(1) => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           ADD_WR(0) => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           ADD_RD1(4) => datapath_i_n9, ADD_RD1(3) => 
                           datapath_i_n10, ADD_RD1(2) => datapath_i_n11, 
                           ADD_RD1(1) => datapath_i_n12, ADD_RD1(0) => 
                           datapath_i_n13, ADD_RD2(4) => 
                           curr_instruction_to_cu_i_20_port, ADD_RD2(3) => 
                           curr_instruction_to_cu_i_19_port, ADD_RD2(2) => 
                           curr_instruction_to_cu_i_18_port, ADD_RD2(1) => 
                           curr_instruction_to_cu_i_17_port, ADD_RD2(0) => 
                           curr_instruction_to_cu_i_16_port, DATAIN(31) => 
                           datapath_i_decode_stage_dp_n12, DATAIN(30) => 
                           datapath_i_decode_stage_dp_n13, DATAIN(29) => 
                           datapath_i_decode_stage_dp_n14, DATAIN(28) => 
                           datapath_i_decode_stage_dp_n15, DATAIN(27) => 
                           datapath_i_decode_stage_dp_n16, DATAIN(26) => 
                           datapath_i_decode_stage_dp_n17, DATAIN(25) => 
                           datapath_i_decode_stage_dp_n18, DATAIN(24) => 
                           datapath_i_decode_stage_dp_n19, DATAIN(23) => 
                           datapath_i_decode_stage_dp_n20, DATAIN(22) => 
                           datapath_i_decode_stage_dp_n21, DATAIN(21) => 
                           datapath_i_decode_stage_dp_n22, DATAIN(20) => 
                           datapath_i_decode_stage_dp_n23, DATAIN(19) => 
                           datapath_i_decode_stage_dp_n24, DATAIN(18) => 
                           datapath_i_decode_stage_dp_n25, DATAIN(17) => 
                           datapath_i_decode_stage_dp_n26, DATAIN(16) => 
                           datapath_i_decode_stage_dp_n27, DATAIN(15) => 
                           datapath_i_decode_stage_dp_n28, DATAIN(14) => 
                           datapath_i_decode_stage_dp_n29, DATAIN(13) => 
                           datapath_i_decode_stage_dp_n30, DATAIN(12) => 
                           datapath_i_decode_stage_dp_n31, DATAIN(11) => 
                           datapath_i_decode_stage_dp_n32, DATAIN(10) => 
                           datapath_i_decode_stage_dp_n33, DATAIN(9) => 
                           datapath_i_decode_stage_dp_n34, DATAIN(8) => 
                           datapath_i_decode_stage_dp_n35, DATAIN(7) => 
                           datapath_i_decode_stage_dp_n36, DATAIN(6) => 
                           datapath_i_decode_stage_dp_n37, DATAIN(5) => 
                           datapath_i_decode_stage_dp_n38, DATAIN(4) => 
                           datapath_i_decode_stage_dp_n39, DATAIN(3) => 
                           datapath_i_decode_stage_dp_n40, DATAIN(2) => 
                           datapath_i_decode_stage_dp_n41, DATAIN(1) => 
                           datapath_i_decode_stage_dp_n42, DATAIN(0) => 
                           datapath_i_decode_stage_dp_n43, OUT1(31) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, 
                           OUT1(30) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, 
                           OUT1(29) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, 
                           OUT1(28) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, 
                           OUT1(27) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, 
                           OUT1(26) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, 
                           OUT1(25) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, 
                           OUT1(24) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, 
                           OUT1(23) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, 
                           OUT1(22) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, 
                           OUT1(21) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, 
                           OUT1(20) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, 
                           OUT1(19) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, 
                           OUT1(18) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, 
                           OUT1(17) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, 
                           OUT1(16) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, 
                           OUT1(15) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, 
                           OUT1(14) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, 
                           OUT1(13) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, 
                           OUT1(12) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, 
                           OUT1(11) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, 
                           OUT1(10) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, 
                           OUT1(9) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, 
                           OUT1(8) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, 
                           OUT1(7) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, 
                           OUT1(6) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, 
                           OUT1(5) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, 
                           OUT1(4) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, 
                           OUT1(3) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, 
                           OUT1(2) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, 
                           OUT1(1) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, 
                           OUT1(0) => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, 
                           OUT2(31) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, 
                           OUT2(30) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, 
                           OUT2(29) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, 
                           OUT2(28) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, 
                           OUT2(27) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, 
                           OUT2(26) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, 
                           OUT2(25) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, 
                           OUT2(24) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, 
                           OUT2(23) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, 
                           OUT2(22) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, 
                           OUT2(21) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, 
                           OUT2(20) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, 
                           OUT2(19) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, 
                           OUT2(18) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, 
                           OUT2(17) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, 
                           OUT2(16) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, 
                           OUT2(15) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, 
                           OUT2(14) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, 
                           OUT2(13) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, 
                           OUT2(12) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, 
                           OUT2(11) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, 
                           OUT2(10) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, 
                           OUT2(9) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, 
                           OUT2(8) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, 
                           OUT2(7) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, 
                           OUT2(6) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, 
                           OUT2(5) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, 
                           OUT2(4) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, 
                           OUT2(3) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, 
                           OUT2(2) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, 
                           OUT2(1) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, 
                           OUT2(0) => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, 
                           RESET_BAR => RST);
   datapath_i_execute_stage_dp_general_alu_i : general_alu_N32 port map( clk =>
                           CLK, zero_mul_detect => n_1414, mul_exeception => 
                           n_1415, FUNC(0) => n1925, FUNC(1) => 
                           datapath_i_execute_stage_dp_n7, FUNC(2) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port, 
                           FUNC(3) => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port, 
                           DATA1(31) => datapath_i_execute_stage_dp_opa_31_port
                           , DATA1(30) => 
                           datapath_i_execute_stage_dp_opa_30_port, DATA1(29) 
                           => datapath_i_execute_stage_dp_opa_29_port, 
                           DATA1(28) => datapath_i_execute_stage_dp_opa_28_port
                           , DATA1(27) => 
                           datapath_i_execute_stage_dp_opa_27_port, DATA1(26) 
                           => datapath_i_execute_stage_dp_opa_26_port, 
                           DATA1(25) => datapath_i_execute_stage_dp_opa_25_port
                           , DATA1(24) => 
                           datapath_i_execute_stage_dp_opa_24_port, DATA1(23) 
                           => datapath_i_execute_stage_dp_opa_23_port, 
                           DATA1(22) => datapath_i_execute_stage_dp_opa_22_port
                           , DATA1(21) => 
                           datapath_i_execute_stage_dp_opa_21_port, DATA1(20) 
                           => datapath_i_execute_stage_dp_opa_20_port, 
                           DATA1(19) => datapath_i_execute_stage_dp_opa_19_port
                           , DATA1(18) => 
                           datapath_i_execute_stage_dp_opa_18_port, DATA1(17) 
                           => datapath_i_execute_stage_dp_opa_17_port, 
                           DATA1(16) => datapath_i_execute_stage_dp_opa_16_port
                           , DATA1(15) => 
                           datapath_i_execute_stage_dp_opa_15_port, DATA1(14) 
                           => datapath_i_execute_stage_dp_opa_14_port, 
                           DATA1(13) => datapath_i_execute_stage_dp_opa_13_port
                           , DATA1(12) => 
                           datapath_i_execute_stage_dp_opa_12_port, DATA1(11) 
                           => datapath_i_execute_stage_dp_opa_11_port, 
                           DATA1(10) => datapath_i_execute_stage_dp_opa_10_port
                           , DATA1(9) => datapath_i_execute_stage_dp_opa_9_port
                           , DATA1(8) => datapath_i_execute_stage_dp_opa_8_port
                           , DATA1(7) => datapath_i_execute_stage_dp_opa_7_port
                           , DATA1(6) => datapath_i_execute_stage_dp_opa_6_port
                           , DATA1(5) => datapath_i_execute_stage_dp_opa_5_port
                           , DATA1(4) => datapath_i_execute_stage_dp_opa_4_port
                           , DATA1(3) => datapath_i_execute_stage_dp_opa_3_port
                           , DATA1(2) => datapath_i_execute_stage_dp_opa_2_port
                           , DATA1(1) => datapath_i_execute_stage_dp_opa_1_port
                           , DATA1(0) => datapath_i_execute_stage_dp_opa_0_port
                           , DATA2(31) => 
                           datapath_i_execute_stage_dp_opb_31_port, DATA2(30) 
                           => datapath_i_execute_stage_dp_opb_30_port, 
                           DATA2(29) => datapath_i_execute_stage_dp_opb_29_port
                           , DATA2(28) => 
                           datapath_i_execute_stage_dp_opb_28_port, DATA2(27) 
                           => datapath_i_execute_stage_dp_opb_27_port, 
                           DATA2(26) => datapath_i_execute_stage_dp_opb_26_port
                           , DATA2(25) => 
                           datapath_i_execute_stage_dp_opb_25_port, DATA2(24) 
                           => datapath_i_execute_stage_dp_opb_24_port, 
                           DATA2(23) => datapath_i_execute_stage_dp_opb_23_port
                           , DATA2(22) => 
                           datapath_i_execute_stage_dp_opb_22_port, DATA2(21) 
                           => datapath_i_execute_stage_dp_opb_21_port, 
                           DATA2(20) => datapath_i_execute_stage_dp_opb_20_port
                           , DATA2(19) => 
                           datapath_i_execute_stage_dp_opb_19_port, DATA2(18) 
                           => datapath_i_execute_stage_dp_opb_18_port, 
                           DATA2(17) => datapath_i_execute_stage_dp_opb_17_port
                           , DATA2(16) => 
                           datapath_i_execute_stage_dp_opb_16_port, DATA2(15) 
                           => datapath_i_execute_stage_dp_opb_15_port, 
                           DATA2(14) => datapath_i_execute_stage_dp_opb_14_port
                           , DATA2(13) => 
                           datapath_i_execute_stage_dp_opb_13_port, DATA2(12) 
                           => datapath_i_execute_stage_dp_opb_12_port, 
                           DATA2(11) => datapath_i_execute_stage_dp_opb_11_port
                           , DATA2(10) => 
                           datapath_i_execute_stage_dp_opb_10_port, DATA2(9) =>
                           datapath_i_execute_stage_dp_opb_9_port, DATA2(8) => 
                           datapath_i_execute_stage_dp_opb_8_port, DATA2(7) => 
                           datapath_i_execute_stage_dp_opb_7_port, DATA2(6) => 
                           datapath_i_execute_stage_dp_opb_6_port, DATA2(5) => 
                           datapath_i_execute_stage_dp_opb_5_port, DATA2(4) => 
                           datapath_i_execute_stage_dp_opb_4_port, DATA2(3) => 
                           datapath_i_execute_stage_dp_opb_3_port, DATA2(2) => 
                           datapath_i_execute_stage_dp_opb_2_port, DATA2(1) => 
                           datapath_i_execute_stage_dp_opb_1_port, DATA2(0) => 
                           datapath_i_execute_stage_dp_opb_0_port, cin => 
                           alu_cin_i, signed_notsigned => 
                           datapath_i_execute_stage_dp_n9, overflow => n_1416, 
                           OUTALU(31) => 
                           datapath_i_execute_stage_dp_alu_out_31_port, 
                           OUTALU(30) => 
                           datapath_i_execute_stage_dp_alu_out_30_port, 
                           OUTALU(29) => 
                           datapath_i_execute_stage_dp_alu_out_29_port, 
                           OUTALU(28) => 
                           datapath_i_execute_stage_dp_alu_out_28_port, 
                           OUTALU(27) => 
                           datapath_i_execute_stage_dp_alu_out_27_port, 
                           OUTALU(26) => 
                           datapath_i_execute_stage_dp_alu_out_26_port, 
                           OUTALU(25) => 
                           datapath_i_execute_stage_dp_alu_out_25_port, 
                           OUTALU(24) => 
                           datapath_i_execute_stage_dp_alu_out_24_port, 
                           OUTALU(23) => 
                           datapath_i_execute_stage_dp_alu_out_23_port, 
                           OUTALU(22) => 
                           datapath_i_execute_stage_dp_alu_out_22_port, 
                           OUTALU(21) => 
                           datapath_i_execute_stage_dp_alu_out_21_port, 
                           OUTALU(20) => 
                           datapath_i_execute_stage_dp_alu_out_20_port, 
                           OUTALU(19) => 
                           datapath_i_execute_stage_dp_alu_out_19_port, 
                           OUTALU(18) => 
                           datapath_i_execute_stage_dp_alu_out_18_port, 
                           OUTALU(17) => 
                           datapath_i_execute_stage_dp_alu_out_17_port, 
                           OUTALU(16) => 
                           datapath_i_execute_stage_dp_alu_out_16_port, 
                           OUTALU(15) => 
                           datapath_i_execute_stage_dp_alu_out_15_port, 
                           OUTALU(14) => 
                           datapath_i_execute_stage_dp_alu_out_14_port, 
                           OUTALU(13) => 
                           datapath_i_execute_stage_dp_alu_out_13_port, 
                           OUTALU(12) => 
                           datapath_i_execute_stage_dp_alu_out_12_port, 
                           OUTALU(11) => 
                           datapath_i_execute_stage_dp_alu_out_11_port, 
                           OUTALU(10) => 
                           datapath_i_execute_stage_dp_alu_out_10_port, 
                           OUTALU(9) => 
                           datapath_i_execute_stage_dp_alu_out_9_port, 
                           OUTALU(8) => 
                           datapath_i_execute_stage_dp_alu_out_8_port, 
                           OUTALU(7) => 
                           datapath_i_execute_stage_dp_alu_out_7_port, 
                           OUTALU(6) => 
                           datapath_i_execute_stage_dp_alu_out_6_port, 
                           OUTALU(5) => 
                           datapath_i_execute_stage_dp_alu_out_5_port, 
                           OUTALU(4) => 
                           datapath_i_execute_stage_dp_alu_out_4_port, 
                           OUTALU(3) => 
                           datapath_i_execute_stage_dp_alu_out_3_port, 
                           OUTALU(2) => 
                           datapath_i_execute_stage_dp_alu_out_2_port, 
                           OUTALU(1) => 
                           datapath_i_execute_stage_dp_alu_out_1_port, 
                           OUTALU(0) => 
                           datapath_i_execute_stage_dp_alu_out_0_port, rst_BAR 
                           => RST);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_31_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_31_port, EN => n309, Z 
                           => DRAM_ADDRESS_31_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_30_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_30_port, EN => n309, Z 
                           => DRAM_ADDRESS_30_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_29_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_29_port, EN => n2321, Z 
                           => DRAM_ADDRESS_29_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_28_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_28_port, EN => n2321, Z 
                           => DRAM_ADDRESS_28_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_27_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_27_port, EN => n2321, Z 
                           => DRAM_ADDRESS_27_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_26_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_26_port, EN => n2321, Z 
                           => DRAM_ADDRESS_26_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_25_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_25_port, EN => n2321, Z 
                           => DRAM_ADDRESS_25_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_24_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_24_port, EN => n2321, Z 
                           => DRAM_ADDRESS_24_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_23_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_23_port, EN => n2321, Z 
                           => DRAM_ADDRESS_23_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_22_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_22_port, EN => n2321, Z 
                           => DRAM_ADDRESS_22_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_21_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_21_port, EN => n2321, Z 
                           => DRAM_ADDRESS_21_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_20_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_20_port, EN => n2321, Z 
                           => DRAM_ADDRESS_20_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_19_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_19_port, EN => n2321, Z 
                           => DRAM_ADDRESS_19_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_18_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_18_port, EN => n2321, Z 
                           => DRAM_ADDRESS_18_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_17_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_17_port, EN => n309, Z 
                           => DRAM_ADDRESS_17_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_16_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_16_port, EN => n2321, Z 
                           => DRAM_ADDRESS_16_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_15_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_15_port, EN => n2321, Z 
                           => DRAM_ADDRESS_15_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_14_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_14_port, EN => n2321, Z 
                           => DRAM_ADDRESS_14_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_13_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_13_port, EN => n309, Z 
                           => DRAM_ADDRESS_13_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_12_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_12_port, EN => n2321, Z 
                           => DRAM_ADDRESS_12_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_11_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_11_port, EN => n2321, Z 
                           => DRAM_ADDRESS_11_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_10_inst : TBUF_X1 port map( A =>
                           datapath_i_alu_output_val_i_10_port, EN => n2321, Z 
                           => DRAM_ADDRESS_10_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_9_port, EN => n309, Z =>
                           DRAM_ADDRESS_9_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_8_port, EN => n309, Z =>
                           DRAM_ADDRESS_8_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_7_port, EN => n2321, Z 
                           => DRAM_ADDRESS_7_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_6_port, EN => n309, Z =>
                           DRAM_ADDRESS_6_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_5_port, EN => n2321, Z 
                           => DRAM_ADDRESS_5_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_4_port, EN => n309, Z =>
                           DRAM_ADDRESS_4_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_3_port, EN => n2321, Z 
                           => DRAM_ADDRESS_3_port);
   datapath_i_memory_stage_dp_DRAM_ADDRESS_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_alu_output_val_i_2_port, EN => n309, Z =>
                           DRAM_ADDRESS_2_port);
   datapath_i_memory_stage_dp_DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_9_port, EN => n2323, Z => 
                           DRAM_DATA(9));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_31_port, EN => n2323, Z =>
                           DRAM_DATA(31));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_30_port, EN => n2323, Z =>
                           DRAM_DATA(30));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_29_port, EN => n2323, Z =>
                           DRAM_DATA(29));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_28_port, EN => n2323, Z =>
                           DRAM_DATA(28));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_27_port, EN => n2323, Z =>
                           DRAM_DATA(27));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_26_port, EN => n2323, Z =>
                           DRAM_DATA(26));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_25_port, EN => n2323, Z =>
                           DRAM_DATA(25));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_24_port, EN => n2323, Z =>
                           DRAM_DATA(24));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_23_port, EN => n2323, Z =>
                           DRAM_DATA(23));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_22_port, EN => n2323, Z =>
                           DRAM_DATA(22));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_21_port, EN => n2323, Z =>
                           DRAM_DATA(21));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_20_port, EN => n2323, Z =>
                           DRAM_DATA(20));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_19_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(19));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_18_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(18));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_17_port, EN => n2323, Z =>
                           DRAM_DATA(17));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_16_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(16));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_15_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(15));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_14_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(14));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_13_port, EN => n2323, Z =>
                           DRAM_DATA(13));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_12_port, EN => n2323, Z =>
                           DRAM_DATA(12));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_11_port, EN => n2323, Z =>
                           DRAM_DATA(11));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_10_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(10));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_8_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(8));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_7_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(7));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_6_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(6));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_5_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(5));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_4_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(4));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_3_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(3));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_2_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(2));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_1_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(1));
   datapath_i_memory_stage_dp_DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => 
                           datapath_i_value_to_mem_i_0_port, EN => 
                           datapath_i_memory_stage_dp_n2, Z => DRAM_DATA(0));
   cu_i_e_reg_D_I_0_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_0_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_0_port, QN => 
                           n_1417);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_0_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_1_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_2_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_3_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_4_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_5_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_6_inst : 
                           DLH_X1 port map( G => n2320, D => datapath_i_n18, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_7_inst : 
                           DLH_X1 port map( G => n2320, D => datapath_i_n17, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_8_inst : 
                           DLH_X1 port map( G => n2320, D => datapath_i_n16, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_9_inst : 
                           DLH_X1 port map( G => n2320, D => datapath_i_n15, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n310, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n310, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_immediate_extended_val_reg_31_inst : 
                           DLH_X1 port map( G => n2320, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_0_inst
                           : DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_0_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_1_inst
                           : DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_1_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_2_inst
                           : DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_2_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_3_inst
                           : DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_3_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_4_inst
                           : DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_4_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_5_inst
                           : DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_5_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_6_inst
                           : DLH_X1 port map( G => n2324, D => datapath_i_n18, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_7_inst
                           : DLH_X1 port map( G => n2324, D => datapath_i_n17, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_8_inst
                           : DLH_X1 port map( G => n2324, D => datapath_i_n16, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port);
   datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_9_inst
                           : DLH_X1 port map( G => n2324, D => datapath_i_n15, 
                           Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_10_inst : 
                           DLH_X1 port map( G => n2324, D => datapath_i_n14, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_11_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_11_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_12_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_12_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_13_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_13_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_14_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_14_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_15_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_15_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_16_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_16_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_17_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_17_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_18_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_18_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_19_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_19_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_20_inst : 
                           DLH_X1 port map( G => n2324, D => 
                           curr_instruction_to_cu_i_20_port, Q => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_21_inst : 
                           DLH_X1 port map( G => n2324, D => datapath_i_n13, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_22_inst : 
                           DLH_X1 port map( G => n2324, D => datapath_i_n12, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_23_inst : 
                           DLH_X1 port map( G => n2324, D => datapath_i_n11, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_24_inst : 
                           DLH_X1 port map( G => n2324, D => datapath_i_n10, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port);
   
                           datapath_i_decode_stage_dp_sign_extension_logic_jump_extended_val_reg_25_inst : 
                           DLH_X1 port map( G => n2324, D => datapath_i_n9, Q 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port);
   cu_i_wb_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n1932, CK => CLK, RN => RST
                           , Q => cu_i_cw3_6_port, QN => n_1418);
   cu_i_wb_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n131, CK => CLK, RN =>
                           RST, Q => n_1419, QN => n699);
   cu_i_m_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_8_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_8_port, QN => n_1420);
   cu_i_m_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_7_port, CK => CLK
                           , RN => RST, Q => cu_i_cw2_7_port, QN => n_1421);
   cu_i_m_reg_D_I_6_Q_reg : DFFR_X1 port map( D => cu_i_n127, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_6_port, QN => n_1422);
   cu_i_m_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_n126, CK => CLK, RN => 
                           RST, Q => cu_i_cw2_5_port, QN => n2318);
   cu_i_m_reg_D_I_4_Q_reg : DFFR_X1 port map( D => cu_i_cw1_i_4_port, CK => CLK
                           , RN => RST, Q => n_1423, QN => n756);
   cu_i_e_reg_D_I_13_Q_reg : DFFR_X1 port map( D => n2320, CK => CLK, RN => RST
                           , Q => n_1424, QN => n2319);
   cu_i_e_reg_D_I_12_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_8_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_12_port, QN => n_1425)
                           ;
   cu_i_e_reg_D_I_11_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_7_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_11_port, QN => n_1426)
                           ;
   cu_i_e_reg_D_I_10_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_6_port, CK =>
                           CLK, RN => RST, Q => cu_i_cw1_10_port, QN => n_1427)
                           ;
   cu_i_e_reg_D_I_8_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_4_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_8_port, QN => n_1428);
   cu_i_e_reg_D_I_7_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_3_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_7_port, QN => n_1429);
   cu_i_e_reg_D_I_6_Q_reg : DFFR_X1 port map( D => n311, CK => CLK, RN => RST, 
                           Q => cu_i_cw1_6_port, QN => n_1430);
   cu_i_e_reg_D_I_5_Q_reg : DFFR_X1 port map( D => cu_i_cmd_word_1_port, CK => 
                           CLK, RN => RST, Q => cu_i_cw1_5_port, QN => n_1431);
   cu_i_e_reg_D_I_4_Q_reg : DFFR_X1 port map( D => n1152, CK => CLK, RN => RST,
                           Q => cu_i_cw1_4_port, QN => n_1432);
   cu_i_e_reg_D_I_3_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_3_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_3_port, QN => 
                           n_1433);
   cu_i_e_reg_D_I_2_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_2_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_2_port, QN => 
                           n_1434);
   cu_i_e_reg_D_I_1_Q_reg : DFFR_X1 port map( D => cu_i_cmd_alu_op_type_1_port,
                           CK => CLK, RN => RST, Q => cu_i_cw1_1_port, QN => 
                           n_1435);
   datapath_i_memory_stage_dp_delay_regg_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_31_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_31_port, QN 
                           => n_1436);
   datapath_i_memory_stage_dp_delay_regg_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_30_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_30_port, QN 
                           => n_1437);
   datapath_i_memory_stage_dp_delay_regg_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_29_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_29_port, QN 
                           => n_1438);
   datapath_i_memory_stage_dp_delay_regg_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_28_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_28_port, QN 
                           => n_1439);
   datapath_i_memory_stage_dp_delay_regg_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_27_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_27_port, QN 
                           => n_1440);
   datapath_i_memory_stage_dp_delay_regg_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_26_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_26_port, QN 
                           => n_1441);
   datapath_i_memory_stage_dp_delay_regg_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_25_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_25_port, QN 
                           => n_1442);
   datapath_i_memory_stage_dp_delay_regg_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_24_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_24_port, QN 
                           => n_1443);
   datapath_i_memory_stage_dp_delay_regg_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_23_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_23_port, QN 
                           => n_1444);
   datapath_i_memory_stage_dp_delay_regg_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_22_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_22_port, QN 
                           => n_1445);
   datapath_i_memory_stage_dp_delay_regg_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_21_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_21_port, QN 
                           => n_1446);
   datapath_i_memory_stage_dp_delay_regg_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_20_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_20_port, QN 
                           => n_1447);
   datapath_i_memory_stage_dp_delay_regg_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_19_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_19_port, QN 
                           => n_1448);
   datapath_i_memory_stage_dp_delay_regg_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_18_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_18_port, QN 
                           => n_1449);
   datapath_i_memory_stage_dp_delay_regg_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_17_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_17_port, QN 
                           => n_1450);
   datapath_i_memory_stage_dp_delay_regg_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_16_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_16_port, QN 
                           => n_1451);
   datapath_i_memory_stage_dp_delay_regg_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_15_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_15_port, QN 
                           => n_1452);
   datapath_i_memory_stage_dp_delay_regg_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_14_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_14_port, QN 
                           => n_1453);
   datapath_i_memory_stage_dp_delay_regg_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_13_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_13_port, QN 
                           => n_1454);
   datapath_i_memory_stage_dp_delay_regg_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_12_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_12_port, QN 
                           => n_1455);
   datapath_i_memory_stage_dp_delay_regg_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_11_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_11_port, QN 
                           => n_1456);
   datapath_i_memory_stage_dp_delay_regg_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_10_port, CK => CLK, RN 
                           => RST, Q => datapath_i_data_from_alu_i_10_port, QN 
                           => n_1457);
   datapath_i_memory_stage_dp_delay_regg_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_9_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_9_port, QN => 
                           n_1458);
   datapath_i_memory_stage_dp_delay_regg_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_8_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_8_port, QN => 
                           n_1459);
   datapath_i_memory_stage_dp_delay_regg_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_7_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_7_port, QN => 
                           n_1460);
   datapath_i_memory_stage_dp_delay_regg_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_6_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_6_port, QN => 
                           n_1461);
   datapath_i_memory_stage_dp_delay_regg_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_5_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_5_port, QN => 
                           n_1462);
   datapath_i_memory_stage_dp_delay_regg_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_4_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_4_port, QN => 
                           n_1463);
   datapath_i_memory_stage_dp_delay_regg_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_3_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_3_port, QN => 
                           n_1464);
   datapath_i_memory_stage_dp_delay_regg_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_2_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_2_port, QN => 
                           n_1465);
   datapath_i_memory_stage_dp_delay_regg_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_1_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_1_port, QN => 
                           n_1466);
   datapath_i_memory_stage_dp_delay_regg_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_alu_output_val_i_0_port, CK => CLK, RN =>
                           RST, Q => datapath_i_data_from_alu_i_0_port, QN => 
                           n_1467);
   datapath_i_memory_stage_dp_lmd_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_31_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_31_port, QN => n_1468)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_30_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_30_port, QN => n_1469)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_29_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_29_port, QN => n_1470)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_28_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_28_port, QN => n_1471)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_27_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_27_port, QN => n_1472)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_26_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_26_port, QN => n_1473)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_25_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_25_port, QN => n_1474)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_24_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_24_port, QN => n_1475)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_23_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_23_port, QN => n_1476)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_22_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_22_port, QN => n_1477)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_21_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_21_port, QN => n_1478)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_20_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_20_port, QN => n_1479)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_19_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_19_port, QN => n_1480)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_18_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_18_port, QN => n_1481)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_17_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_17_port, QN => n_1482)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_16_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_16_port, QN => n_1483)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_15_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_15_port, QN => n_1484)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_14_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_14_port, QN => n_1485)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_13_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_13_port, QN => n_1486)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_12_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_12_port, QN => n_1487)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_11_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_11_port, QN => n_1488)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_10_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_data_from_memory_i_10_port, QN => n_1489)
                           ;
   datapath_i_memory_stage_dp_lmd_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_9_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_9_port, QN => n_1490);
   datapath_i_memory_stage_dp_lmd_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_8_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_8_port, QN => n_1491);
   datapath_i_memory_stage_dp_lmd_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_7_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_7_port, QN => n_1492);
   datapath_i_memory_stage_dp_lmd_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_6_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_6_port, QN => n_1493);
   datapath_i_memory_stage_dp_lmd_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_5_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_5_port, QN => n_1494);
   datapath_i_memory_stage_dp_lmd_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_4_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_4_port, QN => n_1495);
   datapath_i_memory_stage_dp_lmd_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_3_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_3_port, QN => n_1496);
   datapath_i_memory_stage_dp_lmd_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_2_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_2_port, QN => n_1497);
   datapath_i_memory_stage_dp_lmd_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_1_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_1_port, QN => n_1498);
   datapath_i_memory_stage_dp_lmd_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_memory_stage_dp_data_ir_0_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_data_from_memory_i_0_port, QN => n_1499);
   datapath_i_execute_stage_dp_reg_del_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_31_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_31_port, QN => n_1500);
   datapath_i_execute_stage_dp_reg_del_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_30_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_30_port, QN => n_1501);
   datapath_i_execute_stage_dp_reg_del_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_29_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_29_port, QN => n_1502);
   datapath_i_execute_stage_dp_reg_del_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_28_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_28_port, QN => n_1503);
   datapath_i_execute_stage_dp_reg_del_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_27_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_27_port, QN => n_1504);
   datapath_i_execute_stage_dp_reg_del_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_26_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_26_port, QN => n_1505);
   datapath_i_execute_stage_dp_reg_del_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_25_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_25_port, QN => n_1506);
   datapath_i_execute_stage_dp_reg_del_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_24_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_24_port, QN => n_1507);
   datapath_i_execute_stage_dp_reg_del_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_23_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_23_port, QN => n_1508);
   datapath_i_execute_stage_dp_reg_del_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_22_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_22_port, QN => n_1509);
   datapath_i_execute_stage_dp_reg_del_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_21_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_21_port, QN => n_1510);
   datapath_i_execute_stage_dp_reg_del_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_20_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_20_port, QN => n_1511);
   datapath_i_execute_stage_dp_reg_del_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_19_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_19_port, QN => n_1512);
   datapath_i_execute_stage_dp_reg_del_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_18_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_18_port, QN => n_1513);
   datapath_i_execute_stage_dp_reg_del_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_17_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_17_port, QN => n_1514);
   datapath_i_execute_stage_dp_reg_del_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_16_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_16_port, QN => n_1515);
   datapath_i_execute_stage_dp_reg_del_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_15_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_15_port, QN => n_1516);
   datapath_i_execute_stage_dp_reg_del_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_14_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_14_port, QN => n_1517);
   datapath_i_execute_stage_dp_reg_del_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_13_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_13_port, QN => n_1518);
   datapath_i_execute_stage_dp_reg_del_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_12_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_12_port, QN => n_1519);
   datapath_i_execute_stage_dp_reg_del_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_11_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_11_port, QN => n_1520);
   datapath_i_execute_stage_dp_reg_del_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_10_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_10_port, QN => n_1521);
   datapath_i_execute_stage_dp_reg_del_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_9_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_9_port, QN => n_1522);
   datapath_i_execute_stage_dp_reg_del_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_8_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_8_port, QN => n_1523);
   datapath_i_execute_stage_dp_reg_del_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_7_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_7_port, QN => n_1524);
   datapath_i_execute_stage_dp_reg_del_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_6_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_6_port, QN => n_1525);
   datapath_i_execute_stage_dp_reg_del_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_5_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_5_port, QN => n_1526);
   datapath_i_execute_stage_dp_reg_del_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_4_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_4_port, QN => n_1527);
   datapath_i_execute_stage_dp_reg_del_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_3_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_3_port, QN => n_1528);
   datapath_i_execute_stage_dp_reg_del_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_2_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_2_port, QN => n_1529);
   datapath_i_execute_stage_dp_reg_del_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_1_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_1_port, QN => n_1530);
   datapath_i_execute_stage_dp_reg_del_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_val_b_i_0_port, CK => CLK, RN => RST, Q 
                           => datapath_i_value_to_mem_i_0_port, QN => n_1531);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_31_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_31_port, QN => n_1532);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_30_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_30_port, QN => n_1533);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_29_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_29_port, QN => n_1534);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_28_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_28_port, QN => n_1535);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_27_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_27_port, QN => n_1536);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_26_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_26_port, QN => n_1537);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_25_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_25_port, QN => n_1538);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_24_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_24_port, QN => n_1539);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_23_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_23_port, QN => n_1540);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_22_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_22_port, QN => n_1541);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_21_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_21_port, QN => n_1542);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_20_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_20_port, QN => n_1543);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_19_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_19_port, QN => n_1544);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_18_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_18_port, QN => n_1545);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_17_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_17_port, QN => n_1546);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_16_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_16_port, QN => n_1547);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_15_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_15_port, QN => n_1548);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_14_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_14_port, QN => n_1549);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_13_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_13_port, QN => n_1550);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_12_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_12_port, QN => n_1551);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_11_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_11_port, QN => n_1552);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_execute_stage_dp_alu_out_10_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_10_port, QN => n_1553);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_9_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_9_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_9_port, QN => n_1554);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_8_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_8_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_8_port, QN => n_1555);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_7_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_7_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_7_port, QN => n_1556);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_6_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_6_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_6_port, QN => n_1557);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_5_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_5_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_5_port, QN => n_1558);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_4_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_4_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_4_port, QN => n_1559);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_3_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_3_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_3_port, QN => n_1560);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_2_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_2_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_2_port, QN => n_1561);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_1_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_1_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_1_port, QN => n_1562);
   datapath_i_execute_stage_dp_alu_reg_out_D_I_0_Q_reg : DFFR_X1 port map( D =>
                           datapath_i_execute_stage_dp_alu_out_0_port, CK => 
                           CLK, RN => RST, Q => 
                           datapath_i_alu_output_val_i_0_port, QN => n_1563);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_32_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_32_port, CK 
                           => CLK, RN => RST, Q => n_1564, QN => n703);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_31_port, CK 
                           => CLK, RN => RST, Q => n_1565, QN => n727);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_30_port, CK 
                           => CLK, RN => RST, Q => n_1566, QN => n726);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_29_port, CK 
                           => CLK, RN => RST, Q => n_1567, QN => n725);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_28_port, CK 
                           => CLK, RN => RST, Q => n_1568, QN => n724);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_27_port, CK 
                           => CLK, RN => RST, Q => n_1569, QN => n691);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_26_port, CK 
                           => CLK, RN => RST, Q => n_1570, QN => n723);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_25_port, CK 
                           => CLK, RN => RST, Q => n_1571, QN => n722);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_24_port, CK 
                           => CLK, RN => RST, Q => n_1572, QN => n721);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_23_port, CK 
                           => CLK, RN => RST, Q => n_1573, QN => n720);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_22_port, CK 
                           => CLK, RN => RST, Q => n_1574, QN => n719);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_21_port, CK 
                           => CLK, RN => RST, Q => n_1575, QN => n718);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_20_port, CK 
                           => CLK, RN => RST, Q => n_1576, QN => n717);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_19_port, CK 
                           => CLK, RN => RST, Q => n_1577, QN => n716);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_18_port, CK 
                           => CLK, RN => RST, Q => n_1578, QN => n715);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_17_port, CK 
                           => CLK, RN => RST, Q => n_1579, QN => n714);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_16_port, CK 
                           => CLK, RN => RST, Q => n_1580, QN => n713);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_15_port, CK 
                           => CLK, RN => RST, Q => n_1581, QN => n712);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_14_port, CK 
                           => CLK, RN => RST, Q => n_1582, QN => n711);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_13_port, CK 
                           => CLK, RN => RST, Q => n_1583, QN => n710);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_12_port, CK 
                           => CLK, RN => RST, Q => n_1584, QN => n709);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_11_port, CK 
                           => CLK, RN => RST, Q => n_1585, QN => n708);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_decode_stage_dp_pc_delay2_10_port, CK 
                           => CLK, RN => RST, Q => n_1586, QN => n707);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_9_port, CK 
                           => CLK, RN => RST, Q => n_1587, QN => n706);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_8_port, CK 
                           => CLK, RN => RST, Q => n_1588, QN => n705);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_7_port, CK 
                           => CLK, RN => RST, Q => n_1589, QN => n732);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_6_port, CK 
                           => CLK, RN => RST, Q => n_1590, QN => n731);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_5_port, CK 
                           => CLK, RN => RST, Q => n_1591, QN => n730);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_4_port, CK 
                           => CLK, RN => RST, Q => n_1592, QN => n729);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_3_port, CK 
                           => CLK, RN => RST, Q => n_1593, QN => n728);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_2_port, CK 
                           => CLK, RN => RST, Q => n_1594, QN => n734);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_1_port, CK 
                           => CLK, RN => RST, Q => n_1595, QN => n733);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_32_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_31_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_32_port, QN => 
                           n_1596);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_31_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_30_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_31_port, QN => 
                           n_1597);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_30_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_29_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_30_port, QN => 
                           n_1598);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_29_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_28_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_29_port, QN => 
                           n_1599);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_28_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_27_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_28_port, QN => 
                           n_1600);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_27_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_26_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_27_port, QN => 
                           n_1601);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_26_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_25_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_26_port, QN => 
                           n_1602);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_24_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_25_port, QN => 
                           n_1603);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_23_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_24_port, QN => 
                           n_1604);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_22_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_23_port, QN => 
                           n_1605);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_21_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_22_port, QN => 
                           n_1606);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_20_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_21_port, QN => 
                           n_1607);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_19_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_20_port, QN => 
                           n_1608);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_18_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_19_port, QN => 
                           n_1609);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_17_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_18_port, QN => 
                           n_1610);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_16_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_17_port, QN => 
                           n_1611);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_15_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_16_port, QN => 
                           n_1612);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_14_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_15_port, QN => 
                           n_1613);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_13_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_14_port, QN => 
                           n_1614);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_12_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_13_port, QN => 
                           n_1615);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_11_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_12_port, QN => 
                           n_1616);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_10_port, CK => CLK
                           , RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_11_port, QN => 
                           n_1617);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_9_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_10_port, QN => 
                           n_1618);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_8_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_9_port, QN => 
                           n_1619);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_7_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_8_port, QN => 
                           n_1620);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_6_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_7_port, QN => 
                           n_1621);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_5_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_6_port, QN => 
                           n_1622);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_4_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_5_port, QN => 
                           n_1623);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_3_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_4_port, QN => 
                           n_1624);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_2_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_3_port, QN => 
                           n_1625);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_1_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_2_port, QN => 
                           n_1626);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_decode_0_port, CK => CLK,
                           RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_1_port, QN => 
                           n_1627);
   datapath_i_decode_stage_dp_pc_delay_reg1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n2324, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay2_0_port, QN => 
                           n_1628);
   datapath_i_decode_stage_dp_reg_immediate_D_I_25_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_25_port, QN 
                           => n_1629);
   datapath_i_decode_stage_dp_reg_immediate_D_I_24_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_24_port, QN 
                           => n_1630);
   datapath_i_decode_stage_dp_reg_immediate_D_I_23_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_23_port, QN 
                           => n_1631);
   datapath_i_decode_stage_dp_reg_immediate_D_I_22_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_22_port, QN 
                           => n_1632);
   datapath_i_decode_stage_dp_reg_immediate_D_I_21_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_21_port, QN 
                           => n_1633);
   datapath_i_decode_stage_dp_reg_immediate_D_I_20_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_20_port, QN 
                           => n_1634);
   datapath_i_decode_stage_dp_reg_immediate_D_I_19_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_19_port, QN 
                           => n_1635);
   datapath_i_decode_stage_dp_reg_immediate_D_I_18_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_18_port, QN 
                           => n_1636);
   datapath_i_decode_stage_dp_reg_immediate_D_I_17_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_17_port, QN 
                           => n_1637);
   datapath_i_decode_stage_dp_reg_immediate_D_I_16_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_16_port, QN 
                           => n_1638);
   datapath_i_decode_stage_dp_reg_immediate_D_I_15_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_15_port, QN 
                           => n_1639);
   datapath_i_decode_stage_dp_reg_immediate_D_I_14_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_14_port, QN 
                           => n_1640);
   datapath_i_decode_stage_dp_reg_immediate_D_I_13_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_13_port, QN 
                           => n_1641);
   datapath_i_decode_stage_dp_reg_immediate_D_I_12_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_12_port, QN 
                           => n_1642);
   datapath_i_decode_stage_dp_reg_immediate_D_I_11_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_11_port, QN 
                           => n_1643);
   datapath_i_decode_stage_dp_reg_immediate_D_I_10_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           , CK => datapath_i_decode_stage_dp_clk_immediate, RN
                           => RST, Q => datapath_i_val_immediate_i_10_port, QN 
                           => n_1644);
   datapath_i_decode_stage_dp_reg_immediate_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_9_port, QN 
                           => n_1645);
   datapath_i_decode_stage_dp_reg_immediate_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_8_port, QN 
                           => n_1646);
   datapath_i_decode_stage_dp_reg_immediate_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_7_port, QN 
                           => n_1647);
   datapath_i_decode_stage_dp_reg_immediate_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_6_port, QN 
                           => n_1648);
   datapath_i_decode_stage_dp_reg_immediate_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_5_port, QN 
                           => n_1649);
   datapath_i_decode_stage_dp_reg_immediate_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_4_port, QN 
                           => n_1650);
   datapath_i_decode_stage_dp_reg_immediate_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_3_port, QN 
                           => n_1651);
   datapath_i_decode_stage_dp_reg_immediate_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_2_port, QN 
                           => n_1652);
   datapath_i_decode_stage_dp_reg_immediate_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_1_port, QN 
                           => n_1653);
   datapath_i_decode_stage_dp_reg_immediate_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port,
                           CK => datapath_i_decode_stage_dp_clk_immediate, RN 
                           => RST, Q => datapath_i_val_immediate_i_0_port, QN 
                           => n_1654);
   datapath_i_decode_stage_dp_reg_b_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_31_port, 
                           QN => n764);
   datapath_i_decode_stage_dp_reg_b_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_30_port, 
                           QN => n763);
   datapath_i_decode_stage_dp_reg_b_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_29_port, 
                           QN => n762);
   datapath_i_decode_stage_dp_reg_b_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_28_port, 
                           QN => n761);
   datapath_i_decode_stage_dp_reg_b_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_27_port, 
                           QN => n760);
   datapath_i_decode_stage_dp_reg_b_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_26_port, 
                           QN => n759);
   datapath_i_decode_stage_dp_reg_b_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_25_port, 
                           QN => n758);
   datapath_i_decode_stage_dp_reg_b_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_24_port, 
                           QN => n_1655);
   datapath_i_decode_stage_dp_reg_b_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_23_port, 
                           QN => n_1656);
   datapath_i_decode_stage_dp_reg_b_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_22_port, 
                           QN => n_1657);
   datapath_i_decode_stage_dp_reg_b_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_21_port, 
                           QN => n_1658);
   datapath_i_decode_stage_dp_reg_b_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_20_port, 
                           QN => n_1659);
   datapath_i_decode_stage_dp_reg_b_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_19_port, 
                           QN => n_1660);
   datapath_i_decode_stage_dp_reg_b_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_18_port, 
                           QN => n_1661);
   datapath_i_decode_stage_dp_reg_b_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_17_port, 
                           QN => n_1662);
   datapath_i_decode_stage_dp_reg_b_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_16_port, 
                           QN => n_1663);
   datapath_i_decode_stage_dp_reg_b_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_15_port, 
                           QN => n_1664);
   datapath_i_decode_stage_dp_reg_b_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_14_port, 
                           QN => n_1665);
   datapath_i_decode_stage_dp_reg_b_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_13_port, 
                           QN => n_1666);
   datapath_i_decode_stage_dp_reg_b_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_12_port, 
                           QN => n_1667);
   datapath_i_decode_stage_dp_reg_b_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_11_port, 
                           QN => n_1668);
   datapath_i_decode_stage_dp_reg_b_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_b_i_10_port, 
                           QN => n_1669);
   datapath_i_decode_stage_dp_reg_b_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_9_port, QN 
                           => n_1670);
   datapath_i_decode_stage_dp_reg_b_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_8_port, QN 
                           => n_1671);
   datapath_i_decode_stage_dp_reg_b_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_7_port, QN 
                           => n_1672);
   datapath_i_decode_stage_dp_reg_b_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_6_port, QN 
                           => n_1673);
   datapath_i_decode_stage_dp_reg_b_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_5_port, QN 
                           => n_1674);
   datapath_i_decode_stage_dp_reg_b_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_4_port, QN 
                           => n_1675);
   datapath_i_decode_stage_dp_reg_b_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_3_port, QN 
                           => n_1676);
   datapath_i_decode_stage_dp_reg_b_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_2_port, QN 
                           => n_1677);
   datapath_i_decode_stage_dp_reg_b_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_1_port, QN 
                           => n_1678);
   datapath_i_decode_stage_dp_reg_b_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_b_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_b_i_0_port, QN 
                           => n_1679);
   datapath_i_decode_stage_dp_reg_a_D_I_31_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_31_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_31_port, 
                           QN => n_1680);
   datapath_i_decode_stage_dp_reg_a_D_I_30_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_30_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_30_port, 
                           QN => n_1681);
   datapath_i_decode_stage_dp_reg_a_D_I_29_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_29_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_29_port, 
                           QN => n_1682);
   datapath_i_decode_stage_dp_reg_a_D_I_28_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_28_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_28_port, 
                           QN => n_1683);
   datapath_i_decode_stage_dp_reg_a_D_I_27_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_27_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_27_port, 
                           QN => n_1684);
   datapath_i_decode_stage_dp_reg_a_D_I_26_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_26_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_26_port, 
                           QN => n_1685);
   datapath_i_decode_stage_dp_reg_a_D_I_25_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_25_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_25_port, 
                           QN => n_1686);
   datapath_i_decode_stage_dp_reg_a_D_I_24_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_24_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_24_port, 
                           QN => n_1687);
   datapath_i_decode_stage_dp_reg_a_D_I_23_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_23_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_23_port, 
                           QN => n_1688);
   datapath_i_decode_stage_dp_reg_a_D_I_22_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_22_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_22_port, 
                           QN => n_1689);
   datapath_i_decode_stage_dp_reg_a_D_I_21_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_21_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_21_port, 
                           QN => n_1690);
   datapath_i_decode_stage_dp_reg_a_D_I_20_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_20_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_20_port, 
                           QN => n_1691);
   datapath_i_decode_stage_dp_reg_a_D_I_19_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_19_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_19_port, 
                           QN => n_1692);
   datapath_i_decode_stage_dp_reg_a_D_I_18_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_18_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_18_port, 
                           QN => n_1693);
   datapath_i_decode_stage_dp_reg_a_D_I_17_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_17_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_17_port, 
                           QN => n_1694);
   datapath_i_decode_stage_dp_reg_a_D_I_16_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_16_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_16_port, 
                           QN => n_1695);
   datapath_i_decode_stage_dp_reg_a_D_I_15_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_15_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_15_port, 
                           QN => n_1696);
   datapath_i_decode_stage_dp_reg_a_D_I_14_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_14_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_14_port, 
                           QN => n_1697);
   datapath_i_decode_stage_dp_reg_a_D_I_13_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_13_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_13_port, 
                           QN => n_1698);
   datapath_i_decode_stage_dp_reg_a_D_I_12_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_12_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_12_port, 
                           QN => n_1699);
   datapath_i_decode_stage_dp_reg_a_D_I_11_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_11_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_11_port, 
                           QN => n_1700);
   datapath_i_decode_stage_dp_reg_a_D_I_10_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_10_port, CK 
                           => CLK, RN => RST, Q => datapath_i_val_a_i_10_port, 
                           QN => n_1701);
   datapath_i_decode_stage_dp_reg_a_D_I_9_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_9_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_9_port, QN 
                           => n_1702);
   datapath_i_decode_stage_dp_reg_a_D_I_8_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_8_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_8_port, QN 
                           => n_1703);
   datapath_i_decode_stage_dp_reg_a_D_I_7_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_7_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_7_port, QN 
                           => n_1704);
   datapath_i_decode_stage_dp_reg_a_D_I_6_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_6_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_6_port, QN 
                           => n_1705);
   datapath_i_decode_stage_dp_reg_a_D_I_5_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_5_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_5_port, QN 
                           => n_1706);
   datapath_i_decode_stage_dp_reg_a_D_I_4_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_4_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_4_port, QN 
                           => n_1707);
   datapath_i_decode_stage_dp_reg_a_D_I_3_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_3_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_3_port, QN 
                           => n_1708);
   datapath_i_decode_stage_dp_reg_a_D_I_2_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_2_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_2_port, QN 
                           => n_1709);
   datapath_i_decode_stage_dp_reg_a_D_I_1_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_1_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_1_port, QN 
                           => n_1710);
   datapath_i_decode_stage_dp_reg_a_D_I_0_Q_reg : DFFR_X1 port map( D => 
                           datapath_i_decode_stage_dp_val_reg_a_i_0_port, CK =>
                           CLK, RN => RST, Q => datapath_i_val_a_i_0_port, QN 
                           => n_1711);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           QN => n_1712);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           QN => n_1713);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           QN => n_1714);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           QN => n_1715);
   datapath_i_decode_stage_dp_delay_reg_wb_3_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_2_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           QN => n_1716);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_4_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_4_port, QN 
                           => n_1717);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_3_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_3_port, QN 
                           => n_1718);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_2_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_2_port, QN 
                           => n_1719);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_1_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_1_port, QN 
                           => n_1720);
   datapath_i_decode_stage_dp_delay_reg_wb_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_del_reg_wb_1_0_port, 
                           CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_2_0_port, QN 
                           => n_1721);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => n1926, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_4_port, QN 
                           => n_1722);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => n1927, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_3_port, QN 
                           => n_1723);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_n78, CK => CLK, RN => 
                           RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_2_port, QN 
                           => n_1724);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => n1928, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_1_port, QN 
                           => n_1725);
   datapath_i_decode_stage_dp_delay_reg_wb_1_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => n1929, CK => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_del_reg_wb_1_0_port, QN 
                           => n_1726);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n69, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_31_port, QN => 
                           n2316);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n68, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_30_port, QN => 
                           n2304);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n67, CK => CLK, RN => 
                           RST, Q => n2315, QN => n737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n66, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_28_port, QN => 
                           n2307);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n65, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_27_port, QN => 
                           n2305);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n64, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_26_port, QN => 
                           n2302);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n63, CK => CLK, RN => 
                           RST, Q => datapath_i_n9, QN => n_1727);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n62, CK => CLK, RN => 
                           RST, Q => datapath_i_n10, QN => n_1728);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n61, CK => CLK, RN => 
                           RST, Q => datapath_i_n11, QN => n_1729);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n60, CK => CLK, RN => 
                           RST, Q => datapath_i_n12, QN => n_1730);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n59, CK => CLK, RN => 
                           RST, Q => datapath_i_n13, QN => n_1731);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n58, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_20_port, QN => 
                           n_1732);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n57, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_19_port, QN => 
                           n_1733);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n56, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_18_port, QN => 
                           n697);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n55, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_17_port, QN => 
                           n_1734);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n54, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_16_port, QN => 
                           n_1735);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n53, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_15_port, QN => 
                           n_1736);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n52, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_14_port, QN => 
                           n_1737);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n51, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_13_port, QN => 
                           n740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n50, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_12_port, QN => 
                           n_1738);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n49, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_11_port, QN => 
                           n_1739);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_fetch_stage_dp_n48, CK => CLK, RN => 
                           RST, Q => datapath_i_n14, QN => n_1740);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n47, CK => CLK, RN => 
                           RST, Q => datapath_i_n15, QN => n_1741);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n46, CK => CLK, RN => 
                           RST, Q => datapath_i_n16, QN => n_1742);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n45, CK => CLK, RN => 
                           RST, Q => datapath_i_n17, QN => n_1743);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n44, CK => CLK, RN => 
                           RST, Q => datapath_i_n18, QN => n_1744);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n43, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_5_port, QN => 
                           n2310);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n42, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_4_port, QN => 
                           n_1745);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n41, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_3_port, QN => 
                           n2311);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n40, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_2_port, QN => 
                           n_1746);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n39, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_1_port, QN => 
                           n2301);
   datapath_i_fetch_stage_dp_instruction_reg_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_n38, CK => CLK, RN => 
                           RST, Q => curr_instruction_to_cu_i_0_port, QN => 
                           n2309);
   datapath_i_fetch_stage_dp_new_program_counter_D_I_31_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n2, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_31_port, QN => n_1747
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_30_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n3, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_30_port, QN => n_1748
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_29_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n4, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_29_port, QN => n_1749
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_28_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n9, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_28_port, QN => n_1750
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_27_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n10, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_27_port, QN => n_1751
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_26_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n11, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_26_port, QN => n_1752
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_25_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n12, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_25_port, QN => n_1753
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_24_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n13, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_24_port, QN => n_1754
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_23_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n14, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_23_port, QN => n_1755
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_22_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n15, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_22_port, QN => n_1756
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_21_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n16, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_21_port, QN => n_1757
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_20_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n17, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_20_port, QN => n_1758
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_19_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n18, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_19_port, QN => n_1759
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_18_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n19, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_18_port, QN => n_1760
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_17_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n20, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_17_port, QN => n_1761
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_16_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n21, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_16_port, QN => n_1762
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_15_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n22, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_15_port, QN => n_1763
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_14_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n23, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_14_port, QN => n_1764
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_13_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n24, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_13_port, QN => n_1765
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_12_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n25, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_12_port, QN => n_1766
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_11_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n26, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_11_port, QN => n_1767
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_10_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n27, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_10_port, QN => n_1768
                           );
   datapath_i_fetch_stage_dp_new_program_counter_D_I_9_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n28, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_9_port, QN => n_1769)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_8_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n29, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_8_port, QN => n_1770)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_7_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n30, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_7_port, QN => n_1771)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_6_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n31, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_6_port, QN => n_1772)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_5_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n32, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_5_port, QN => n_1773)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_4_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n33, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_4_port, QN => n_1774)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_3_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n34, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_3_port, QN => n_1775)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_2_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n35, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_2_port, QN => n_1776)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_1_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n36, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_1_port, QN => n_1777)
                           ;
   datapath_i_fetch_stage_dp_new_program_counter_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => datapath_i_fetch_stage_dp_n37, CK => CLK, 
                           RN => RST, Q => 
                           datapath_i_new_pc_value_decode_0_port, QN => n_1778)
                           ;
   datapath_i_fetch_stage_dp_program_counter_D_I_31_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_31_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_31_port, QN => 
                           n_1779);
   datapath_i_fetch_stage_dp_program_counter_D_I_30_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_30_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_30_port, QN => 
                           n_1780);
   datapath_i_fetch_stage_dp_program_counter_D_I_29_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_29_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_29_port, QN => 
                           n753);
   datapath_i_fetch_stage_dp_program_counter_D_I_28_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_28_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_28_port, QN => 
                           n_1781);
   datapath_i_fetch_stage_dp_program_counter_D_I_27_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_27_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_27_port, QN => 
                           n751);
   datapath_i_fetch_stage_dp_program_counter_D_I_26_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_26_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_26_port, QN => 
                           n_1782);
   datapath_i_fetch_stage_dp_program_counter_D_I_25_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_25_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_25_port, QN => 
                           n750);
   datapath_i_fetch_stage_dp_program_counter_D_I_24_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_24_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_24_port, QN => 
                           n_1783);
   datapath_i_fetch_stage_dp_program_counter_D_I_23_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_23_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_23_port, QN => 
                           n749);
   datapath_i_fetch_stage_dp_program_counter_D_I_22_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_22_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_22_port, QN => 
                           n_1784);
   datapath_i_fetch_stage_dp_program_counter_D_I_21_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_21_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_21_port, QN => 
                           n748);
   datapath_i_fetch_stage_dp_program_counter_D_I_20_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_20_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_20_port, QN => 
                           n_1785);
   datapath_i_fetch_stage_dp_program_counter_D_I_19_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_19_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_19_port, QN => 
                           n747);
   datapath_i_fetch_stage_dp_program_counter_D_I_18_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_18_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_18_port, QN => 
                           n_1786);
   datapath_i_fetch_stage_dp_program_counter_D_I_17_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_17_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_17_port, QN => 
                           n746);
   datapath_i_fetch_stage_dp_program_counter_D_I_16_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_16_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_16_port, QN => 
                           n_1787);
   datapath_i_fetch_stage_dp_program_counter_D_I_15_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_15_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_15_port, QN => 
                           n745);
   datapath_i_fetch_stage_dp_program_counter_D_I_14_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_14_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_14_port, QN => 
                           n_1788);
   datapath_i_fetch_stage_dp_program_counter_D_I_13_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_13_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_13_port, QN => 
                           n752);
   datapath_i_fetch_stage_dp_program_counter_D_I_12_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_12_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_12_port, QN => 
                           n_1789);
   datapath_i_fetch_stage_dp_program_counter_D_I_11_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_11_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_11_port, QN => 
                           n744);
   datapath_i_fetch_stage_dp_program_counter_D_I_10_Q_reg : DFFR_X1 port map( D
                           => datapath_i_new_pc_value_mem_stage_i_10_port, CK 
                           => CLK, RN => RST, Q => IRAM_ADDRESS_10_port, QN => 
                           n_1790);
   datapath_i_fetch_stage_dp_program_counter_D_I_9_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_9_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_9_port, QN => n743
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_8_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_8_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_8_port, QN => 
                           n_1791);
   datapath_i_fetch_stage_dp_program_counter_D_I_7_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_7_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_7_port, QN => n742
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_6_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_6_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_6_port, QN => 
                           n_1792);
   datapath_i_fetch_stage_dp_program_counter_D_I_5_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_5_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_5_port, QN => n741
                           );
   datapath_i_fetch_stage_dp_program_counter_D_I_4_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_4_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_4_port, QN => 
                           n_1793);
   datapath_i_fetch_stage_dp_program_counter_D_I_3_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_3_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_3_port, QN => 
                           n_1794);
   datapath_i_fetch_stage_dp_program_counter_D_I_2_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_new_pc_value_mem_stage_i_2_port, CK =>
                           CLK, RN => RST, Q => IRAM_ADDRESS_2_port, QN => 
                           n_1795);
   datapath_i_fetch_stage_dp_program_counter_D_I_1_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N6, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N40_port, QN => 
                           n_1796);
   datapath_i_fetch_stage_dp_program_counter_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_fetch_stage_dp_N5, CK => CLK, RN => 
                           RST, Q => datapath_i_fetch_stage_dp_N39_port, QN => 
                           n_1797);
   cu_i_cmd_alu_op_type_reg_0_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N264, Q => cu_i_cmd_alu_op_type_0_port);
   datapath_i_execute_stage_dp_condition_delay_reg_D_I_0_Q_reg : DFFR_X1 port 
                           map( D => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port, 
                           CK => CLK, RN => RST, Q => n2306, QN => n1534);
   datapath_i_decode_stage_dp_pc_delay_reg_2_D_I_0_Q_reg : DFFR_X1 port map( D 
                           => datapath_i_decode_stage_dp_pc_delay2_0_port, CK 
                           => CLK, RN => RST, Q => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, QN => 
                           n_1798);
   cu_i_cmd_alu_op_type_reg_1_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N265, Q => cu_i_cmd_alu_op_type_1_port);
   cu_i_counter_mul_reg_1_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_1_port, CK => CLK, RN => 
                           RST, Q => n2312, QN => cu_i_n26);
   U1922 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(9), ZN => 
                           datapath_i_memory_stage_dp_data_ir_9_port);
   U1923 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(8), ZN => 
                           datapath_i_memory_stage_dp_data_ir_8_port);
   U1924 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(7), ZN => 
                           datapath_i_memory_stage_dp_data_ir_7_port);
   U1925 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(6), ZN => 
                           datapath_i_memory_stage_dp_data_ir_6_port);
   U1926 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(5), ZN => 
                           datapath_i_memory_stage_dp_data_ir_5_port);
   U1927 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(4), ZN => 
                           datapath_i_memory_stage_dp_data_ir_4_port);
   U1928 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(3), ZN => 
                           datapath_i_memory_stage_dp_data_ir_3_port);
   U1929 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(31), ZN => 
                           datapath_i_memory_stage_dp_data_ir_31_port);
   U1930 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(30), ZN => 
                           datapath_i_memory_stage_dp_data_ir_30_port);
   U1931 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(2), ZN => 
                           datapath_i_memory_stage_dp_data_ir_2_port);
   U1932 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(29), ZN => 
                           datapath_i_memory_stage_dp_data_ir_29_port);
   U1933 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(28), ZN => 
                           datapath_i_memory_stage_dp_data_ir_28_port);
   U1934 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(27), ZN => 
                           datapath_i_memory_stage_dp_data_ir_27_port);
   U1935 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(26), ZN => 
                           datapath_i_memory_stage_dp_data_ir_26_port);
   U1936 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(25), ZN => 
                           datapath_i_memory_stage_dp_data_ir_25_port);
   U1937 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(24), ZN => 
                           datapath_i_memory_stage_dp_data_ir_24_port);
   U1938 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(23), ZN => 
                           datapath_i_memory_stage_dp_data_ir_23_port);
   U1939 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(22), ZN => 
                           datapath_i_memory_stage_dp_data_ir_22_port);
   U1940 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(21), ZN => 
                           datapath_i_memory_stage_dp_data_ir_21_port);
   U1941 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(20), ZN => 
                           datapath_i_memory_stage_dp_data_ir_20_port);
   U1942 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(1), ZN => 
                           datapath_i_memory_stage_dp_data_ir_1_port);
   U1943 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(19), ZN => 
                           datapath_i_memory_stage_dp_data_ir_19_port);
   U1944 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(18), ZN => 
                           datapath_i_memory_stage_dp_data_ir_18_port);
   U1945 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(17), ZN => 
                           datapath_i_memory_stage_dp_data_ir_17_port);
   U1946 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(16), ZN => 
                           datapath_i_memory_stage_dp_data_ir_16_port);
   U1947 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(15), ZN => 
                           datapath_i_memory_stage_dp_data_ir_15_port);
   U1948 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(14), ZN => 
                           datapath_i_memory_stage_dp_data_ir_14_port);
   U1949 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(13), ZN => 
                           datapath_i_memory_stage_dp_data_ir_13_port);
   U1950 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(12), ZN => 
                           datapath_i_memory_stage_dp_data_ir_12_port);
   U1951 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(11), ZN => 
                           datapath_i_memory_stage_dp_data_ir_11_port);
   U1952 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(10), ZN => 
                           datapath_i_memory_stage_dp_data_ir_10_port);
   U1953 : AND2_X1 port map( A1 => DRAM_READY, A2 => DRAM_DATA(0), ZN => 
                           datapath_i_memory_stage_dp_data_ir_0_port);
   cu_i_cmd_alu_op_type_reg_2_inst : DLH_X1 port map( G => cu_i_N278, D => 
                           cu_i_N266, Q => cu_i_cmd_alu_op_type_2_port);
   cu_i_counter_mul_reg_2_inst : DFFR_X1 port map( D => 
                           cu_i_next_val_counter_mul_2_port, CK => CLK, RN => 
                           RST, Q => n2317, QN => cu_i_n25);
   cu_i_curr_state_reg_0_inst : DFFS_X1 port map( D => cu_i_n210, CK => CLK, SN
                           => RST, Q => n2314, QN => cu_i_n23);
   cu_i_stall_reg : DFFR_X2 port map( D => cu_i_next_stall, CK => CLK, RN => 
                           RST, Q => n704, QN => n2308);
   U1954 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           curr_instruction_to_cu_i_28_port, A3 => 
                           curr_instruction_to_cu_i_30_port, A4 => n2015, ZN =>
                           n2074);
   U1955 : AOI21_X1 port map( B1 => n2192, B2 => n2191, A => cu_i_cw3_6_port, 
                           ZN => n2193);
   U1956 : CLKBUF_X1 port map( A => n2228, Z => n2219);
   U1957 : OAI21_X1 port map( B1 => n2059, B2 => n2060, A => n699, ZN => 
                           write_rf_i);
   U1958 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_0_port, B1
                           => cu_i_cw1_0_port, B2 => n2308, ZN => n2021);
   U1959 : NAND2_X1 port map( A1 => cu_i_n25, A2 => cu_i_n26, ZN => n1964);
   U1960 : OR2_X1 port map( A1 => enable_rf_i, A2 => write_rf_i, ZN => 
                           datapath_i_decode_stage_dp_enable_rf_i);
   U1961 : NAND2_X1 port map( A1 => n1964, A2 => n2313, ZN => n2059);
   U1962 : NOR2_X1 port map( A1 => cu_i_n123, A2 => n2314, ZN => n2064);
   U1963 : CLKBUF_X1 port map( A => n2138, Z => n2186);
   U1964 : AOI21_X1 port map( B1 => n2008, B2 => n2017, A => n2066, ZN => n2189
                           );
   U1965 : NOR3_X1 port map( A1 => n2301, A2 => n2309, A3 => n1965, ZN => n2017
                           );
   U1966 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           curr_instruction_to_cu_i_30_port, A3 => n1933, ZN =>
                           cu_i_cmd_word_4_port);
   U1967 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           curr_instruction_to_cu_i_31_port, A3 => n2064, A4 =>
                           curr_instruction_to_cu_i_26_port, ZN => n1933);
   U1968 : OAI22_X1 port map( A1 => n2308, A2 => cu_i_cmd_word_4_port, B1 => 
                           cu_i_cw2_8_port, B2 => n704, ZN => n309);
   U1969 : INV_X1 port map( A => n309, ZN => DRAM_ENABLE_port);
   U1970 : INV_X1 port map( A => cu_i_cmd_word_4_port, ZN => n2187);
   U1971 : NOR2_X1 port map( A1 => n2315, A2 => n2187, ZN => 
                           cu_i_cmd_word_3_port);
   U1972 : OAI22_X1 port map( A1 => n2308, A2 => cu_i_cmd_word_3_port, B1 => 
                           cu_i_cw2_7_port, B2 => n704, ZN => n2019);
   U1973 : NAND2_X1 port map( A1 => DRAM_ENABLE_port, A2 => n2019, ZN => 
                           datapath_i_memory_stage_dp_n2);
   U1974 : CLKBUF_X1 port map( A => datapath_i_memory_stage_dp_n2, Z => n2323);
   U1975 : INV_X1 port map( A => DRAM_ENABLE_port, ZN => n2321);
   U1976 : NAND2_X2 port map( A1 => n1534, A2 => 
                           datapath_i_decode_stage_dp_pc_delay3_0_port, ZN => 
                           n2180);
   U1977 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n2306, ZN => n2178);
   U1978 : CLKBUF_X1 port map( A => n2306, Z => n2177);
   U1979 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_29_port,
                           B2 => n2177, ZN => n1934);
   U1980 : OAI21_X1 port map( B1 => n726, B2 => n2180, A => n1934, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_29_port);
   U1981 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_27_port,
                           B2 => n2177, ZN => n1935);
   U1982 : OAI21_X1 port map( B1 => n724, B2 => n2180, A => n1935, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_27_port);
   U1983 : CLKBUF_X1 port map( A => n2178, Z => n1959);
   U1984 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_25_port,
                           B2 => n2306, ZN => n1936);
   U1985 : OAI21_X1 port map( B1 => n723, B2 => n2180, A => n1936, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_25_port);
   U1986 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_23_port,
                           B2 => n2306, ZN => n1937);
   U1987 : OAI21_X1 port map( B1 => n721, B2 => n2180, A => n1937, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_23_port);
   U1988 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_21_port,
                           B2 => n2306, ZN => n1938);
   U1989 : OAI21_X1 port map( B1 => n719, B2 => n2180, A => n1938, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_21_port);
   U1990 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_19_port,
                           B2 => n2306, ZN => n1939);
   U1991 : OAI21_X1 port map( B1 => n717, B2 => n2180, A => n1939, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_19_port);
   U1992 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_17_port,
                           B2 => n2306, ZN => n1940);
   U1993 : OAI21_X1 port map( B1 => n715, B2 => n2180, A => n1940, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_17_port);
   U1994 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_15_port,
                           B2 => n2306, ZN => n1941);
   U1995 : OAI21_X1 port map( B1 => n713, B2 => n2180, A => n1941, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_15_port);
   U1996 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_13_port,
                           B2 => n2306, ZN => n1942);
   U1997 : OAI21_X1 port map( B1 => n711, B2 => n2180, A => n1942, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_13_port);
   U1998 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_11_port,
                           B2 => n2177, ZN => n1943);
   U1999 : OAI21_X1 port map( B1 => n709, B2 => n2180, A => n1943, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_11_port);
   U2000 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_9_port, 
                           B2 => n2177, ZN => n1944);
   U2001 : OAI21_X1 port map( B1 => n707, B2 => n2180, A => n1944, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_9_port);
   U2002 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_7_port, 
                           B2 => n2177, ZN => n1945);
   U2003 : OAI21_X1 port map( B1 => n705, B2 => n2180, A => n1945, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_7_port);
   U2004 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_5_port, 
                           B2 => n2177, ZN => n1946);
   U2005 : OAI21_X1 port map( B1 => n731, B2 => n2180, A => n1946, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_5_port);
   U2006 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_4_port, 
                           B2 => n2306, ZN => n1947);
   U2007 : OAI21_X1 port map( B1 => n730, B2 => n2180, A => n1947, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_4_port);
   U2008 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_2_port, 
                           B2 => n2177, ZN => n1948);
   U2009 : OAI21_X1 port map( B1 => n728, B2 => n2180, A => n1948, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_2_port);
   U2010 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_3_port, 
                           B2 => n2306, ZN => n1949);
   U2011 : OAI21_X1 port map( B1 => n729, B2 => n2180, A => n1949, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_3_port);
   U2012 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_6_port, 
                           B2 => n2306, ZN => n1950);
   U2013 : OAI21_X1 port map( B1 => n732, B2 => n2180, A => n1950, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_6_port);
   U2014 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_8_port, 
                           B2 => n2306, ZN => n1951);
   U2015 : OAI21_X1 port map( B1 => n706, B2 => n2180, A => n1951, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_8_port);
   U2016 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_10_port,
                           B2 => n2306, ZN => n1952);
   U2017 : OAI21_X1 port map( B1 => n708, B2 => n2180, A => n1952, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_10_port);
   U2018 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_12_port,
                           B2 => n2177, ZN => n1953);
   U2019 : OAI21_X1 port map( B1 => n710, B2 => n2180, A => n1953, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_12_port);
   U2020 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_14_port,
                           B2 => n2177, ZN => n1954);
   U2021 : OAI21_X1 port map( B1 => n712, B2 => n2180, A => n1954, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_14_port);
   U2022 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_16_port,
                           B2 => n2177, ZN => n1955);
   U2023 : OAI21_X1 port map( B1 => n714, B2 => n2180, A => n1955, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_16_port);
   U2024 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_18_port,
                           B2 => n2306, ZN => n1956);
   U2025 : OAI21_X1 port map( B1 => n716, B2 => n2180, A => n1956, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_18_port);
   U2026 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_20_port,
                           B2 => n2306, ZN => n1957);
   U2027 : OAI21_X1 port map( B1 => n718, B2 => n2180, A => n1957, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_20_port);
   U2028 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_22_port,
                           B2 => n2306, ZN => n1958);
   U2029 : OAI21_X1 port map( B1 => n720, B2 => n2180, A => n1958, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_22_port);
   U2030 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n1959, B1 => datapath_i_alu_output_val_i_24_port,
                           B2 => n2177, ZN => n1960);
   U2031 : OAI21_X1 port map( B1 => n722, B2 => n2180, A => n1960, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_24_port);
   U2032 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_26_port,
                           B2 => n2177, ZN => n1961);
   U2033 : OAI21_X1 port map( B1 => n691, B2 => n2180, A => n1961, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_26_port);
   U2034 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_28_port,
                           B2 => n2177, ZN => n1962);
   U2035 : OAI21_X1 port map( B1 => n725, B2 => n2180, A => n1962, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_28_port);
   U2036 : NAND4_X1 port map( A1 => n737, A2 => n2064, A3 => n2316, A4 => n2304
                           , ZN => n1963);
   U2037 : OR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n2305
                           , A3 => n1963, ZN => n2232);
   U2038 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n2305, ZN => n2051);
   U2039 : OR2_X1 port map( A1 => n1963, A2 => n2051, ZN => n2233);
   U2040 : NAND2_X1 port map( A1 => n2232, A2 => n2233, ZN => n1152);
   U2041 : NAND4_X1 port map( A1 => cu_i_n26, A2 => cu_i_n25, A3 => n2303, A4 
                           => n2313, ZN => cu_i_n145);
   U2042 : NAND2_X1 port map( A1 => cu_i_n145, A2 => n2059, ZN => n2008);
   U2043 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           curr_instruction_to_cu_i_2_port, A3 => 
                           curr_instruction_to_cu_i_5_port, A4 => 
                           curr_instruction_to_cu_i_4_port, ZN => n1965);
   U2044 : NAND3_X1 port map( A1 => n737, A2 => n2316, A3 => n2302, ZN => n2015
                           );
   U2045 : NAND2_X1 port map( A1 => n2017, A2 => n2074, ZN => n2034);
   U2046 : OAI21_X1 port map( B1 => n2008, B2 => n2034, A => n2064, ZN => n1966
                           );
   U2047 : NAND2_X1 port map( A1 => cu_i_n123, A2 => n2314, ZN => n2078);
   U2048 : AOI21_X1 port map( B1 => n1966, B2 => n2078, A => n704, ZN => 
                           IRAM_ENABLE_port);
   U2049 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_29_port, 
                           ZN => n1967);
   U2050 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_27_port, 
                           ZN => n1970);
   U2051 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_25_port, 
                           ZN => n1973);
   U2052 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_23_port, 
                           ZN => n1976);
   U2053 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_21_port, 
                           ZN => n1979);
   U2054 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_19_port, 
                           ZN => n1982);
   U2055 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_17_port, 
                           ZN => n1985);
   U2056 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_15_port, 
                           ZN => n1988);
   U2057 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_13_port, 
                           ZN => n1991);
   U2058 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_11_port, 
                           ZN => n1994);
   U2059 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_9_port, ZN
                           => n1997);
   U2060 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_7_port, ZN
                           => n2000);
   U2061 : INV_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_5_port, ZN
                           => n2003);
   U2062 : NAND3_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_4_port,
                           A2 => datapath_i_new_pc_value_mem_stage_i_2_port, A3
                           => datapath_i_new_pc_value_mem_stage_i_3_port, ZN =>
                           n2093);
   U2063 : NOR2_X1 port map( A1 => n2003, A2 => n2093, ZN => n2100);
   U2064 : NAND2_X1 port map( A1 => n2100, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, ZN => 
                           n2099);
   U2065 : NOR2_X1 port map( A1 => n2000, A2 => n2099, ZN => n2106);
   U2066 : NAND2_X1 port map( A1 => n2106, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, ZN => 
                           n2105);
   U2067 : NOR2_X1 port map( A1 => n1997, A2 => n2105, ZN => n2112);
   U2068 : NAND2_X1 port map( A1 => n2112, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, ZN => 
                           n2111);
   U2069 : NOR2_X1 port map( A1 => n1994, A2 => n2111, ZN => n2118);
   U2070 : NAND2_X1 port map( A1 => n2118, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, ZN => 
                           n2117);
   U2071 : NOR2_X1 port map( A1 => n1991, A2 => n2117, ZN => n2124);
   U2072 : NAND2_X1 port map( A1 => n2124, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, ZN => 
                           n2123);
   U2073 : NOR2_X1 port map( A1 => n1988, A2 => n2123, ZN => n2130);
   U2074 : NAND2_X1 port map( A1 => n2130, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, ZN => 
                           n2129);
   U2075 : NOR2_X1 port map( A1 => n1985, A2 => n2129, ZN => n2136);
   U2076 : NAND2_X1 port map( A1 => n2136, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, ZN => 
                           n2135);
   U2077 : NOR2_X1 port map( A1 => n1982, A2 => n2135, ZN => n2143);
   U2078 : NAND2_X1 port map( A1 => n2143, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, ZN => 
                           n2142);
   U2079 : NOR2_X1 port map( A1 => n1979, A2 => n2142, ZN => n2149);
   U2080 : NAND2_X1 port map( A1 => n2149, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, ZN => 
                           n2148);
   U2081 : NOR2_X1 port map( A1 => n1976, A2 => n2148, ZN => n2155);
   U2082 : NAND2_X1 port map( A1 => n2155, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, ZN => 
                           n2154);
   U2083 : NOR2_X1 port map( A1 => n1973, A2 => n2154, ZN => n2161);
   U2084 : NAND2_X1 port map( A1 => n2161, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, ZN => 
                           n2160);
   U2085 : NOR2_X1 port map( A1 => n1970, A2 => n2160, ZN => n2167);
   U2086 : NAND2_X1 port map( A1 => n2167, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, ZN => 
                           n2166);
   U2087 : INV_X1 port map( A => n1152, ZN => n2079);
   U2088 : OAI221_X1 port map( B1 => n2308, B2 => n2079, C1 => n704, C2 => n756
                           , A => n1534, ZN => n2090);
   U2089 : INV_X1 port map( A => n2090, ZN => n2138);
   U2090 : NOR2_X1 port map( A1 => n1967, A2 => n2166, ZN => n2173);
   U2091 : AOI211_X1 port map( C1 => n1967, C2 => n2166, A => n2138, B => n2173
                           , ZN => n1969);
   U2092 : NAND2_X1 port map( A1 => IRAM_ENABLE_port, A2 => IRAM_ADDRESS_2_port
                           , ZN => n2087);
   U2093 : INV_X1 port map( A => n2087, ZN => n2089);
   U2094 : AND2_X1 port map( A1 => n2089, A2 => IRAM_ADDRESS_3_port, ZN => 
                           n2096);
   U2095 : NAND2_X1 port map( A1 => n2096, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n2095);
   U2096 : NOR2_X1 port map( A1 => n741, A2 => n2095, ZN => n2102);
   U2097 : NAND2_X1 port map( A1 => n2102, A2 => IRAM_ADDRESS_6_port, ZN => 
                           n2101);
   U2098 : NOR2_X1 port map( A1 => n742, A2 => n2101, ZN => n2108);
   U2099 : NAND2_X1 port map( A1 => n2108, A2 => IRAM_ADDRESS_8_port, ZN => 
                           n2107);
   U2100 : NOR2_X1 port map( A1 => n743, A2 => n2107, ZN => n2114);
   U2101 : NAND2_X1 port map( A1 => n2114, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n2113);
   U2102 : NOR2_X1 port map( A1 => n744, A2 => n2113, ZN => n2120);
   U2103 : NAND2_X1 port map( A1 => n2120, A2 => IRAM_ADDRESS_12_port, ZN => 
                           n2119);
   U2104 : NOR2_X1 port map( A1 => n752, A2 => n2119, ZN => n2126);
   U2105 : NAND2_X1 port map( A1 => n2126, A2 => IRAM_ADDRESS_14_port, ZN => 
                           n2125);
   U2106 : NOR2_X1 port map( A1 => n745, A2 => n2125, ZN => n2132);
   U2107 : NAND2_X1 port map( A1 => n2132, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n2131);
   U2108 : NOR2_X1 port map( A1 => n746, A2 => n2131, ZN => n2139);
   U2109 : NAND2_X1 port map( A1 => n2139, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n2137);
   U2110 : NOR2_X1 port map( A1 => n747, A2 => n2137, ZN => n2145);
   U2111 : NAND2_X1 port map( A1 => n2145, A2 => IRAM_ADDRESS_20_port, ZN => 
                           n2144);
   U2112 : NOR2_X1 port map( A1 => n748, A2 => n2144, ZN => n2151);
   U2113 : NAND2_X1 port map( A1 => n2151, A2 => IRAM_ADDRESS_22_port, ZN => 
                           n2150);
   U2114 : NOR2_X1 port map( A1 => n749, A2 => n2150, ZN => n2157);
   U2115 : NAND2_X1 port map( A1 => n2157, A2 => IRAM_ADDRESS_24_port, ZN => 
                           n2156);
   U2116 : NOR2_X1 port map( A1 => n750, A2 => n2156, ZN => n2163);
   U2117 : NAND2_X1 port map( A1 => n2163, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n2162);
   U2118 : NOR2_X1 port map( A1 => n751, A2 => n2162, ZN => n2169);
   U2119 : NAND2_X1 port map( A1 => n2169, A2 => IRAM_ADDRESS_28_port, ZN => 
                           n2168);
   U2120 : NOR2_X1 port map( A1 => n753, A2 => n2168, ZN => n2174);
   U2121 : INV_X1 port map( A => n2186, ZN => n2183);
   U2122 : AOI211_X1 port map( C1 => n753, C2 => n2168, A => n2174, B => n2183,
                           ZN => n1968);
   U2123 : OR2_X1 port map( A1 => n1969, A2 => n1968, ZN => 
                           datapath_i_fetch_stage_dp_n4);
   U2124 : AOI211_X1 port map( C1 => n1970, C2 => n2160, A => n2138, B => n2167
                           , ZN => n1972);
   U2125 : AOI211_X1 port map( C1 => n751, C2 => n2162, A => n2169, B => n2090,
                           ZN => n1971);
   U2126 : OR2_X1 port map( A1 => n1972, A2 => n1971, ZN => 
                           datapath_i_fetch_stage_dp_n10);
   U2127 : AOI211_X1 port map( C1 => n1973, C2 => n2154, A => n2138, B => n2161
                           , ZN => n1975);
   U2128 : AOI211_X1 port map( C1 => n750, C2 => n2156, A => n2163, B => n2183,
                           ZN => n1974);
   U2129 : OR2_X1 port map( A1 => n1975, A2 => n1974, ZN => 
                           datapath_i_fetch_stage_dp_n12);
   U2130 : AOI211_X1 port map( C1 => n1976, C2 => n2148, A => n2186, B => n2155
                           , ZN => n1978);
   U2131 : AOI211_X1 port map( C1 => n749, C2 => n2150, A => n2157, B => n2183,
                           ZN => n1977);
   U2132 : OR2_X1 port map( A1 => n1978, A2 => n1977, ZN => 
                           datapath_i_fetch_stage_dp_n14);
   U2133 : AOI211_X1 port map( C1 => n1979, C2 => n2142, A => n2186, B => n2149
                           , ZN => n1981);
   U2134 : AOI211_X1 port map( C1 => n748, C2 => n2144, A => n2151, B => n2090,
                           ZN => n1980);
   U2135 : OR2_X1 port map( A1 => n1981, A2 => n1980, ZN => 
                           datapath_i_fetch_stage_dp_n16);
   U2136 : AOI211_X1 port map( C1 => n1982, C2 => n2135, A => n2186, B => n2143
                           , ZN => n1984);
   U2137 : AOI211_X1 port map( C1 => n747, C2 => n2137, A => n2145, B => n2090,
                           ZN => n1983);
   U2138 : OR2_X1 port map( A1 => n1984, A2 => n1983, ZN => 
                           datapath_i_fetch_stage_dp_n18);
   U2139 : AOI211_X1 port map( C1 => n1985, C2 => n2129, A => n2138, B => n2136
                           , ZN => n1987);
   U2140 : AOI211_X1 port map( C1 => n746, C2 => n2131, A => n2139, B => n2090,
                           ZN => n1986);
   U2141 : OR2_X1 port map( A1 => n1987, A2 => n1986, ZN => 
                           datapath_i_fetch_stage_dp_n20);
   U2142 : AOI211_X1 port map( C1 => n1988, C2 => n2123, A => n2138, B => n2130
                           , ZN => n1990);
   U2143 : AOI211_X1 port map( C1 => n745, C2 => n2125, A => n2132, B => n2183,
                           ZN => n1989);
   U2144 : OR2_X1 port map( A1 => n1990, A2 => n1989, ZN => 
                           datapath_i_fetch_stage_dp_n22);
   U2145 : AOI211_X1 port map( C1 => n1991, C2 => n2117, A => n2138, B => n2124
                           , ZN => n1993);
   U2146 : AOI211_X1 port map( C1 => n752, C2 => n2119, A => n2126, B => n2183,
                           ZN => n1992);
   U2147 : OR2_X1 port map( A1 => n1993, A2 => n1992, ZN => 
                           datapath_i_fetch_stage_dp_n24);
   U2148 : AOI211_X1 port map( C1 => n1994, C2 => n2111, A => n2138, B => n2118
                           , ZN => n1996);
   U2149 : AOI211_X1 port map( C1 => n744, C2 => n2113, A => n2120, B => n2183,
                           ZN => n1995);
   U2150 : OR2_X1 port map( A1 => n1996, A2 => n1995, ZN => 
                           datapath_i_fetch_stage_dp_n26);
   U2151 : AOI211_X1 port map( C1 => n1997, C2 => n2105, A => n2138, B => n2112
                           , ZN => n1999);
   U2152 : AOI211_X1 port map( C1 => n743, C2 => n2107, A => n2114, B => n2183,
                           ZN => n1998);
   U2153 : OR2_X1 port map( A1 => n1999, A2 => n1998, ZN => 
                           datapath_i_fetch_stage_dp_n28);
   U2154 : AOI211_X1 port map( C1 => n2000, C2 => n2099, A => n2186, B => n2106
                           , ZN => n2002);
   U2155 : AOI211_X1 port map( C1 => n742, C2 => n2101, A => n2108, B => n2090,
                           ZN => n2001);
   U2156 : OR2_X1 port map( A1 => n2002, A2 => n2001, ZN => 
                           datapath_i_fetch_stage_dp_n30);
   U2157 : AOI211_X1 port map( C1 => n2003, C2 => n2093, A => n2138, B => n2100
                           , ZN => n2005);
   U2158 : AOI211_X1 port map( C1 => n741, C2 => n2095, A => n2102, B => n2090,
                           ZN => n2004);
   U2159 : OR2_X1 port map( A1 => n2005, A2 => n2004, ZN => 
                           datapath_i_fetch_stage_dp_n32);
   U2160 : INV_X1 port map( A => n704, ZN => n2084);
   U2161 : OAI22_X1 port map( A1 => n2084, A2 => cu_i_cw3_6_port, B1 => 
                           cu_i_cw2_6_port, B2 => n704, ZN => n2006);
   U2162 : INV_X1 port map( A => n2006, ZN => n1932);
   U2163 : NAND2_X1 port map( A1 => n2064, A2 => n2074, ZN => n2066);
   U2164 : INV_X1 port map( A => n2064, ZN => n2080);
   U2165 : NOR3_X1 port map( A1 => n2307, A2 => n2304, A3 => n2015, ZN => n2045
                           );
   U2166 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_31_port, A2 => n737
                           , ZN => n2043);
   U2167 : NAND2_X1 port map( A1 => n2043, A2 => n2304, ZN => n2050);
   U2168 : AOI21_X1 port map( B1 => curr_instruction_to_cu_i_26_port, B2 => 
                           n2051, A => n2050, ZN => n2007);
   U2169 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_30_port, A2 => 
                           n2043, A3 => n2305, ZN => n2032);
   U2170 : AOI21_X1 port map( B1 => n2307, B2 => n2302, A => n2032, ZN => n2036
                           );
   U2171 : NOR3_X1 port map( A1 => n2045, A2 => n2007, A3 => n2036, ZN => n2071
                           );
   U2172 : OAI222_X1 port map( A1 => n2302, A2 => n2232, B1 => n2066, B2 => 
                           n2017, C1 => n2080, C2 => n2071, ZN => n311);
   U2173 : OR2_X1 port map( A1 => cu_i_cmd_word_3_port, A2 => n311, ZN => 
                           cu_i_cmd_word_1_port);
   U2174 : INV_X1 port map( A => n2232, ZN => n2324);
   U2175 : INV_X1 port map( A => n2189, ZN => n2188);
   U2176 : AOI221_X1 port map( B1 => n2188, B2 => 
                           curr_instruction_to_cu_i_20_port, C1 => n2189, C2 =>
                           curr_instruction_to_cu_i_15_port, A => n2324, ZN => 
                           n2009);
   U2177 : INV_X1 port map( A => n2009, ZN => n1926);
   U2178 : AOI221_X1 port map( B1 => n2188, B2 => 
                           curr_instruction_to_cu_i_19_port, C1 => n2189, C2 =>
                           curr_instruction_to_cu_i_14_port, A => n2324, ZN => 
                           n2010);
   U2179 : INV_X1 port map( A => n2010, ZN => n1927);
   U2180 : AOI221_X1 port map( B1 => n2188, B2 => 
                           curr_instruction_to_cu_i_17_port, C1 => n2189, C2 =>
                           curr_instruction_to_cu_i_12_port, A => n2324, ZN => 
                           n2011);
   U2181 : INV_X1 port map( A => n2011, ZN => n1928);
   U2182 : AOI221_X1 port map( B1 => n2188, B2 => 
                           curr_instruction_to_cu_i_16_port, C1 => n2189, C2 =>
                           curr_instruction_to_cu_i_11_port, A => n2324, ZN => 
                           n2012);
   U2183 : INV_X1 port map( A => n2012, ZN => n1929);
   U2184 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_2_port, B1
                           => cu_i_cw1_2_port, B2 => n2084, ZN => n2025);
   U2185 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_1_port, B1
                           => cu_i_cw1_1_port, B2 => n2308, ZN => n2023);
   U2186 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_alu_op_type_3_port, B1
                           => cu_i_cw1_3_port, B2 => n2308, ZN => n2020);
   U2187 : AOI21_X1 port map( B1 => n2025, B2 => n2023, A => n2020, ZN => n2013
                           );
   U2188 : NOR2_X1 port map( A1 => n2021, A2 => n2013, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_0_port);
   U2189 : INV_X1 port map( A => n2020, ZN => n2024);
   U2190 : OAI211_X1 port map( C1 => n2021, C2 => n2023, A => n2024, B => n2025
                           , ZN => n2014);
   U2191 : INV_X1 port map( A => n2014, ZN => n1925);
   U2192 : NOR2_X1 port map( A1 => n2233, A2 => n2302, ZN => 
                           cu_i_cmd_word_7_port);
   U2193 : OAI21_X1 port map( B1 => n2051, B2 => n2015, A => n2071, ZN => n2069
                           );
   U2194 : AOI211_X1 port map( C1 => n2064, C2 => n2069, A => 
                           cu_i_cmd_word_4_port, B => cu_i_cmd_word_7_port, ZN 
                           => n2018);
   U2195 : NAND2_X1 port map( A1 => n2018, A2 => n2188, ZN => enable_rf_i);
   U2196 : INV_X1 port map( A => n2066, ZN => n2016);
   U2197 : NAND2_X1 port map( A1 => n2017, A2 => n2016, ZN => n2060);
   U2198 : NAND2_X1 port map( A1 => n2018, A2 => n2232, ZN => n310);
   U2199 : INV_X1 port map( A => n310, ZN => n2260);
   U2200 : INV_X1 port map( A => n2260, ZN => n2320);
   U2201 : AND2_X1 port map( A1 => n2320, A2 => CLK, ZN => 
                           datapath_i_decode_stage_dp_clk_immediate);
   U2202 : INV_X1 port map( A => n2019, ZN => DRAM_READNOTWRITE);
   U2203 : OAI22_X1 port map( A1 => n2308, A2 => n2260, B1 => n2319, B2 => n704
                           , ZN => n2261);
   U2204 : CLKBUF_X1 port map( A => n2261, Z => n2263);
   U2205 : MUX2_X1 port map( A => datapath_i_val_b_i_2_port, B => 
                           datapath_i_val_immediate_i_2_port, S => n2263, Z => 
                           datapath_i_execute_stage_dp_opb_2_port);
   U2206 : MUX2_X1 port map( A => datapath_i_val_b_i_0_port, B => 
                           datapath_i_val_immediate_i_0_port, S => n2261, Z => 
                           datapath_i_execute_stage_dp_opb_0_port);
   U2207 : MUX2_X1 port map( A => datapath_i_val_b_i_1_port, B => 
                           datapath_i_val_immediate_i_1_port, S => n2263, Z => 
                           datapath_i_execute_stage_dp_opb_1_port);
   U2208 : AOI21_X1 port map( B1 => n2025, B2 => n2021, A => n2020, ZN => n2022
                           );
   U2209 : NOR2_X1 port map( A1 => n2023, A2 => n2022, ZN => 
                           datapath_i_execute_stage_dp_alu_op_type_i_1_port);
   U2210 : NOR2_X1 port map( A1 => n2025, A2 => n2024, ZN => 
                           datapath_i_execute_stage_dp_n7);
   U2211 : NOR2_X1 port map( A1 => n2303, A2 => n2060, ZN => cu_i_N273);
   U2212 : INV_X1 port map( A => n2060, ZN => n2191);
   U2213 : AOI221_X1 port map( B1 => cu_i_n25, B2 => n2191, C1 => cu_i_n26, C2 
                           => n2191, A => cu_i_N273, ZN => n2026);
   U2214 : INV_X1 port map( A => n2026, ZN => n2029);
   U2215 : NOR2_X1 port map( A1 => cu_i_n125, A2 => n2060, ZN => n2027);
   U2216 : NAND2_X1 port map( A1 => n2027, A2 => n2312, ZN => n2058);
   U2217 : NOR2_X1 port map( A1 => cu_i_n25, A2 => n2058, ZN => n2028);
   U2218 : MUX2_X1 port map( A => n2029, B => n2028, S => cu_i_n124, Z => 
                           cu_i_N277);
   datapath_i_execute_stage_dp_n9 <= '0';
   U2220 : NAND2_X1 port map( A1 => n2260, A2 => n2066, ZN => cu_i_N278);
   U2221 : INV_X1 port map( A => n2074, ZN => n2076);
   U2222 : NAND2_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => 
                           n2311, ZN => n2056);
   U2223 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => 
                           curr_instruction_to_cu_i_4_port, A3 => n2076, A4 => 
                           n2056, ZN => n2044);
   U2224 : AOI21_X1 port map( B1 => n2044, B2 => n2310, A => n2045, ZN => n2054
                           );
   U2225 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => 
                           n2051, A3 => n2050, ZN => n2031);
   U2226 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => n2310
                           , A3 => n2076, ZN => n2049);
   U2227 : NAND3_X1 port map( A1 => curr_instruction_to_cu_i_3_port, A2 => 
                           n2049, A3 => n2301, ZN => n2038);
   U2228 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_2_port, A2 => n2309
                           , A3 => n2038, ZN => n2030);
   U2229 : AOI211_X1 port map( C1 => n2044, C2 => n2301, A => n2031, B => n2030
                           , ZN => n2035);
   U2230 : OR3_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => n2302
                           , A3 => n2032, ZN => n2033);
   U2231 : NAND4_X1 port map( A1 => n2054, A2 => n2035, A3 => n2034, A4 => 
                           n2033, ZN => cu_i_N265);
   U2232 : MUX2_X1 port map( A => datapath_i_val_b_i_3_port, B => 
                           datapath_i_val_immediate_i_3_port, S => n2263, Z => 
                           datapath_i_execute_stage_dp_opb_3_port);
   U2233 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_0_port, A2 => 
                           curr_instruction_to_cu_i_2_port, ZN => n2061);
   U2234 : INV_X1 port map( A => n2036, ZN => n2037);
   U2235 : OAI21_X1 port map( B1 => n2061, B2 => n2038, A => n2037, ZN => 
                           cu_i_N267);
   U2236 : NOR2_X1 port map( A1 => n2308, A2 => n1152, ZN => n2039);
   U2237 : NOR2_X1 port map( A1 => n704, A2 => cu_i_cw1_4_port, ZN => n2068);
   U2238 : NOR2_X1 port map( A1 => n2039, A2 => n2068, ZN => n2040);
   U2239 : NAND2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port
                           , A2 => n2040, ZN => n2300);
   U2240 : CLKBUF_X1 port map( A => n2300, Z => n2289);
   U2241 : INV_X1 port map( A => n2040, ZN => n2285);
   U2242 : NOR2_X1 port map( A1 => datapath_i_decode_stage_dp_pc_delay3_0_port,
                           A2 => n2285, ZN => n2298);
   U2243 : CLKBUF_X1 port map( A => n2298, Z => n2287);
   U2244 : CLKBUF_X1 port map( A => n2285, Z => n2297);
   U2245 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_26_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_26_port, B2 => 
                           n2297, ZN => n2041);
   U2246 : OAI21_X1 port map( B1 => n691, B2 => n2289, A => n2041, ZN => 
                           datapath_i_execute_stage_dp_opa_26_port);
   U2247 : OAI221_X1 port map( B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           curr_instruction_to_cu_i_2_port, C1 => n2301, C2 => 
                           n2311, A => n2049, ZN => n2048);
   U2248 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => 
                           n2051, ZN => n2042);
   U2249 : NOR3_X1 port map( A1 => curr_instruction_to_cu_i_26_port, A2 => 
                           n2305, A3 => n2050, ZN => n2063);
   U2250 : AOI21_X1 port map( B1 => n2043, B2 => n2042, A => n2063, ZN => n2047
                           );
   U2251 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_27_port, A2 => 
                           n2045, B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           n2044, ZN => n2046);
   U2252 : OAI211_X1 port map( C1 => curr_instruction_to_cu_i_0_port, C2 => 
                           n2048, A => n2047, B => n2046, ZN => cu_i_N264);
   U2253 : OAI221_X1 port map( B1 => curr_instruction_to_cu_i_1_port, B2 => 
                           curr_instruction_to_cu_i_0_port, C1 => n2301, C2 => 
                           n2309, A => n2049, ZN => n2055);
   U2254 : NOR2_X1 port map( A1 => n2051, A2 => n2050, ZN => n2052);
   U2255 : AOI22_X1 port map( A1 => curr_instruction_to_cu_i_28_port, A2 => 
                           n2063, B1 => curr_instruction_to_cu_i_26_port, B2 =>
                           n2052, ZN => n2053);
   U2256 : OAI211_X1 port map( C1 => n2056, C2 => n2055, A => n2054, B => n2053
                           , ZN => cu_i_N266);
   U2257 : NAND2_X1 port map( A1 => n704, A2 => n2060, ZN => cu_i_N274);
   U2258 : AOI221_X1 port map( B1 => cu_i_n125, B2 => cu_i_n26, C1 => n2303, C2
                           => n2312, A => n2060, ZN => cu_i_N275);
   U2259 : OAI21_X1 port map( B1 => cu_i_n26, B2 => cu_i_n125, A => n2191, ZN 
                           => n2057);
   U2260 : AOI22_X1 port map( A1 => cu_i_n25, A2 => n2058, B1 => n2057, B2 => 
                           n2317, ZN => cu_i_N276);
   U2261 : INV_X1 port map( A => n2059, ZN => n2192);
   U2262 : AOI211_X1 port map( C1 => n704, C2 => cu_i_n145, A => n2192, B => 
                           n2060, ZN => cu_i_N279);
   U2263 : NOR2_X1 port map( A1 => curr_instruction_to_cu_i_4_port, A2 => n2310
                           , ZN => n2062);
   U2264 : NAND4_X1 port map( A1 => curr_instruction_to_cu_i_1_port, A2 => 
                           n2062, A3 => n2061, A4 => n2311, ZN => n2067);
   U2265 : NAND3_X1 port map( A1 => n2064, A2 => n2063, A3 => n2307, ZN => 
                           n2065);
   U2266 : OAI21_X1 port map( B1 => n2067, B2 => n2066, A => n2065, ZN => 
                           cu_i_cmd_word_8_port);
   U2267 : MUX2_X1 port map( A => cu_i_cmd_word_8_port, B => cu_i_cw1_12_port, 
                           S => n2084, Z => alu_cin_i);
   U2268 : AOI21_X1 port map( B1 => n756, B2 => n704, A => n2068, ZN => 
                           cu_i_cw1_i_4_port);
   U2269 : MUX2_X1 port map( A => cu_i_cw2_7_port, B => cu_i_cw1_7_port, S => 
                           n2308, Z => cu_i_cw1_i_7_port);
   U2270 : MUX2_X1 port map( A => cu_i_cw2_8_port, B => cu_i_cw1_8_port, S => 
                           n2308, Z => cu_i_cw1_i_8_port);
   U2271 : INV_X1 port map( A => n2069, ZN => n2077);
   U2272 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_12_port, A2 => 
                           curr_instruction_to_cu_i_11_port, A3 => 
                           curr_instruction_to_cu_i_15_port, A4 => 
                           curr_instruction_to_cu_i_14_port, ZN => n2070);
   U2273 : NAND2_X1 port map( A1 => n740, A2 => n2070, ZN => n2075);
   U2274 : NOR4_X1 port map( A1 => curr_instruction_to_cu_i_17_port, A2 => 
                           curr_instruction_to_cu_i_16_port, A3 => 
                           curr_instruction_to_cu_i_20_port, A4 => 
                           curr_instruction_to_cu_i_19_port, ZN => n2072);
   U2275 : AOI21_X1 port map( B1 => n697, B2 => n2072, A => n2071, ZN => n2073)
                           ;
   U2276 : AOI221_X1 port map( B1 => n2077, B2 => n2076, C1 => n2075, C2 => 
                           n2074, A => n2073, ZN => n2081);
   U2277 : OAI211_X1 port map( C1 => n2081, C2 => n2080, A => n2079, B => n2078
                           , ZN => cu_i_n209);
   U2278 : NOR2_X1 port map( A1 => cu_i_n123, A2 => cu_i_n23, ZN => cu_i_n210);
   U2279 : AOI22_X1 port map( A1 => n704, A2 => n699, B1 => n2318, B2 => n2084,
                           ZN => cu_i_n131);
   U2280 : MUX2_X1 port map( A => cu_i_cw2_6_port, B => cu_i_cw1_6_port, S => 
                           n2084, Z => cu_i_n127);
   U2281 : MUX2_X1 port map( A => cu_i_cw2_5_port, B => cu_i_cw1_5_port, S => 
                           n2084, Z => cu_i_n126);
   U2282 : MUX2_X1 port map( A => curr_instruction_to_cu_i_31_port, B => 
                           IRAM_DATA(31), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n69);
   U2283 : MUX2_X1 port map( A => curr_instruction_to_cu_i_30_port, B => 
                           IRAM_DATA(30), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n68);
   U2284 : MUX2_X1 port map( A => n2315, B => IRAM_DATA(29), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n67);
   U2285 : MUX2_X1 port map( A => curr_instruction_to_cu_i_28_port, B => 
                           IRAM_DATA(28), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n66);
   U2286 : MUX2_X1 port map( A => curr_instruction_to_cu_i_27_port, B => 
                           IRAM_DATA(27), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n65);
   U2287 : MUX2_X1 port map( A => curr_instruction_to_cu_i_26_port, B => 
                           IRAM_DATA(26), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n64);
   U2288 : MUX2_X1 port map( A => datapath_i_n9, B => IRAM_DATA(25), S => n2084
                           , Z => datapath_i_fetch_stage_dp_n63);
   U2289 : MUX2_X1 port map( A => datapath_i_n10, B => IRAM_DATA(24), S => 
                           n2308, Z => datapath_i_fetch_stage_dp_n62);
   U2290 : MUX2_X1 port map( A => datapath_i_n11, B => IRAM_DATA(23), S => 
                           n2084, Z => datapath_i_fetch_stage_dp_n61);
   U2291 : MUX2_X1 port map( A => datapath_i_n12, B => IRAM_DATA(22), S => 
                           n2084, Z => datapath_i_fetch_stage_dp_n60);
   U2292 : MUX2_X1 port map( A => datapath_i_n13, B => IRAM_DATA(21), S => 
                           n2084, Z => datapath_i_fetch_stage_dp_n59);
   U2293 : MUX2_X1 port map( A => curr_instruction_to_cu_i_20_port, B => 
                           IRAM_DATA(20), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n58);
   U2294 : MUX2_X1 port map( A => curr_instruction_to_cu_i_19_port, B => 
                           IRAM_DATA(19), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n57);
   U2295 : NAND2_X1 port map( A1 => n2308, A2 => IRAM_DATA(18), ZN => n2082);
   U2296 : OAI21_X1 port map( B1 => n2308, B2 => n697, A => n2082, ZN => 
                           datapath_i_fetch_stage_dp_n56);
   U2297 : MUX2_X1 port map( A => curr_instruction_to_cu_i_17_port, B => 
                           IRAM_DATA(17), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n55);
   U2298 : MUX2_X1 port map( A => curr_instruction_to_cu_i_16_port, B => 
                           IRAM_DATA(16), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n54);
   U2299 : MUX2_X1 port map( A => curr_instruction_to_cu_i_15_port, B => 
                           IRAM_DATA(15), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n53);
   U2300 : MUX2_X1 port map( A => curr_instruction_to_cu_i_14_port, B => 
                           IRAM_DATA(14), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n52);
   U2301 : NAND2_X1 port map( A1 => n2308, A2 => IRAM_DATA(13), ZN => n2083);
   U2302 : OAI21_X1 port map( B1 => n2308, B2 => n740, A => n2083, ZN => 
                           datapath_i_fetch_stage_dp_n51);
   U2303 : MUX2_X1 port map( A => curr_instruction_to_cu_i_12_port, B => 
                           IRAM_DATA(12), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n50);
   U2304 : MUX2_X1 port map( A => curr_instruction_to_cu_i_11_port, B => 
                           IRAM_DATA(11), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n49);
   U2305 : MUX2_X1 port map( A => datapath_i_n14, B => IRAM_DATA(10), S => 
                           n2084, Z => datapath_i_fetch_stage_dp_n48);
   U2306 : MUX2_X1 port map( A => datapath_i_n15, B => IRAM_DATA(9), S => n2084
                           , Z => datapath_i_fetch_stage_dp_n47);
   U2307 : MUX2_X1 port map( A => datapath_i_n16, B => IRAM_DATA(8), S => n2308
                           , Z => datapath_i_fetch_stage_dp_n46);
   U2308 : MUX2_X1 port map( A => datapath_i_n17, B => IRAM_DATA(7), S => n2084
                           , Z => datapath_i_fetch_stage_dp_n45);
   U2309 : MUX2_X1 port map( A => datapath_i_n18, B => IRAM_DATA(6), S => n2084
                           , Z => datapath_i_fetch_stage_dp_n44);
   U2310 : MUX2_X1 port map( A => curr_instruction_to_cu_i_5_port, B => 
                           IRAM_DATA(5), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n43);
   U2311 : MUX2_X1 port map( A => curr_instruction_to_cu_i_4_port, B => 
                           IRAM_DATA(4), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n42);
   U2312 : MUX2_X1 port map( A => curr_instruction_to_cu_i_3_port, B => 
                           IRAM_DATA(3), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n41);
   U2313 : MUX2_X1 port map( A => curr_instruction_to_cu_i_2_port, B => 
                           IRAM_DATA(2), S => n2308, Z => 
                           datapath_i_fetch_stage_dp_n40);
   U2314 : MUX2_X1 port map( A => curr_instruction_to_cu_i_1_port, B => 
                           IRAM_DATA(1), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n39);
   U2315 : MUX2_X1 port map( A => curr_instruction_to_cu_i_0_port, B => 
                           IRAM_DATA(0), S => n2084, Z => 
                           datapath_i_fetch_stage_dp_n38);
   U2316 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_0_port, 
                           B2 => n2177, ZN => n2085);
   U2317 : OAI21_X1 port map( B1 => n733, B2 => n2180, A => n2085, ZN => 
                           datapath_i_fetch_stage_dp_N5);
   U2318 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N39_port, B => 
                           datapath_i_fetch_stage_dp_N5, S => n2090, Z => 
                           datapath_i_fetch_stage_dp_n37);
   U2319 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_1_port, 
                           B2 => n2177, ZN => n2086);
   U2320 : OAI21_X1 port map( B1 => n734, B2 => n2180, A => n2086, ZN => 
                           datapath_i_fetch_stage_dp_N6);
   U2321 : MUX2_X1 port map( A => datapath_i_fetch_stage_dp_N40_port, B => 
                           datapath_i_fetch_stage_dp_N6, S => n2090, Z => 
                           datapath_i_fetch_stage_dp_n36);
   U2322 : OAI21_X1 port map( B1 => IRAM_ENABLE_port, B2 => IRAM_ADDRESS_2_port
                           , A => n2087, ZN => n2088);
   U2323 : AOI22_X1 port map( A1 => n2186, A2 => n2088, B1 => 
                           datapath_i_new_pc_value_mem_stage_i_2_port, B2 => 
                           n2183, ZN => datapath_i_fetch_stage_dp_n35);
   U2324 : OAI21_X1 port map( B1 => n2089, B2 => IRAM_ADDRESS_3_port, A => 
                           n2138, ZN => n2092);
   U2325 : AND2_X1 port map( A1 => datapath_i_new_pc_value_mem_stage_i_2_port, 
                           A2 => datapath_i_new_pc_value_mem_stage_i_3_port, ZN
                           => n2094);
   U2326 : OAI21_X1 port map( B1 => datapath_i_new_pc_value_mem_stage_i_2_port,
                           B2 => datapath_i_new_pc_value_mem_stage_i_3_port, A 
                           => n2090, ZN => n2091);
   U2327 : OAI22_X1 port map( A1 => n2096, A2 => n2092, B1 => n2094, B2 => 
                           n2091, ZN => datapath_i_fetch_stage_dp_n34);
   U2328 : OAI211_X1 port map( C1 => n2094, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_4_port, A => 
                           n2183, B => n2093, ZN => n2098);
   U2329 : OAI211_X1 port map( C1 => n2096, C2 => IRAM_ADDRESS_4_port, A => 
                           n2186, B => n2095, ZN => n2097);
   U2330 : NAND2_X1 port map( A1 => n2098, A2 => n2097, ZN => 
                           datapath_i_fetch_stage_dp_n33);
   U2331 : OAI211_X1 port map( C1 => n2100, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_6_port, A => 
                           n2183, B => n2099, ZN => n2104);
   U2332 : OAI211_X1 port map( C1 => n2102, C2 => IRAM_ADDRESS_6_port, A => 
                           n2186, B => n2101, ZN => n2103);
   U2333 : NAND2_X1 port map( A1 => n2104, A2 => n2103, ZN => 
                           datapath_i_fetch_stage_dp_n31);
   U2334 : OAI211_X1 port map( C1 => n2106, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_8_port, A => 
                           n2183, B => n2105, ZN => n2110);
   U2335 : OAI211_X1 port map( C1 => n2108, C2 => IRAM_ADDRESS_8_port, A => 
                           n2186, B => n2107, ZN => n2109);
   U2336 : NAND2_X1 port map( A1 => n2110, A2 => n2109, ZN => 
                           datapath_i_fetch_stage_dp_n29);
   U2337 : OAI211_X1 port map( C1 => n2112, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_10_port, A => 
                           n2183, B => n2111, ZN => n2116);
   U2338 : OAI211_X1 port map( C1 => n2114, C2 => IRAM_ADDRESS_10_port, A => 
                           n2186, B => n2113, ZN => n2115);
   U2339 : NAND2_X1 port map( A1 => n2116, A2 => n2115, ZN => 
                           datapath_i_fetch_stage_dp_n27);
   U2340 : OAI211_X1 port map( C1 => n2118, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_12_port, A => 
                           n2183, B => n2117, ZN => n2122);
   U2341 : OAI211_X1 port map( C1 => n2120, C2 => IRAM_ADDRESS_12_port, A => 
                           n2138, B => n2119, ZN => n2121);
   U2342 : NAND2_X1 port map( A1 => n2122, A2 => n2121, ZN => 
                           datapath_i_fetch_stage_dp_n25);
   U2343 : OAI211_X1 port map( C1 => n2124, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_14_port, A => 
                           n2183, B => n2123, ZN => n2128);
   U2344 : OAI211_X1 port map( C1 => n2126, C2 => IRAM_ADDRESS_14_port, A => 
                           n2138, B => n2125, ZN => n2127);
   U2345 : NAND2_X1 port map( A1 => n2128, A2 => n2127, ZN => 
                           datapath_i_fetch_stage_dp_n23);
   U2346 : OAI211_X1 port map( C1 => n2130, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_16_port, A => 
                           n2183, B => n2129, ZN => n2134);
   U2347 : OAI211_X1 port map( C1 => n2132, C2 => IRAM_ADDRESS_16_port, A => 
                           n2138, B => n2131, ZN => n2133);
   U2348 : NAND2_X1 port map( A1 => n2134, A2 => n2133, ZN => 
                           datapath_i_fetch_stage_dp_n21);
   U2349 : OAI211_X1 port map( C1 => n2136, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_18_port, A => 
                           n2183, B => n2135, ZN => n2141);
   U2350 : OAI211_X1 port map( C1 => n2139, C2 => IRAM_ADDRESS_18_port, A => 
                           n2138, B => n2137, ZN => n2140);
   U2351 : NAND2_X1 port map( A1 => n2141, A2 => n2140, ZN => 
                           datapath_i_fetch_stage_dp_n19);
   U2352 : OAI211_X1 port map( C1 => n2143, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_20_port, A => 
                           n2183, B => n2142, ZN => n2147);
   U2353 : OAI211_X1 port map( C1 => n2145, C2 => IRAM_ADDRESS_20_port, A => 
                           n2186, B => n2144, ZN => n2146);
   U2354 : NAND2_X1 port map( A1 => n2147, A2 => n2146, ZN => 
                           datapath_i_fetch_stage_dp_n17);
   U2355 : OAI211_X1 port map( C1 => n2149, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_22_port, A => 
                           n2183, B => n2148, ZN => n2153);
   U2356 : OAI211_X1 port map( C1 => n2151, C2 => IRAM_ADDRESS_22_port, A => 
                           n2186, B => n2150, ZN => n2152);
   U2357 : NAND2_X1 port map( A1 => n2153, A2 => n2152, ZN => 
                           datapath_i_fetch_stage_dp_n15);
   U2358 : OAI211_X1 port map( C1 => n2155, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_24_port, A => 
                           n2183, B => n2154, ZN => n2159);
   U2359 : OAI211_X1 port map( C1 => n2157, C2 => IRAM_ADDRESS_24_port, A => 
                           n2186, B => n2156, ZN => n2158);
   U2360 : NAND2_X1 port map( A1 => n2159, A2 => n2158, ZN => 
                           datapath_i_fetch_stage_dp_n13);
   U2361 : OAI211_X1 port map( C1 => n2161, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_26_port, A => 
                           n2183, B => n2160, ZN => n2165);
   U2362 : OAI211_X1 port map( C1 => n2163, C2 => IRAM_ADDRESS_26_port, A => 
                           n2186, B => n2162, ZN => n2164);
   U2363 : NAND2_X1 port map( A1 => n2165, A2 => n2164, ZN => 
                           datapath_i_fetch_stage_dp_n11);
   U2364 : OAI211_X1 port map( C1 => n2167, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_28_port, A => 
                           n2183, B => n2166, ZN => n2171);
   U2365 : OAI211_X1 port map( C1 => n2169, C2 => IRAM_ADDRESS_28_port, A => 
                           n2186, B => n2168, ZN => n2170);
   U2366 : NAND2_X1 port map( A1 => n2171, A2 => n2170, ZN => 
                           datapath_i_fetch_stage_dp_n9);
   U2367 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n2178, B1 => datapath_i_alu_output_val_i_30_port,
                           B2 => n2177, ZN => n2172);
   U2368 : OAI21_X1 port map( B1 => n727, B2 => n2180, A => n2172, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_30_port);
   U2369 : NAND2_X1 port map( A1 => n2173, A2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, ZN => 
                           n2182);
   U2370 : OAI211_X1 port map( C1 => n2173, C2 => 
                           datapath_i_new_pc_value_mem_stage_i_30_port, A => 
                           n2183, B => n2182, ZN => n2176);
   U2371 : NAND2_X1 port map( A1 => n2174, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n2181);
   U2372 : OAI211_X1 port map( C1 => n2174, C2 => IRAM_ADDRESS_30_port, A => 
                           n2186, B => n2181, ZN => n2175);
   U2373 : NAND2_X1 port map( A1 => n2176, A2 => n2175, ZN => 
                           datapath_i_fetch_stage_dp_n3);
   U2374 : AOI22_X1 port map( A1 => n2178, A2 => 
                           datapath_i_new_pc_value_decode_31_port, B1 => 
                           datapath_i_alu_output_val_i_31_port, B2 => n2177, ZN
                           => n2179);
   U2375 : OAI21_X1 port map( B1 => n703, B2 => n2180, A => n2179, ZN => 
                           datapath_i_new_pc_value_mem_stage_i_31_port);
   U2376 : XOR2_X1 port map( A => IRAM_ADDRESS_31_port, B => n2181, Z => n2185)
                           ;
   U2377 : XOR2_X1 port map( A => datapath_i_new_pc_value_mem_stage_i_31_port, 
                           B => n2182, Z => n2184);
   U2378 : AOI22_X1 port map( A1 => n2186, A2 => n2185, B1 => n2184, B2 => 
                           n2183, ZN => datapath_i_fetch_stage_dp_n2);
   U2379 : OAI21_X1 port map( B1 => n737, B2 => n2187, A => n2188, ZN => 
                           read_rf_p2_i);
   U2380 : OAI221_X1 port map( B1 => n2189, B2 => n697, C1 => n2188, C2 => n740
                           , A => n2232, ZN => datapath_i_decode_stage_dp_n78);
   U2381 : AND4_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_3_port, 
                           A2 => 
                           datapath_i_decode_stage_dp_address_rf_write_1_port, 
                           A3 => 
                           datapath_i_decode_stage_dp_address_rf_write_0_port, 
                           A4 => 
                           datapath_i_decode_stage_dp_address_rf_write_2_port, 
                           ZN => n2190);
   U2382 : AND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_address_rf_write_4_port, 
                           A2 => n2190, ZN => n2206);
   U2383 : INV_X1 port map( A => n2206, ZN => n2215);
   U2384 : AND2_X2 port map( A1 => n2215, A2 => n2193, ZN => n2229);
   U2385 : NOR2_X1 port map( A1 => n2206, A2 => n2193, ZN => n2228);
   U2386 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_0_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_0_port, ZN => n2194
                           );
   U2387 : OAI21_X1 port map( B1 => n733, B2 => n2215, A => n2194, ZN => 
                           datapath_i_decode_stage_dp_n43);
   U2388 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_1_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_1_port, ZN => n2195
                           );
   U2389 : OAI21_X1 port map( B1 => n734, B2 => n2215, A => n2195, ZN => 
                           datapath_i_decode_stage_dp_n42);
   U2390 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_2_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_2_port, ZN => n2196
                           );
   U2391 : OAI21_X1 port map( B1 => n728, B2 => n2215, A => n2196, ZN => 
                           datapath_i_decode_stage_dp_n41);
   U2392 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_3_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_3_port, ZN => n2197
                           );
   U2393 : OAI21_X1 port map( B1 => n729, B2 => n2215, A => n2197, ZN => 
                           datapath_i_decode_stage_dp_n40);
   U2394 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_4_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_4_port, ZN => n2198
                           );
   U2395 : OAI21_X1 port map( B1 => n730, B2 => n2215, A => n2198, ZN => 
                           datapath_i_decode_stage_dp_n39);
   U2396 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_5_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_5_port, ZN => n2199
                           );
   U2397 : OAI21_X1 port map( B1 => n731, B2 => n2215, A => n2199, ZN => 
                           datapath_i_decode_stage_dp_n38);
   U2398 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_6_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_6_port, ZN => n2200
                           );
   U2399 : OAI21_X1 port map( B1 => n732, B2 => n2215, A => n2200, ZN => 
                           datapath_i_decode_stage_dp_n37);
   U2400 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_7_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_7_port, ZN => n2201
                           );
   U2401 : OAI21_X1 port map( B1 => n705, B2 => n2215, A => n2201, ZN => 
                           datapath_i_decode_stage_dp_n36);
   U2402 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_8_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_8_port, ZN => n2202
                           );
   U2403 : OAI21_X1 port map( B1 => n706, B2 => n2215, A => n2202, ZN => 
                           datapath_i_decode_stage_dp_n35);
   U2404 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_9_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_9_port, ZN => n2203
                           );
   U2405 : OAI21_X1 port map( B1 => n707, B2 => n2215, A => n2203, ZN => 
                           datapath_i_decode_stage_dp_n34);
   U2406 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_10_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_10_port, ZN => 
                           n2204);
   U2407 : OAI21_X1 port map( B1 => n708, B2 => n2215, A => n2204, ZN => 
                           datapath_i_decode_stage_dp_n33);
   U2408 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_11_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_11_port, ZN => 
                           n2205);
   U2409 : OAI21_X1 port map( B1 => n709, B2 => n2215, A => n2205, ZN => 
                           datapath_i_decode_stage_dp_n32);
   U2410 : INV_X1 port map( A => n2206, ZN => n2231);
   U2411 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_12_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_12_port, ZN => 
                           n2207);
   U2412 : OAI21_X1 port map( B1 => n710, B2 => n2231, A => n2207, ZN => 
                           datapath_i_decode_stage_dp_n31);
   U2413 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_13_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_13_port, ZN => 
                           n2208);
   U2414 : OAI21_X1 port map( B1 => n711, B2 => n2215, A => n2208, ZN => 
                           datapath_i_decode_stage_dp_n30);
   U2415 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_14_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_14_port, ZN => 
                           n2209);
   U2416 : OAI21_X1 port map( B1 => n712, B2 => n2231, A => n2209, ZN => 
                           datapath_i_decode_stage_dp_n29);
   U2417 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_15_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_15_port, ZN => 
                           n2210);
   U2418 : OAI21_X1 port map( B1 => n713, B2 => n2215, A => n2210, ZN => 
                           datapath_i_decode_stage_dp_n28);
   U2419 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_16_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_16_port, ZN => 
                           n2211);
   U2420 : OAI21_X1 port map( B1 => n714, B2 => n2231, A => n2211, ZN => 
                           datapath_i_decode_stage_dp_n27);
   U2421 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_17_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_17_port, ZN => 
                           n2212);
   U2422 : OAI21_X1 port map( B1 => n715, B2 => n2215, A => n2212, ZN => 
                           datapath_i_decode_stage_dp_n26);
   U2423 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_18_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_18_port, ZN => 
                           n2213);
   U2424 : OAI21_X1 port map( B1 => n716, B2 => n2231, A => n2213, ZN => 
                           datapath_i_decode_stage_dp_n25);
   U2425 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_19_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_19_port, ZN => 
                           n2214);
   U2426 : OAI21_X1 port map( B1 => n717, B2 => n2215, A => n2214, ZN => 
                           datapath_i_decode_stage_dp_n24);
   U2427 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_20_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_20_port, ZN => 
                           n2216);
   U2428 : OAI21_X1 port map( B1 => n718, B2 => n2231, A => n2216, ZN => 
                           datapath_i_decode_stage_dp_n23);
   U2429 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_21_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_21_port, ZN => 
                           n2217);
   U2430 : OAI21_X1 port map( B1 => n719, B2 => n2231, A => n2217, ZN => 
                           datapath_i_decode_stage_dp_n22);
   U2431 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_22_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_22_port, ZN => 
                           n2218);
   U2432 : OAI21_X1 port map( B1 => n720, B2 => n2231, A => n2218, ZN => 
                           datapath_i_decode_stage_dp_n21);
   U2433 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_23_port, B1 => n2219, 
                           B2 => datapath_i_data_from_alu_i_23_port, ZN => 
                           n2220);
   U2434 : OAI21_X1 port map( B1 => n721, B2 => n2231, A => n2220, ZN => 
                           datapath_i_decode_stage_dp_n20);
   U2435 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_24_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_24_port, ZN => 
                           n2221);
   U2436 : OAI21_X1 port map( B1 => n722, B2 => n2231, A => n2221, ZN => 
                           datapath_i_decode_stage_dp_n19);
   U2437 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_25_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_25_port, ZN => 
                           n2222);
   U2438 : OAI21_X1 port map( B1 => n723, B2 => n2231, A => n2222, ZN => 
                           datapath_i_decode_stage_dp_n18);
   U2439 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_26_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_26_port, ZN => 
                           n2223);
   U2440 : OAI21_X1 port map( B1 => n691, B2 => n2231, A => n2223, ZN => 
                           datapath_i_decode_stage_dp_n17);
   U2441 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_27_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_27_port, ZN => 
                           n2224);
   U2442 : OAI21_X1 port map( B1 => n724, B2 => n2231, A => n2224, ZN => 
                           datapath_i_decode_stage_dp_n16);
   U2443 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_28_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_28_port, ZN => 
                           n2225);
   U2444 : OAI21_X1 port map( B1 => n725, B2 => n2231, A => n2225, ZN => 
                           datapath_i_decode_stage_dp_n15);
   U2445 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_29_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_29_port, ZN => 
                           n2226);
   U2446 : OAI21_X1 port map( B1 => n726, B2 => n2231, A => n2226, ZN => 
                           datapath_i_decode_stage_dp_n14);
   U2447 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_30_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_30_port, ZN => 
                           n2227);
   U2448 : OAI21_X1 port map( B1 => n727, B2 => n2231, A => n2227, ZN => 
                           datapath_i_decode_stage_dp_n13);
   U2449 : AOI22_X1 port map( A1 => n2229, A2 => 
                           datapath_i_data_from_memory_i_31_port, B1 => n2228, 
                           B2 => datapath_i_data_from_alu_i_31_port, ZN => 
                           n2230);
   U2450 : OAI21_X1 port map( B1 => n703, B2 => n2231, A => n2230, ZN => 
                           datapath_i_decode_stage_dp_n12);
   U2451 : OAI21_X1 port map( B1 => curr_instruction_to_cu_i_26_port, B2 => 
                           n2233, A => n2232, ZN => cu_i_cmd_word_6_port);
   U2452 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_6_port, B1 => 
                           cu_i_cw1_10_port, B2 => n2308, ZN => n2247);
   U2453 : NOR4_X1 port map( A1 => datapath_i_val_a_i_14_port, A2 => 
                           datapath_i_val_a_i_15_port, A3 => 
                           datapath_i_val_a_i_16_port, A4 => 
                           datapath_i_val_a_i_17_port, ZN => n2237);
   U2454 : NOR4_X1 port map( A1 => datapath_i_val_a_i_18_port, A2 => 
                           datapath_i_val_a_i_19_port, A3 => 
                           datapath_i_val_a_i_20_port, A4 => 
                           datapath_i_val_a_i_21_port, ZN => n2236);
   U2455 : NOR4_X1 port map( A1 => datapath_i_val_a_i_26_port, A2 => 
                           datapath_i_val_a_i_7_port, A3 => 
                           datapath_i_val_a_i_8_port, A4 => 
                           datapath_i_val_a_i_9_port, ZN => n2235);
   U2456 : NOR4_X1 port map( A1 => datapath_i_val_a_i_10_port, A2 => 
                           datapath_i_val_a_i_11_port, A3 => 
                           datapath_i_val_a_i_12_port, A4 => 
                           datapath_i_val_a_i_13_port, ZN => n2234);
   U2457 : NAND4_X1 port map( A1 => n2237, A2 => n2236, A3 => n2235, A4 => 
                           n2234, ZN => n2243);
   U2458 : NOR4_X1 port map( A1 => datapath_i_val_a_i_30_port, A2 => 
                           datapath_i_val_a_i_31_port, A3 => 
                           datapath_i_val_a_i_1_port, A4 => 
                           datapath_i_val_a_i_2_port, ZN => n2241);
   U2459 : NOR4_X1 port map( A1 => datapath_i_val_a_i_3_port, A2 => 
                           datapath_i_val_a_i_4_port, A3 => 
                           datapath_i_val_a_i_5_port, A4 => 
                           datapath_i_val_a_i_6_port, ZN => n2240);
   U2460 : NOR4_X1 port map( A1 => datapath_i_val_a_i_22_port, A2 => 
                           datapath_i_val_a_i_23_port, A3 => 
                           datapath_i_val_a_i_24_port, A4 => 
                           datapath_i_val_a_i_25_port, ZN => n2239);
   U2461 : NOR4_X1 port map( A1 => datapath_i_val_a_i_0_port, A2 => 
                           datapath_i_val_a_i_27_port, A3 => 
                           datapath_i_val_a_i_28_port, A4 => 
                           datapath_i_val_a_i_29_port, ZN => n2238);
   U2462 : NAND4_X1 port map( A1 => n2241, A2 => n2240, A3 => n2239, A4 => 
                           n2238, ZN => n2242);
   U2463 : NOR2_X1 port map( A1 => n2243, A2 => n2242, ZN => n2245);
   U2464 : AOI22_X1 port map( A1 => n704, A2 => cu_i_cmd_word_7_port, B1 => 
                           cu_i_cw1_11_port, B2 => n2308, ZN => n2244);
   U2465 : NAND2_X1 port map( A1 => n2245, A2 => n2244, ZN => n2246);
   U2466 : OAI22_X1 port map( A1 => n2247, A2 => n2246, B1 => n2245, B2 => 
                           n2244, ZN => 
                           datapath_i_execute_stage_dp_branch_taken_reg_q_0_port);
   U2467 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_7_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_7_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_7_port)
                           ;
   U2468 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_8_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_8_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_8_port)
                           ;
   U2469 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_9_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_9_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_9_port)
                           ;
   U2470 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_10_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_10_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_10_port
                           );
   U2471 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_11_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_11_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_11_port
                           );
   U2472 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_12_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_12_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_12_port
                           );
   U2473 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_13_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_13_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_13_port
                           );
   U2474 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_14_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_14_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_14_port
                           );
   U2475 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_15_port, 
                           ZN => n2248);
   U2476 : NAND2_X1 port map( A1 => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_31_port, 
                           A2 => n310, ZN => n2258);
   U2477 : OAI21_X1 port map( B1 => n310, B2 => n2248, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_15_port
                           );
   U2478 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_16_port, 
                           ZN => n2249);
   U2479 : OAI21_X1 port map( B1 => n2320, B2 => n2249, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_16_port
                           );
   U2480 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_17_port, 
                           ZN => n2250);
   U2481 : OAI21_X1 port map( B1 => n310, B2 => n2250, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_17_port
                           );
   U2482 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_18_port, 
                           ZN => n2251);
   U2483 : OAI21_X1 port map( B1 => n2320, B2 => n2251, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_18_port
                           );
   U2484 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_19_port, 
                           ZN => n2252);
   U2485 : OAI21_X1 port map( B1 => n310, B2 => n2252, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_19_port
                           );
   U2486 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_20_port, 
                           ZN => n2253);
   U2487 : OAI21_X1 port map( B1 => n2320, B2 => n2253, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_20_port
                           );
   U2488 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_21_port, 
                           ZN => n2254);
   U2489 : OAI21_X1 port map( B1 => n310, B2 => n2254, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_21_port
                           );
   U2490 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_22_port, 
                           ZN => n2255);
   U2491 : OAI21_X1 port map( B1 => n2320, B2 => n2255, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_22_port
                           );
   U2492 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_23_port, 
                           ZN => n2256);
   U2493 : OAI21_X1 port map( B1 => n310, B2 => n2256, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_23_port
                           );
   U2494 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_24_port, 
                           ZN => n2257);
   U2495 : OAI21_X1 port map( B1 => n2320, B2 => n2257, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_24_port
                           );
   U2496 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_0_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_0_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_0_port)
                           ;
   U2497 : INV_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_25_port, 
                           ZN => n2259);
   U2498 : OAI21_X1 port map( B1 => n310, B2 => n2259, A => n2258, ZN => 
                           datapath_i_decode_stage_dp_val_reg_immediate_31_port
                           );
   U2499 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_1_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_1_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_1_port)
                           ;
   U2500 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_2_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_2_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_2_port)
                           ;
   U2501 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_3_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_3_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_3_port)
                           ;
   U2502 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_4_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_4_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_4_port)
                           ;
   U2503 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_5_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_5_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_5_port)
                           ;
   U2504 : MUX2_X1 port map( A => 
                           datapath_i_decode_stage_dp_val_reg_immediate_i_6_port, B 
                           => 
                           datapath_i_decode_stage_dp_val_reg_immediate_j_6_port, S 
                           => n2260, Z => 
                           datapath_i_decode_stage_dp_val_reg_immediate_6_port)
                           ;
   U2505 : MUX2_X1 port map( A => datapath_i_val_b_i_7_port, B => 
                           datapath_i_val_immediate_i_7_port, S => n2261, Z => 
                           datapath_i_execute_stage_dp_opb_7_port);
   U2506 : MUX2_X1 port map( A => datapath_i_val_b_i_8_port, B => 
                           datapath_i_val_immediate_i_8_port, S => n2261, Z => 
                           datapath_i_execute_stage_dp_opb_8_port);
   U2507 : MUX2_X1 port map( A => datapath_i_val_b_i_9_port, B => 
                           datapath_i_val_immediate_i_9_port, S => n2261, Z => 
                           datapath_i_execute_stage_dp_opb_9_port);
   U2508 : MUX2_X1 port map( A => datapath_i_val_b_i_10_port, B => 
                           datapath_i_val_immediate_i_10_port, S => n2261, Z =>
                           datapath_i_execute_stage_dp_opb_10_port);
   U2509 : MUX2_X1 port map( A => datapath_i_val_b_i_11_port, B => 
                           datapath_i_val_immediate_i_11_port, S => n2261, Z =>
                           datapath_i_execute_stage_dp_opb_11_port);
   U2510 : MUX2_X1 port map( A => datapath_i_val_b_i_12_port, B => 
                           datapath_i_val_immediate_i_12_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_12_port);
   U2511 : MUX2_X1 port map( A => datapath_i_val_b_i_13_port, B => 
                           datapath_i_val_immediate_i_13_port, S => n2261, Z =>
                           datapath_i_execute_stage_dp_opb_13_port);
   U2512 : MUX2_X1 port map( A => datapath_i_val_b_i_14_port, B => 
                           datapath_i_val_immediate_i_14_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_14_port);
   U2513 : MUX2_X1 port map( A => datapath_i_val_b_i_15_port, B => 
                           datapath_i_val_immediate_i_15_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_15_port);
   U2514 : MUX2_X1 port map( A => datapath_i_val_b_i_16_port, B => 
                           datapath_i_val_immediate_i_16_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_16_port);
   U2515 : MUX2_X1 port map( A => datapath_i_val_b_i_17_port, B => 
                           datapath_i_val_immediate_i_17_port, S => n2261, Z =>
                           datapath_i_execute_stage_dp_opb_17_port);
   U2516 : MUX2_X1 port map( A => datapath_i_val_b_i_18_port, B => 
                           datapath_i_val_immediate_i_18_port, S => n2261, Z =>
                           datapath_i_execute_stage_dp_opb_18_port);
   U2517 : MUX2_X1 port map( A => datapath_i_val_b_i_19_port, B => 
                           datapath_i_val_immediate_i_19_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_19_port);
   U2518 : MUX2_X1 port map( A => datapath_i_val_b_i_20_port, B => 
                           datapath_i_val_immediate_i_20_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_20_port);
   U2519 : MUX2_X1 port map( A => datapath_i_val_b_i_21_port, B => 
                           datapath_i_val_immediate_i_21_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_21_port);
   U2520 : MUX2_X1 port map( A => datapath_i_val_b_i_22_port, B => 
                           datapath_i_val_immediate_i_22_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_22_port);
   U2521 : MUX2_X1 port map( A => datapath_i_val_b_i_23_port, B => 
                           datapath_i_val_immediate_i_23_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_23_port);
   U2522 : MUX2_X1 port map( A => datapath_i_val_b_i_24_port, B => 
                           datapath_i_val_immediate_i_24_port, S => n2263, Z =>
                           datapath_i_execute_stage_dp_opb_24_port);
   U2523 : NAND2_X1 port map( A1 => datapath_i_val_immediate_i_25_port, A2 => 
                           n2263, ZN => n2262);
   U2524 : OAI21_X1 port map( B1 => n758, B2 => n2263, A => n2262, ZN => 
                           datapath_i_execute_stage_dp_opb_25_port);
   U2525 : OAI21_X1 port map( B1 => n759, B2 => n2263, A => n2262, ZN => 
                           datapath_i_execute_stage_dp_opb_26_port);
   U2526 : OAI21_X1 port map( B1 => n760, B2 => n2263, A => n2262, ZN => 
                           datapath_i_execute_stage_dp_opb_27_port);
   U2527 : OAI21_X1 port map( B1 => n761, B2 => n2263, A => n2262, ZN => 
                           datapath_i_execute_stage_dp_opb_28_port);
   U2528 : OAI21_X1 port map( B1 => n762, B2 => n2263, A => n2262, ZN => 
                           datapath_i_execute_stage_dp_opb_29_port);
   U2529 : OAI21_X1 port map( B1 => n763, B2 => n2263, A => n2262, ZN => 
                           datapath_i_execute_stage_dp_opb_30_port);
   U2530 : OAI21_X1 port map( B1 => n764, B2 => n2263, A => n2262, ZN => 
                           datapath_i_execute_stage_dp_opb_31_port);
   U2531 : MUX2_X1 port map( A => datapath_i_val_b_i_4_port, B => 
                           datapath_i_val_immediate_i_4_port, S => n2263, Z => 
                           datapath_i_execute_stage_dp_opb_4_port);
   U2532 : MUX2_X1 port map( A => datapath_i_val_b_i_5_port, B => 
                           datapath_i_val_immediate_i_5_port, S => n2263, Z => 
                           datapath_i_execute_stage_dp_opb_5_port);
   U2533 : MUX2_X1 port map( A => datapath_i_val_b_i_6_port, B => 
                           datapath_i_val_immediate_i_6_port, S => n2263, Z => 
                           datapath_i_execute_stage_dp_opb_6_port);
   U2534 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_7_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_7_port, B2 => 
                           n2285, ZN => n2264);
   U2535 : OAI21_X1 port map( B1 => n705, B2 => n2300, A => n2264, ZN => 
                           datapath_i_execute_stage_dp_opa_7_port);
   U2536 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_8_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_8_port, B2 => 
                           n2297, ZN => n2265);
   U2537 : OAI21_X1 port map( B1 => n706, B2 => n2289, A => n2265, ZN => 
                           datapath_i_execute_stage_dp_opa_8_port);
   U2538 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_9_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_9_port, B2 => 
                           n2285, ZN => n2266);
   U2539 : OAI21_X1 port map( B1 => n707, B2 => n2300, A => n2266, ZN => 
                           datapath_i_execute_stage_dp_opa_9_port);
   U2540 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_10_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_10_port, B2 => 
                           n2297, ZN => n2267);
   U2541 : OAI21_X1 port map( B1 => n708, B2 => n2289, A => n2267, ZN => 
                           datapath_i_execute_stage_dp_opa_10_port);
   U2542 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_11_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_11_port, B2 => 
                           n2285, ZN => n2268);
   U2543 : OAI21_X1 port map( B1 => n709, B2 => n2300, A => n2268, ZN => 
                           datapath_i_execute_stage_dp_opa_11_port);
   U2544 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_12_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_12_port, B2 => 
                           n2297, ZN => n2269);
   U2545 : OAI21_X1 port map( B1 => n710, B2 => n2289, A => n2269, ZN => 
                           datapath_i_execute_stage_dp_opa_12_port);
   U2546 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_13_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_13_port, B2 => 
                           n2285, ZN => n2270);
   U2547 : OAI21_X1 port map( B1 => n711, B2 => n2300, A => n2270, ZN => 
                           datapath_i_execute_stage_dp_opa_13_port);
   U2548 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_14_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_14_port, B2 => 
                           n2297, ZN => n2271);
   U2549 : OAI21_X1 port map( B1 => n712, B2 => n2289, A => n2271, ZN => 
                           datapath_i_execute_stage_dp_opa_14_port);
   U2550 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_15_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_15_port, B2 => 
                           n2285, ZN => n2272);
   U2551 : OAI21_X1 port map( B1 => n713, B2 => n2300, A => n2272, ZN => 
                           datapath_i_execute_stage_dp_opa_15_port);
   U2552 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_16_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_16_port, B2 => 
                           n2285, ZN => n2273);
   U2553 : OAI21_X1 port map( B1 => n714, B2 => n2300, A => n2273, ZN => 
                           datapath_i_execute_stage_dp_opa_16_port);
   U2554 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_17_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_17_port, B2 => 
                           n2297, ZN => n2274);
   U2555 : OAI21_X1 port map( B1 => n715, B2 => n2300, A => n2274, ZN => 
                           datapath_i_execute_stage_dp_opa_17_port);
   U2556 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_18_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_18_port, B2 => 
                           n2285, ZN => n2275);
   U2557 : OAI21_X1 port map( B1 => n716, B2 => n2289, A => n2275, ZN => 
                           datapath_i_execute_stage_dp_opa_18_port);
   U2558 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_19_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_19_port, B2 => 
                           n2297, ZN => n2276);
   U2559 : OAI21_X1 port map( B1 => n717, B2 => n2289, A => n2276, ZN => 
                           datapath_i_execute_stage_dp_opa_19_port);
   U2560 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_20_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_20_port, B2 => 
                           n2285, ZN => n2277);
   U2561 : OAI21_X1 port map( B1 => n718, B2 => n2289, A => n2277, ZN => 
                           datapath_i_execute_stage_dp_opa_20_port);
   U2562 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_21_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_21_port, B2 => 
                           n2297, ZN => n2278);
   U2563 : OAI21_X1 port map( B1 => n719, B2 => n2289, A => n2278, ZN => 
                           datapath_i_execute_stage_dp_opa_21_port);
   U2564 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_22_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_22_port, B2 => 
                           n2285, ZN => n2279);
   U2565 : OAI21_X1 port map( B1 => n720, B2 => n2289, A => n2279, ZN => 
                           datapath_i_execute_stage_dp_opa_22_port);
   U2566 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_23_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_23_port, B2 => 
                           n2285, ZN => n2280);
   U2567 : OAI21_X1 port map( B1 => n721, B2 => n2289, A => n2280, ZN => 
                           datapath_i_execute_stage_dp_opa_23_port);
   U2568 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_24_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_24_port, B2 => 
                           n2285, ZN => n2281);
   U2569 : OAI21_X1 port map( B1 => n722, B2 => n2289, A => n2281, ZN => 
                           datapath_i_execute_stage_dp_opa_24_port);
   U2570 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_25_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_25_port, B2 => 
                           n2285, ZN => n2282);
   U2571 : OAI21_X1 port map( B1 => n723, B2 => n2289, A => n2282, ZN => 
                           datapath_i_execute_stage_dp_opa_25_port);
   U2572 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_0_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_0_port, B2 => 
                           n2285, ZN => n2283);
   U2573 : OAI21_X1 port map( B1 => n733, B2 => n2289, A => n2283, ZN => 
                           datapath_i_execute_stage_dp_opa_0_port);
   U2574 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_27_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_27_port, B2 => 
                           n2285, ZN => n2284);
   U2575 : OAI21_X1 port map( B1 => n724, B2 => n2289, A => n2284, ZN => 
                           datapath_i_execute_stage_dp_opa_27_port);
   U2576 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_28_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_28_port, B2 => 
                           n2285, ZN => n2286);
   U2577 : OAI21_X1 port map( B1 => n725, B2 => n2289, A => n2286, ZN => 
                           datapath_i_execute_stage_dp_opa_28_port);
   U2578 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_29_port, A2 
                           => n2287, B1 => datapath_i_val_a_i_29_port, B2 => 
                           n2297, ZN => n2288);
   U2579 : OAI21_X1 port map( B1 => n726, B2 => n2289, A => n2288, ZN => 
                           datapath_i_execute_stage_dp_opa_29_port);
   U2580 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_30_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_30_port, B2 => 
                           n2297, ZN => n2290);
   U2581 : OAI21_X1 port map( B1 => n727, B2 => n2300, A => n2290, ZN => 
                           datapath_i_execute_stage_dp_opa_30_port);
   U2582 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_31_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_31_port, B2 => 
                           n2297, ZN => n2291);
   U2583 : OAI21_X1 port map( B1 => n703, B2 => n2300, A => n2291, ZN => 
                           datapath_i_execute_stage_dp_opa_31_port);
   U2584 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_1_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_1_port, B2 => 
                           n2297, ZN => n2292);
   U2585 : OAI21_X1 port map( B1 => n734, B2 => n2300, A => n2292, ZN => 
                           datapath_i_execute_stage_dp_opa_1_port);
   U2586 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_2_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_2_port, B2 => 
                           n2297, ZN => n2293);
   U2587 : OAI21_X1 port map( B1 => n728, B2 => n2300, A => n2293, ZN => 
                           datapath_i_execute_stage_dp_opa_2_port);
   U2588 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_3_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_3_port, B2 => 
                           n2297, ZN => n2294);
   U2589 : OAI21_X1 port map( B1 => n729, B2 => n2300, A => n2294, ZN => 
                           datapath_i_execute_stage_dp_opa_3_port);
   U2590 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_4_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_4_port, B2 => 
                           n2297, ZN => n2295);
   U2591 : OAI21_X1 port map( B1 => n730, B2 => n2300, A => n2295, ZN => 
                           datapath_i_execute_stage_dp_opa_4_port);
   U2592 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_5_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_5_port, B2 => 
                           n2297, ZN => n2296);
   U2593 : OAI21_X1 port map( B1 => n731, B2 => n2300, A => n2296, ZN => 
                           datapath_i_execute_stage_dp_opa_5_port);
   U2594 : AOI22_X1 port map( A1 => datapath_i_new_pc_value_decode_6_port, A2 
                           => n2298, B1 => datapath_i_val_a_i_6_port, B2 => 
                           n2297, ZN => n2299);
   U2595 : OAI21_X1 port map( B1 => n732, B2 => n2300, A => n2299, ZN => 
                           datapath_i_execute_stage_dp_opa_6_port);

end SYN_dlx_rtl;
