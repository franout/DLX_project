//
//					\\\ Sapere Aude ///
//
// -----------------------------------------------------------------------------
// Copyright (c) 2014-2020 All rights reserved
// -----------------------------------------------------------------------------
// Author : Angione Francesco s262620@studenti.polito.it franout@Github.com
// File   : dlx_driver.sv
// Create : 2020-09-01 21:57:00
// Revise : 2020-09-01 22:05:14
// Editor : sublime text3, tab size (4)
// Description :
// -----------------------------------------------------------------------------



`ifndef __DLX_DRIVER_SV
`define __DLX_DRIVER_SV

class driver extends uvm_driver #(reg_item);
  `uvm_component_utils(driver)
  function new(string name = "driver", uvm_component parent=null);
    super.new(name, parent);
  endfunction

  virtual reg_if vif;

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if (!uvm_config_db#(virtual reg_if)::get(this, "", "reg_vif", vif))
      `uvm_fatal("DRV", "Could not get vif")
  endfunction

  virtual task run_phase(uvm_phase phase);
    super.run_phase(phase);
    forever begin
      reg_item m_item;
      `uvm_info("DRV", $sformatf("Wait for item from sequencer"), UVM_LOW)
      seq_item_port.get_next_item(m_item);
      drive_item(m_item);
      seq_item_port.item_done();
    end
  endtask

  virtual task drive_item(reg_item m_item);
      vif.sel <= 1;
      vif.addr 	<= m_item.addr;
      vif.wr 	<= m_item.wr;
      vif.wdata <= m_item.wdata;
      @ (posedge vif.clk);
      while (!vif.ready)  begin
        `uvm_info("DRV", "Wait until ready is high", UVM_LOW)
        @(posedge vif.clk);
      end

      vif.sel <= 0;
  endtask
endclass

// data are usually generated by a generator class
class my_driver extends uvm_driver;
	`uvm_component_utils (my_driver)

	int unsigned      n_times;
	my_data           data_obj;
	virtual  dut_if   vif;

	function new (string name, uvm_component parent);
		super.new (name, parent);
	endfunction

	virtual function void build_phase (uvm_phase phase);
		super.build_phase (phase);
		if (! uvm_config_db #(virtual dut_if) :: get (this, "", "vif", vif)) begin
			`uvm_fatal (get_type_name (), "Didn't get handle to virtual interface dut_if")
		end
	endfunction

	// reset phase 
	task reset_phase (uvm_phase phase);
   super.reset_phase (phase);
   `uvm_info (get_type_name (), $sformatf ("Applying initial reset"), UVM_MEDIUM)
   this.vif.rstn = 0;
   repeat (20) @ (posedge vif.clk);
   this.vif.rstn = 1;
   `uvm_info (get_type_name (), $sformatf ("DUT is now out of reset"), UVM_MEDIUM)
endtask


task main_phase (uvm_phase phase);
	super.main_phase (phase);
	phase.raise_objection (phase);
	`uvm_info (get_type_name (), $sformatf ("Inside Main phase"), UVM_MEDIUM)

	// Let's create a data object, randomize it and send it to the DUT
	n_times = 5;
	repeat (n_times) begin
		`uvm_info (get_type_name (), $sformatf ("Generate and randomize data packet"), UVM_DEBUG)
		data_obj = my_data::type_id::create ("data_obj", this);
		assert(data_obj.randomize ());
		@(posedge vif.clk);
		`uvm_info (get_type_name (), $sformatf ("Drive data packet to DUT"), UVM_DEBUG)
		this.vif.en    = 1;
		this.vif.wr    = 1;
 			this.vif.addr  = data_obj.addr;
		this.vif.wdata = data_obj.data;
 			data_obj.display ();
 		end
	phase.drop_objection (phase);
endtask

`endif