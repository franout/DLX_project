--------------------------------------------------------------------------------
-- Title       : Fetch stage of datapath
-- Project     : DLX for Microelectronic Systems
--------------------------------------------------------------------------------
-- File        : a.b.a-Fetch.stage.vhd
-- Author      : Francesco Angione <s262620@studenti.polito.it>
-- Company     : Politecnico di Torino, Italy
-- Created     : Wed Jul 22 20:57:16 2020
-- Last update : Wed Jul 22 20:57:24 2020
-- Platform    : Default Part Number
-- Standard    : VHDL-2008 
--------------------------------------------------------------------------------
-- Copyright (c) 2020 Politecnico di Torino, Italy
-------------------------------------------------------------------------------
-- Description: 
--------------------------------------------------------------------------------

library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity fetch_stage is
  port (
	clock
  ) ;
end entity ; -- fetch_stage

architecture arch of fetch_stage is

begin

end architecture ; -- arch